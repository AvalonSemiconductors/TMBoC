magic
tech sky130B
magscale 1 2
timestamp 1677505263
<< viali >>
rect 35633 42313 35667 42347
rect 26617 42245 26651 42279
rect 27905 42245 27939 42279
rect 29837 42245 29871 42279
rect 41705 42245 41739 42279
rect 14289 42177 14323 42211
rect 15485 42177 15519 42211
rect 20637 42177 20671 42211
rect 22753 42177 22787 42211
rect 25421 42177 25455 42211
rect 27353 42177 27387 42211
rect 28365 42177 28399 42211
rect 30665 42177 30699 42211
rect 32321 42177 32355 42211
rect 34897 42177 34931 42211
rect 43361 42177 43395 42211
rect 19993 42109 20027 42143
rect 33793 42109 33827 42143
rect 37565 42109 37599 42143
rect 39129 42109 39163 42143
rect 43085 42109 43119 42143
rect 21465 42041 21499 42075
rect 31401 42041 31435 42075
rect 41153 42041 41187 42075
rect 20453 41973 20487 42007
rect 22109 41973 22143 42007
rect 22569 41973 22603 42007
rect 23397 41973 23431 42007
rect 23949 41973 23983 42007
rect 24777 41973 24811 42007
rect 25237 41973 25271 42007
rect 26065 41973 26099 42007
rect 27169 41973 27203 42007
rect 29101 41973 29135 42007
rect 30849 41973 30883 42007
rect 32505 41973 32539 42007
rect 33241 41973 33275 42007
rect 34253 41973 34287 42007
rect 35081 41973 35115 42007
rect 36093 41973 36127 42007
rect 36645 41973 36679 42007
rect 38117 41973 38151 42007
rect 38669 41973 38703 42007
rect 40141 41973 40175 42007
rect 40601 41973 40635 42007
rect 42073 41769 42107 41803
rect 38853 41701 38887 41735
rect 29745 41633 29779 41667
rect 31585 41633 31619 41667
rect 40141 41633 40175 41667
rect 19993 41565 20027 41599
rect 22293 41565 22327 41599
rect 22560 41565 22594 41599
rect 25053 41565 25087 41599
rect 25320 41565 25354 41599
rect 26893 41565 26927 41599
rect 27160 41565 27194 41599
rect 28733 41565 28767 41599
rect 31841 41565 31875 41599
rect 36010 41565 36044 41599
rect 36277 41565 36311 41599
rect 36921 41565 36955 41599
rect 37473 41565 37507 41599
rect 38669 41565 38703 41599
rect 42165 41565 42199 41599
rect 20260 41497 20294 41531
rect 29990 41497 30024 41531
rect 33517 41497 33551 41531
rect 33885 41497 33919 41531
rect 21373 41429 21407 41463
rect 23673 41429 23707 41463
rect 26433 41429 26467 41463
rect 28273 41429 28307 41463
rect 28917 41429 28951 41463
rect 31125 41429 31159 41463
rect 32965 41429 32999 41463
rect 34897 41429 34931 41463
rect 36737 41429 36771 41463
rect 37657 41429 37691 41463
rect 38209 41429 38243 41463
rect 39313 41429 39347 41463
rect 40325 41429 40359 41463
rect 40417 41429 40451 41463
rect 40785 41429 40819 41463
rect 41245 41429 41279 41463
rect 42625 41429 42659 41463
rect 43177 41429 43211 41463
rect 19717 41225 19751 41259
rect 22845 41225 22879 41259
rect 25329 41225 25363 41259
rect 27169 41225 27203 41259
rect 27537 41225 27571 41259
rect 29101 41225 29135 41259
rect 30665 41225 30699 41259
rect 33701 41225 33735 41259
rect 35081 41225 35115 41259
rect 40693 41225 40727 41259
rect 43177 41225 43211 41259
rect 21097 41157 21131 41191
rect 31033 41157 31067 41191
rect 39558 41157 39592 41191
rect 21189 41089 21223 41123
rect 23213 41089 23247 41123
rect 25697 41089 25731 41123
rect 28733 41089 28767 41123
rect 32321 41089 32355 41123
rect 32588 41089 32622 41123
rect 34713 41089 34747 41123
rect 35808 41089 35842 41123
rect 37740 41089 37774 41123
rect 41153 41089 41187 41123
rect 20269 41021 20303 41055
rect 21373 41021 21407 41055
rect 23305 41021 23339 41055
rect 23489 41021 23523 41055
rect 25789 41021 25823 41055
rect 25973 41021 26007 41055
rect 27629 41021 27663 41055
rect 27813 41021 27847 41055
rect 28457 41021 28491 41055
rect 28641 41021 28675 41055
rect 29653 41021 29687 41055
rect 31125 41021 31159 41055
rect 31309 41021 31343 41055
rect 34437 41021 34471 41055
rect 34621 41021 34655 41055
rect 35541 41021 35575 41055
rect 37473 41021 37507 41055
rect 39313 41021 39347 41055
rect 20729 40953 20763 40987
rect 24133 40953 24167 40987
rect 22385 40885 22419 40919
rect 24869 40885 24903 40919
rect 26617 40885 26651 40919
rect 30113 40885 30147 40919
rect 36921 40885 36955 40919
rect 38853 40885 38887 40919
rect 41337 40885 41371 40919
rect 41797 40885 41831 40919
rect 42625 40885 42659 40919
rect 19993 40681 20027 40715
rect 32229 40681 32263 40715
rect 35541 40681 35575 40715
rect 36921 40681 36955 40715
rect 37381 40681 37415 40715
rect 38577 40681 38611 40715
rect 40049 40681 40083 40715
rect 20729 40545 20763 40579
rect 24041 40545 24075 40579
rect 31585 40545 31619 40579
rect 36277 40545 36311 40579
rect 38025 40545 38059 40579
rect 39221 40545 39255 40579
rect 20637 40477 20671 40511
rect 25053 40477 25087 40511
rect 30849 40477 30883 40511
rect 31861 40477 31895 40511
rect 34069 40477 34103 40511
rect 35725 40477 35759 40511
rect 36553 40477 36587 40511
rect 41173 40477 41207 40511
rect 41429 40477 41463 40511
rect 23774 40409 23808 40443
rect 25298 40409 25332 40443
rect 26893 40409 26927 40443
rect 28733 40409 28767 40443
rect 28917 40409 28951 40443
rect 29101 40409 29135 40443
rect 31769 40409 31803 40443
rect 33824 40409 33858 40443
rect 34989 40409 35023 40443
rect 37841 40409 37875 40443
rect 18797 40341 18831 40375
rect 21005 40341 21039 40375
rect 21465 40341 21499 40375
rect 22201 40341 22235 40375
rect 22661 40341 22695 40375
rect 26433 40341 26467 40375
rect 27813 40341 27847 40375
rect 29837 40341 29871 40375
rect 30389 40341 30423 40375
rect 32689 40341 32723 40375
rect 36461 40341 36495 40375
rect 37749 40341 37783 40375
rect 38945 40341 38979 40375
rect 39037 40341 39071 40375
rect 41889 40341 41923 40375
rect 42441 40341 42475 40375
rect 42993 40341 43027 40375
rect 21465 40137 21499 40171
rect 30297 40137 30331 40171
rect 33609 40137 33643 40171
rect 34069 40137 34103 40171
rect 35357 40137 35391 40171
rect 41337 40137 41371 40171
rect 25329 40069 25363 40103
rect 25513 40069 25547 40103
rect 30941 40069 30975 40103
rect 31125 40069 31159 40103
rect 18981 40001 19015 40035
rect 19441 40001 19475 40035
rect 19625 40001 19659 40035
rect 20341 40001 20375 40035
rect 22937 40001 22971 40035
rect 24501 40001 24535 40035
rect 28724 40001 28758 40035
rect 30849 40001 30883 40035
rect 31585 40001 31619 40035
rect 31769 40001 31803 40035
rect 33149 40001 33183 40035
rect 33241 40001 33275 40035
rect 34253 40001 34287 40035
rect 36470 40001 36504 40035
rect 40877 40001 40911 40035
rect 41889 40001 41923 40035
rect 19533 39933 19567 39967
rect 20085 39933 20119 39967
rect 23029 39933 23063 39967
rect 23305 39933 23339 39967
rect 23765 39933 23799 39967
rect 24593 39933 24627 39967
rect 24869 39933 24903 39967
rect 28457 39933 28491 39967
rect 33057 39933 33091 39967
rect 36737 39933 36771 39967
rect 32413 39865 32447 39899
rect 39681 39865 39715 39899
rect 40325 39865 40359 39899
rect 22293 39797 22327 39831
rect 25697 39797 25731 39831
rect 26249 39797 26283 39831
rect 27261 39797 27295 39831
rect 27721 39797 27755 39831
rect 29837 39797 29871 39831
rect 31125 39797 31159 39831
rect 31585 39797 31619 39831
rect 34713 39797 34747 39831
rect 37565 39797 37599 39831
rect 38025 39797 38059 39831
rect 38669 39797 38703 39831
rect 39221 39797 39255 39831
rect 42625 39797 42659 39831
rect 43361 39797 43395 39831
rect 17785 39593 17819 39627
rect 18337 39593 18371 39627
rect 18889 39593 18923 39627
rect 20085 39593 20119 39627
rect 23121 39593 23155 39627
rect 23581 39593 23615 39627
rect 28641 39593 28675 39627
rect 36084 39593 36118 39627
rect 43269 39593 43303 39627
rect 20269 39525 20303 39559
rect 32229 39525 32263 39559
rect 35449 39525 35483 39559
rect 36737 39525 36771 39559
rect 26525 39457 26559 39491
rect 26801 39457 26835 39491
rect 28365 39457 28399 39491
rect 29837 39457 29871 39491
rect 35173 39457 35207 39491
rect 39221 39457 39255 39491
rect 39497 39457 39531 39491
rect 19625 39389 19659 39423
rect 21005 39389 21039 39423
rect 21261 39389 21295 39423
rect 23305 39389 23339 39423
rect 23673 39389 23707 39423
rect 24869 39389 24903 39423
rect 25053 39389 25087 39423
rect 25237 39389 25271 39423
rect 26433 39389 26467 39423
rect 27445 39389 27479 39423
rect 27629 39389 27663 39423
rect 28273 39389 28307 39423
rect 31421 39389 31455 39423
rect 31677 39389 31711 39423
rect 32873 39389 32907 39423
rect 33241 39389 33275 39423
rect 35081 39389 35115 39423
rect 36921 39389 36955 39423
rect 37013 39389 37047 39423
rect 38025 39389 38059 39423
rect 39129 39389 39163 39423
rect 40049 39389 40083 39423
rect 40305 39389 40339 39423
rect 41889 39389 41923 39423
rect 20545 39321 20579 39355
rect 27261 39321 27295 39355
rect 33057 39321 33091 39355
rect 33149 39321 33183 39355
rect 35909 39321 35943 39355
rect 36737 39321 36771 39355
rect 42134 39321 42168 39355
rect 19441 39253 19475 39287
rect 22385 39253 22419 39287
rect 25697 39253 25731 39287
rect 29101 39253 29135 39287
rect 30297 39253 30331 39287
rect 33425 39253 33459 39287
rect 33977 39253 34011 39287
rect 36109 39253 36143 39287
rect 36277 39253 36311 39287
rect 37565 39253 37599 39287
rect 41429 39253 41463 39287
rect 20361 39049 20395 39083
rect 24225 39049 24259 39083
rect 25046 39049 25080 39083
rect 29745 39049 29779 39083
rect 31033 39049 31067 39083
rect 31585 39049 31619 39083
rect 39313 39049 39347 39083
rect 41153 39049 41187 39083
rect 41797 39049 41831 39083
rect 43177 39049 43211 39083
rect 18788 38981 18822 39015
rect 20821 38981 20855 39015
rect 22385 38981 22419 39015
rect 27414 38981 27448 39015
rect 32873 38981 32907 39015
rect 34805 38981 34839 39015
rect 36829 38981 36863 39015
rect 38586 38981 38620 39015
rect 40049 38981 40083 39015
rect 40265 38981 40299 39015
rect 17509 38913 17543 38947
rect 22155 38913 22189 38947
rect 22293 38913 22327 38947
rect 22568 38913 22602 38947
rect 22661 38913 22695 38947
rect 24133 38913 24167 38947
rect 24409 38913 24443 38947
rect 24869 38913 24903 38947
rect 24961 38913 24995 38947
rect 25145 38913 25179 38947
rect 29009 38913 29043 38947
rect 29193 38913 29227 38947
rect 29285 38913 29319 38947
rect 30665 38913 30699 38947
rect 30849 38913 30883 38947
rect 31493 38913 31527 38947
rect 31677 38913 31711 38947
rect 33333 38913 33367 38947
rect 33609 38913 33643 38947
rect 33701 38913 33735 38947
rect 33977 38913 34011 38947
rect 34253 38913 34287 38947
rect 35265 38913 35299 38947
rect 35541 38913 35575 38947
rect 35633 38913 35667 38947
rect 35909 38913 35943 38947
rect 36093 38913 36127 38947
rect 36737 38913 36771 38947
rect 36921 38913 36955 38947
rect 41061 38913 41095 38947
rect 41245 38913 41279 38947
rect 18521 38845 18555 38879
rect 27169 38845 27203 38879
rect 38853 38845 38887 38879
rect 16957 38777 16991 38811
rect 19901 38777 19935 38811
rect 20545 38777 20579 38811
rect 22017 38777 22051 38811
rect 24409 38777 24443 38811
rect 29009 38777 29043 38811
rect 40417 38777 40451 38811
rect 42625 38777 42659 38811
rect 18061 38709 18095 38743
rect 21373 38709 21407 38743
rect 23213 38709 23247 38743
rect 25605 38709 25639 38743
rect 26433 38709 26467 38743
rect 28549 38709 28583 38743
rect 32321 38709 32355 38743
rect 37473 38709 37507 38743
rect 40233 38709 40267 38743
rect 16497 38505 16531 38539
rect 19441 38505 19475 38539
rect 21373 38505 21407 38539
rect 24593 38505 24627 38539
rect 28641 38505 28675 38539
rect 29193 38505 29227 38539
rect 29745 38505 29779 38539
rect 30573 38505 30607 38539
rect 31309 38505 31343 38539
rect 32781 38505 32815 38539
rect 35449 38505 35483 38539
rect 36645 38505 36679 38539
rect 38577 38505 38611 38539
rect 40325 38505 40359 38539
rect 27353 38437 27387 38471
rect 19993 38369 20027 38403
rect 22293 38369 22327 38403
rect 22753 38369 22787 38403
rect 23765 38369 23799 38403
rect 31493 38369 31527 38403
rect 41061 38369 41095 38403
rect 41521 38369 41555 38403
rect 17509 38301 17543 38335
rect 19809 38301 19843 38335
rect 19901 38301 19935 38335
rect 20729 38301 20763 38335
rect 20822 38301 20856 38335
rect 21005 38301 21039 38335
rect 21097 38301 21131 38335
rect 21235 38301 21269 38335
rect 21833 38301 21867 38335
rect 22477 38301 22511 38335
rect 22845 38301 22879 38335
rect 23949 38301 23983 38335
rect 24772 38301 24806 38335
rect 24961 38301 24995 38335
rect 25089 38301 25123 38335
rect 25237 38301 25271 38335
rect 26387 38301 26421 38335
rect 26745 38301 26779 38335
rect 26893 38301 26927 38335
rect 27997 38301 28031 38335
rect 28145 38301 28179 38335
rect 28365 38301 28399 38335
rect 28503 38301 28537 38335
rect 31677 38301 31711 38335
rect 31769 38301 31803 38335
rect 33333 38301 33367 38335
rect 33425 38301 33459 38335
rect 33701 38301 33735 38335
rect 33793 38301 33827 38335
rect 34897 38301 34931 38335
rect 35265 38301 35299 38335
rect 37013 38301 37047 38335
rect 37105 38301 37139 38335
rect 37381 38301 37415 38335
rect 37657 38301 37691 38335
rect 37841 38301 37875 38335
rect 40049 38301 40083 38335
rect 40141 38301 40175 38335
rect 41153 38301 41187 38335
rect 41981 38301 42015 38335
rect 42237 38301 42271 38335
rect 17776 38233 17810 38267
rect 24869 38233 24903 38267
rect 26525 38233 26559 38267
rect 26617 38233 26651 38267
rect 28273 38233 28307 38267
rect 29929 38233 29963 38267
rect 30113 38233 30147 38267
rect 35081 38233 35115 38267
rect 35173 38233 35207 38267
rect 39037 38233 39071 38267
rect 40325 38233 40359 38267
rect 17049 38165 17083 38199
rect 18889 38165 18923 38199
rect 25697 38165 25731 38199
rect 26249 38165 26283 38199
rect 36001 38165 36035 38199
rect 43361 38165 43395 38199
rect 18245 37961 18279 37995
rect 18889 37961 18923 37995
rect 19257 37961 19291 37995
rect 30665 37961 30699 37995
rect 31769 37961 31803 37995
rect 32321 37961 32355 37995
rect 34529 37961 34563 37995
rect 35817 37961 35851 37995
rect 36829 37961 36863 37995
rect 39497 37961 39531 37995
rect 40693 37961 40727 37995
rect 15209 37893 15243 37927
rect 20269 37893 20303 37927
rect 22293 37893 22327 37927
rect 22385 37893 22419 37927
rect 23581 37893 23615 37927
rect 25513 37893 25547 37927
rect 25605 37893 25639 37927
rect 26341 37893 26375 37927
rect 27629 37893 27663 37927
rect 28641 37893 28675 37927
rect 28733 37893 28767 37927
rect 34253 37893 34287 37927
rect 40417 37893 40451 37927
rect 41153 37893 41187 37927
rect 41353 37893 41387 37927
rect 18429 37825 18463 37859
rect 20913 37825 20947 37859
rect 21281 37825 21315 37859
rect 21465 37825 21499 37859
rect 22155 37825 22189 37859
rect 22513 37825 22547 37859
rect 22661 37825 22695 37859
rect 24225 37825 24259 37859
rect 24593 37825 24627 37859
rect 24777 37825 24811 37859
rect 25416 37825 25450 37859
rect 25733 37825 25767 37859
rect 25881 37825 25915 37859
rect 26525 37825 26559 37859
rect 26617 37825 26651 37859
rect 27261 37825 27295 37859
rect 27409 37825 27443 37859
rect 27537 37825 27571 37859
rect 27767 37825 27801 37859
rect 28365 37825 28399 37859
rect 28485 37825 28519 37859
rect 28830 37825 28864 37859
rect 29653 37825 29687 37859
rect 30481 37825 30515 37859
rect 30757 37825 30791 37859
rect 31217 37825 31251 37859
rect 31401 37825 31435 37859
rect 31493 37825 31527 37859
rect 31585 37825 31619 37859
rect 32505 37825 32539 37859
rect 32597 37825 32631 37859
rect 32781 37825 32815 37859
rect 32873 37825 32907 37859
rect 33885 37825 33919 37859
rect 33978 37825 34012 37859
rect 34161 37825 34195 37859
rect 34391 37825 34425 37859
rect 35173 37825 35207 37859
rect 35293 37825 35327 37859
rect 35449 37825 35483 37859
rect 35541 37825 35575 37859
rect 35679 37825 35713 37859
rect 36277 37825 36311 37859
rect 36461 37825 36495 37859
rect 36553 37825 36587 37859
rect 36645 37825 36679 37859
rect 38209 37825 38243 37859
rect 38485 37825 38519 37859
rect 38761 37825 38795 37859
rect 39037 37825 39071 37859
rect 39129 37825 39163 37859
rect 40049 37825 40083 37859
rect 40197 37825 40231 37859
rect 40325 37825 40359 37859
rect 40555 37825 40589 37859
rect 19349 37757 19383 37791
rect 19441 37757 19475 37791
rect 21005 37757 21039 37791
rect 24041 37757 24075 37791
rect 29745 37757 29779 37791
rect 41981 37757 42015 37791
rect 15761 37689 15795 37723
rect 17785 37689 17819 37723
rect 25237 37689 25271 37723
rect 26341 37689 26375 37723
rect 30481 37689 30515 37723
rect 33425 37689 33459 37723
rect 43177 37689 43211 37723
rect 16221 37621 16255 37655
rect 17141 37621 17175 37655
rect 22017 37621 22051 37655
rect 27905 37621 27939 37655
rect 29009 37621 29043 37655
rect 30021 37621 30055 37655
rect 37565 37621 37599 37655
rect 41337 37621 41371 37655
rect 41521 37621 41555 37655
rect 42625 37621 42659 37655
rect 14473 37417 14507 37451
rect 15577 37417 15611 37451
rect 16129 37417 16163 37451
rect 16681 37417 16715 37451
rect 17233 37417 17267 37451
rect 17785 37417 17819 37451
rect 24041 37417 24075 37451
rect 32965 37417 32999 37451
rect 36921 37417 36955 37451
rect 37473 37417 37507 37451
rect 40693 37417 40727 37451
rect 15025 37349 15059 37383
rect 18337 37349 18371 37383
rect 18889 37349 18923 37383
rect 41429 37349 41463 37383
rect 20821 37281 20855 37315
rect 21925 37281 21959 37315
rect 24593 37281 24627 37315
rect 25237 37281 25271 37315
rect 28089 37281 28123 37315
rect 28549 37281 28583 37315
rect 39313 37281 39347 37315
rect 19625 37213 19659 37247
rect 22017 37213 22051 37247
rect 22385 37213 22419 37247
rect 22569 37213 22603 37247
rect 23397 37213 23431 37247
rect 23490 37213 23524 37247
rect 23862 37213 23896 37247
rect 24869 37213 24903 37247
rect 25421 37213 25455 37247
rect 26433 37213 26467 37247
rect 26617 37213 26651 37247
rect 26985 37213 27019 37247
rect 27169 37213 27203 37247
rect 27629 37213 27663 37247
rect 28273 37213 28307 37247
rect 28641 37213 28675 37247
rect 29929 37213 29963 37247
rect 30185 37213 30219 37247
rect 31907 37213 31941 37247
rect 32045 37213 32079 37247
rect 32265 37213 32299 37247
rect 32413 37213 32447 37247
rect 33609 37213 33643 37247
rect 33702 37213 33736 37247
rect 33885 37213 33919 37247
rect 34115 37213 34149 37247
rect 34897 37213 34931 37247
rect 35045 37213 35079 37247
rect 35173 37213 35207 37247
rect 35265 37213 35299 37247
rect 35403 37213 35437 37247
rect 36369 37213 36403 37247
rect 36737 37213 36771 37247
rect 37841 37213 37875 37247
rect 38117 37213 38151 37247
rect 38209 37213 38243 37247
rect 38485 37213 38519 37247
rect 38669 37213 38703 37247
rect 40049 37213 40083 37247
rect 40197 37213 40231 37247
rect 40417 37213 40451 37247
rect 40555 37213 40589 37247
rect 41153 37213 41187 37247
rect 41245 37213 41279 37247
rect 41889 37213 41923 37247
rect 21373 37145 21407 37179
rect 23673 37145 23707 37179
rect 23765 37145 23799 37179
rect 25053 37145 25087 37179
rect 25973 37145 26007 37179
rect 32137 37145 32171 37179
rect 33977 37145 34011 37179
rect 36553 37145 36587 37179
rect 36645 37145 36679 37179
rect 40325 37145 40359 37179
rect 41429 37145 41463 37179
rect 42134 37145 42168 37179
rect 19441 37077 19475 37111
rect 20269 37077 20303 37111
rect 31309 37077 31343 37111
rect 31769 37077 31803 37111
rect 34253 37077 34287 37111
rect 35541 37077 35575 37111
rect 43269 37077 43303 37111
rect 14657 36873 14691 36907
rect 16313 36873 16347 36907
rect 18245 36873 18279 36907
rect 22753 36873 22787 36907
rect 23949 36873 23983 36907
rect 26433 36873 26467 36907
rect 28549 36873 28583 36907
rect 30481 36873 30515 36907
rect 33057 36873 33091 36907
rect 35633 36873 35667 36907
rect 36921 36873 36955 36907
rect 40785 36873 40819 36907
rect 41981 36873 42015 36907
rect 15761 36805 15795 36839
rect 24225 36805 24259 36839
rect 26065 36805 26099 36839
rect 26157 36805 26191 36839
rect 27445 36805 27479 36839
rect 33977 36805 34011 36839
rect 35265 36805 35299 36839
rect 36553 36805 36587 36839
rect 39681 36805 39715 36839
rect 40509 36805 40543 36839
rect 16865 36737 16899 36771
rect 17121 36737 17155 36771
rect 18797 36737 18831 36771
rect 19064 36737 19098 36771
rect 22477 36737 22511 36771
rect 24128 36737 24162 36771
rect 24317 36737 24351 36771
rect 24500 36737 24534 36771
rect 24593 36737 24627 36771
rect 25053 36737 25087 36771
rect 25237 36737 25271 36771
rect 25789 36737 25823 36771
rect 25882 36737 25916 36771
rect 26295 36737 26329 36771
rect 27353 36737 27387 36771
rect 27537 36737 27571 36771
rect 27721 36737 27755 36771
rect 28917 36737 28951 36771
rect 29285 36737 29319 36771
rect 29469 36737 29503 36771
rect 29929 36737 29963 36771
rect 30113 36737 30147 36771
rect 30205 36737 30239 36771
rect 30297 36737 30331 36771
rect 32505 36737 32539 36771
rect 32689 36737 32723 36771
rect 32781 36737 32815 36771
rect 32873 36737 32907 36771
rect 33701 36737 33735 36771
rect 33794 36737 33828 36771
rect 34069 36737 34103 36771
rect 34166 36737 34200 36771
rect 34989 36737 35023 36771
rect 35082 36737 35116 36771
rect 35357 36737 35391 36771
rect 35495 36737 35529 36771
rect 36369 36737 36403 36771
rect 36645 36737 36679 36771
rect 36737 36737 36771 36771
rect 38393 36737 38427 36771
rect 38577 36737 38611 36771
rect 38853 36737 38887 36771
rect 39129 36737 39163 36771
rect 39221 36737 39255 36771
rect 40141 36737 40175 36771
rect 40234 36737 40268 36771
rect 40417 36737 40451 36771
rect 40606 36737 40640 36771
rect 41245 36737 41279 36771
rect 41429 36737 41463 36771
rect 41889 36737 41923 36771
rect 42073 36737 42107 36771
rect 43361 36737 43395 36771
rect 21465 36669 21499 36703
rect 22109 36669 22143 36703
rect 22201 36669 22235 36703
rect 22569 36669 22603 36703
rect 28825 36669 28859 36703
rect 14105 36601 14139 36635
rect 15209 36601 15243 36635
rect 20913 36601 20947 36635
rect 34345 36601 34379 36635
rect 37565 36601 37599 36635
rect 20177 36533 20211 36567
rect 23489 36533 23523 36567
rect 25145 36533 25179 36567
rect 27169 36533 27203 36567
rect 31033 36533 31067 36567
rect 31585 36533 31619 36567
rect 41337 36533 41371 36567
rect 42625 36533 42659 36567
rect 43177 36533 43211 36567
rect 9689 36329 9723 36363
rect 17785 36329 17819 36363
rect 19441 36329 19475 36363
rect 21373 36329 21407 36363
rect 31309 36329 31343 36363
rect 32689 36329 32723 36363
rect 33701 36329 33735 36363
rect 35081 36329 35115 36363
rect 38945 36329 38979 36363
rect 40693 36329 40727 36363
rect 43361 36329 43395 36363
rect 21925 36261 21959 36295
rect 23489 36261 23523 36295
rect 26065 36261 26099 36295
rect 28457 36261 28491 36295
rect 37381 36261 37415 36295
rect 38485 36261 38519 36295
rect 16221 36193 16255 36227
rect 19901 36193 19935 36227
rect 20085 36193 20119 36227
rect 22569 36193 22603 36227
rect 31401 36193 31435 36227
rect 33793 36193 33827 36227
rect 9873 36125 9907 36159
rect 14289 36125 14323 36159
rect 16497 36125 16531 36159
rect 19809 36125 19843 36159
rect 22477 36125 22511 36159
rect 22845 36125 22879 36159
rect 23029 36125 23063 36159
rect 23673 36125 23707 36159
rect 24041 36125 24075 36159
rect 25237 36125 25271 36159
rect 25605 36125 25639 36159
rect 26249 36125 26283 36159
rect 26433 36125 26467 36159
rect 26617 36125 26651 36159
rect 27261 36125 27295 36159
rect 27629 36125 27663 36159
rect 29929 36125 29963 36159
rect 30297 36125 30331 36159
rect 30481 36125 30515 36159
rect 30757 36125 30791 36159
rect 31217 36125 31251 36159
rect 31585 36125 31619 36159
rect 33885 36125 33919 36159
rect 34897 36125 34931 36159
rect 35909 36125 35943 36159
rect 36737 36125 36771 36159
rect 36830 36125 36864 36159
rect 37013 36125 37047 36159
rect 37243 36125 37277 36159
rect 37841 36125 37875 36159
rect 37989 36125 38023 36159
rect 38209 36125 38243 36159
rect 38306 36125 38340 36159
rect 39129 36125 39163 36159
rect 39497 36125 39531 36159
rect 40049 36125 40083 36159
rect 40142 36125 40176 36159
rect 40417 36125 40451 36159
rect 40514 36125 40548 36159
rect 41153 36125 41187 36159
rect 41337 36125 41371 36159
rect 41981 36125 42015 36159
rect 14534 36057 14568 36091
rect 23765 36057 23799 36091
rect 23857 36057 23891 36091
rect 25329 36057 25363 36091
rect 25421 36057 25455 36091
rect 26341 36057 26375 36091
rect 27353 36057 27387 36091
rect 27445 36057 27479 36091
rect 28181 36057 28215 36091
rect 30665 36057 30699 36091
rect 32781 36057 32815 36091
rect 37105 36057 37139 36091
rect 38117 36057 38151 36091
rect 39221 36057 39255 36091
rect 39313 36057 39347 36091
rect 40325 36057 40359 36091
rect 42248 36057 42282 36091
rect 10425 35989 10459 36023
rect 15669 35989 15703 36023
rect 18797 35989 18831 36023
rect 20821 35989 20855 36023
rect 25053 35989 25087 36023
rect 27077 35989 27111 36023
rect 29101 35989 29135 36023
rect 33517 35989 33551 36023
rect 35725 35989 35759 36023
rect 41521 35989 41555 36023
rect 14565 35785 14599 35819
rect 16129 35785 16163 35819
rect 19993 35785 20027 35819
rect 20913 35785 20947 35819
rect 21465 35785 21499 35819
rect 23949 35785 23983 35819
rect 29193 35785 29227 35819
rect 30849 35785 30883 35819
rect 41153 35785 41187 35819
rect 42625 35785 42659 35819
rect 43269 35785 43303 35819
rect 22017 35717 22051 35751
rect 24593 35717 24627 35751
rect 25329 35717 25363 35751
rect 30021 35717 30055 35751
rect 32873 35717 32907 35751
rect 37749 35717 37783 35751
rect 38669 35717 38703 35751
rect 39681 35717 39715 35751
rect 15025 35649 15059 35683
rect 15945 35649 15979 35683
rect 17049 35649 17083 35683
rect 17141 35649 17175 35683
rect 17325 35649 17359 35683
rect 17785 35649 17819 35683
rect 18705 35649 18739 35683
rect 22293 35649 22327 35683
rect 22661 35649 22695 35683
rect 23029 35649 23063 35683
rect 23489 35649 23523 35683
rect 24225 35649 24259 35683
rect 26065 35649 26099 35683
rect 27445 35649 27479 35683
rect 28917 35649 28951 35683
rect 29791 35649 29825 35683
rect 29929 35649 29963 35683
rect 30204 35649 30238 35683
rect 30297 35649 30331 35683
rect 31309 35649 31343 35683
rect 31677 35649 31711 35683
rect 32689 35649 32723 35683
rect 32781 35649 32815 35683
rect 33057 35649 33091 35683
rect 34253 35649 34287 35683
rect 34897 35649 34931 35683
rect 35173 35649 35207 35683
rect 35817 35649 35851 35683
rect 36001 35649 36035 35683
rect 37473 35649 37507 35683
rect 37621 35649 37655 35683
rect 37841 35649 37875 35683
rect 37979 35649 38013 35683
rect 39405 35649 39439 35683
rect 39498 35649 39532 35683
rect 39773 35649 39807 35683
rect 39911 35649 39945 35683
rect 40509 35649 40543 35683
rect 40647 35649 40681 35683
rect 40785 35649 40819 35683
rect 40877 35649 40911 35683
rect 40974 35649 41008 35683
rect 41797 35649 41831 35683
rect 41981 35649 42015 35683
rect 42809 35649 42843 35683
rect 13461 35581 13495 35615
rect 18429 35581 18463 35615
rect 24133 35581 24167 35615
rect 24501 35581 24535 35615
rect 27353 35581 27387 35615
rect 27721 35581 27755 35615
rect 27813 35581 27847 35615
rect 28549 35581 28583 35615
rect 28641 35581 28675 35615
rect 29009 35581 29043 35615
rect 33977 35581 34011 35615
rect 34989 35581 35023 35615
rect 41613 35581 41647 35615
rect 15209 35513 15243 35547
rect 17969 35513 18003 35547
rect 26617 35513 26651 35547
rect 35357 35513 35391 35547
rect 35909 35513 35943 35547
rect 38117 35513 38151 35547
rect 14013 35445 14047 35479
rect 27169 35445 27203 35479
rect 29653 35445 29687 35479
rect 32505 35445 32539 35479
rect 34069 35445 34103 35479
rect 34437 35445 34471 35479
rect 34897 35445 34931 35479
rect 36645 35445 36679 35479
rect 40049 35445 40083 35479
rect 15485 35241 15519 35275
rect 16221 35241 16255 35275
rect 20177 35241 20211 35275
rect 21925 35241 21959 35275
rect 23673 35241 23707 35275
rect 23857 35241 23891 35275
rect 30849 35241 30883 35275
rect 33333 35241 33367 35275
rect 36277 35241 36311 35275
rect 37749 35241 37783 35275
rect 42901 35241 42935 35275
rect 34897 35173 34931 35207
rect 16129 35105 16163 35139
rect 23581 35105 23615 35139
rect 24593 35105 24627 35139
rect 25789 35105 25823 35139
rect 28733 35105 28767 35139
rect 35081 35105 35115 35139
rect 38301 35105 38335 35139
rect 40601 35105 40635 35139
rect 41521 35105 41555 35139
rect 14381 35037 14415 35071
rect 15117 35037 15151 35071
rect 15301 35037 15335 35071
rect 16405 35037 16439 35071
rect 16589 35037 16623 35071
rect 17969 35037 18003 35071
rect 18061 35037 18095 35071
rect 18245 35037 18279 35071
rect 18337 35037 18371 35071
rect 20729 35037 20763 35071
rect 21465 35037 21499 35071
rect 22109 35037 22143 35071
rect 22201 35037 22235 35071
rect 23673 35037 23707 35071
rect 25145 35037 25179 35071
rect 25329 35037 25363 35071
rect 25605 35037 25639 35071
rect 26663 35037 26697 35071
rect 27076 35037 27110 35071
rect 27169 35037 27203 35071
rect 28273 35037 28307 35071
rect 28365 35037 28399 35071
rect 29929 35037 29963 35071
rect 30113 35037 30147 35071
rect 30297 35037 30331 35071
rect 31125 35037 31159 35071
rect 32229 35037 32263 35071
rect 32413 35037 32447 35071
rect 32689 35037 32723 35071
rect 33517 35037 33551 35071
rect 33609 35037 33643 35071
rect 33793 35037 33827 35071
rect 33885 35037 33919 35071
rect 35173 35037 35207 35071
rect 35449 35037 35483 35071
rect 35541 35037 35575 35071
rect 37105 35037 37139 35071
rect 37198 35037 37232 35071
rect 37381 35037 37415 35071
rect 37611 35037 37645 35071
rect 38393 35037 38427 35071
rect 38945 35037 38979 35071
rect 40693 35037 40727 35071
rect 14473 34969 14507 35003
rect 14657 34969 14691 35003
rect 16497 34969 16531 35003
rect 21005 34969 21039 35003
rect 22477 34969 22511 35003
rect 22569 34969 22603 35003
rect 23397 34969 23431 35003
rect 26801 34969 26835 35003
rect 26893 34969 26927 35003
rect 28641 34969 28675 35003
rect 30021 34969 30055 35003
rect 36001 34969 36035 35003
rect 36185 34969 36219 35003
rect 37473 34969 37507 35003
rect 39497 34969 39531 35003
rect 41766 34969 41800 35003
rect 13737 34901 13771 34935
rect 14565 34901 14599 34935
rect 16865 34901 16899 34935
rect 17325 34901 17359 34935
rect 17877 34901 17911 34935
rect 18797 34901 18831 34935
rect 19717 34901 19751 34935
rect 26525 34901 26559 34935
rect 28089 34901 28123 34935
rect 29745 34901 29779 34935
rect 32597 34901 32631 34935
rect 41061 34901 41095 34935
rect 14013 34697 14047 34731
rect 16313 34697 16347 34731
rect 22109 34697 22143 34731
rect 29009 34697 29043 34731
rect 31769 34697 31803 34731
rect 41981 34697 42015 34731
rect 43269 34697 43303 34731
rect 24225 34629 24259 34663
rect 27353 34629 27387 34663
rect 33885 34629 33919 34663
rect 34621 34629 34655 34663
rect 35081 34629 35115 34663
rect 37841 34629 37875 34663
rect 40325 34629 40359 34663
rect 41429 34629 41463 34663
rect 13829 34561 13863 34595
rect 14473 34561 14507 34595
rect 14565 34561 14599 34595
rect 14749 34561 14783 34595
rect 15853 34561 15887 34595
rect 15945 34561 15979 34595
rect 16129 34561 16163 34595
rect 17141 34561 17175 34595
rect 17325 34561 17359 34595
rect 17417 34561 17451 34595
rect 17877 34561 17911 34595
rect 19533 34561 19567 34595
rect 20545 34561 20579 34595
rect 20913 34561 20947 34595
rect 22293 34561 22327 34595
rect 22385 34561 22419 34595
rect 24869 34561 24903 34595
rect 25421 34561 25455 34595
rect 25605 34561 25639 34595
rect 25697 34561 25731 34595
rect 25881 34561 25915 34595
rect 27997 34561 28031 34595
rect 28089 34561 28123 34595
rect 28365 34561 28399 34595
rect 29377 34561 29411 34595
rect 30573 34561 30607 34595
rect 30757 34561 30791 34595
rect 31401 34561 31435 34595
rect 32321 34561 32355 34595
rect 36461 34561 36495 34595
rect 36645 34561 36679 34595
rect 36829 34561 36863 34595
rect 37657 34561 37691 34595
rect 37749 34561 37783 34595
rect 38025 34561 38059 34595
rect 39598 34561 39632 34595
rect 40877 34561 40911 34595
rect 42809 34561 42843 34595
rect 13645 34493 13679 34527
rect 14933 34493 14967 34527
rect 16957 34493 16991 34527
rect 18153 34493 18187 34527
rect 21373 34493 21407 34527
rect 22661 34493 22695 34527
rect 23397 34493 23431 34527
rect 28457 34493 28491 34527
rect 29285 34493 29319 34527
rect 29837 34493 29871 34527
rect 30849 34493 30883 34527
rect 31493 34493 31527 34527
rect 33057 34493 33091 34527
rect 35909 34493 35943 34527
rect 36921 34493 36955 34527
rect 39865 34493 39899 34527
rect 42717 34493 42751 34527
rect 20545 34425 20579 34459
rect 30389 34425 30423 34459
rect 22569 34357 22603 34391
rect 26525 34357 26559 34391
rect 29285 34357 29319 34391
rect 31401 34357 31435 34391
rect 37473 34357 37507 34391
rect 38485 34357 38519 34391
rect 13737 34153 13771 34187
rect 14473 34153 14507 34187
rect 16865 34153 16899 34187
rect 17785 34153 17819 34187
rect 22201 34153 22235 34187
rect 24041 34153 24075 34187
rect 29101 34153 29135 34187
rect 29745 34153 29779 34187
rect 38945 34153 38979 34187
rect 14381 34085 14415 34119
rect 20545 34085 20579 34119
rect 25145 34085 25179 34119
rect 26985 34085 27019 34119
rect 27537 34085 27571 34119
rect 41429 34085 41463 34119
rect 12725 34017 12759 34051
rect 22937 34017 22971 34051
rect 23857 34017 23891 34051
rect 37473 34017 37507 34051
rect 13185 33949 13219 33983
rect 13277 33949 13311 33983
rect 13461 33949 13495 33983
rect 13553 33949 13587 33983
rect 14289 33949 14323 33983
rect 14565 33949 14599 33983
rect 14657 33949 14691 33983
rect 16681 33949 16715 33983
rect 16773 33949 16807 33983
rect 17969 33949 18003 33983
rect 18061 33949 18095 33983
rect 18245 33949 18279 33983
rect 18337 33949 18371 33983
rect 18889 33949 18923 33983
rect 21649 33949 21683 33983
rect 22017 33949 22051 33983
rect 23765 33949 23799 33983
rect 25324 33949 25358 33983
rect 25696 33949 25730 33983
rect 25789 33949 25823 33983
rect 26555 33949 26589 33983
rect 27077 33949 27111 33983
rect 27696 33949 27730 33983
rect 27905 33949 27939 33983
rect 28033 33949 28067 33983
rect 28174 33949 28208 33983
rect 29745 33949 29779 33983
rect 29929 33949 29963 33983
rect 31585 33949 31619 33983
rect 31769 33949 31803 33983
rect 32045 33949 32079 33983
rect 33052 33949 33086 33983
rect 33149 33949 33183 33983
rect 33424 33949 33458 33983
rect 33517 33949 33551 33983
rect 35909 33949 35943 33983
rect 36737 33949 36771 33983
rect 37197 33949 37231 33983
rect 38117 33949 38151 33983
rect 38485 33949 38519 33983
rect 39129 33949 39163 33983
rect 39405 33949 39439 33983
rect 40049 33949 40083 33983
rect 43269 33949 43303 33983
rect 15393 33881 15427 33915
rect 16037 33881 16071 33915
rect 16221 33881 16255 33915
rect 16957 33881 16991 33915
rect 20913 33881 20947 33915
rect 21833 33881 21867 33915
rect 21925 33881 21959 33915
rect 23397 33881 23431 33915
rect 23489 33881 23523 33915
rect 25421 33881 25455 33915
rect 25513 33881 25547 33915
rect 27813 33881 27847 33915
rect 28825 33881 28859 33915
rect 31401 33881 31435 33915
rect 33241 33881 33275 33915
rect 33977 33881 34011 33915
rect 35173 33881 35207 33915
rect 38209 33881 38243 33915
rect 38301 33881 38335 33915
rect 40294 33881 40328 33915
rect 43002 33881 43036 33915
rect 15853 33813 15887 33847
rect 19993 33813 20027 33847
rect 20453 33813 20487 33847
rect 24593 33813 24627 33847
rect 26433 33813 26467 33847
rect 26617 33813 26651 33847
rect 30481 33813 30515 33847
rect 32873 33813 32907 33847
rect 37933 33813 37967 33847
rect 39313 33813 39347 33847
rect 41889 33813 41923 33847
rect 13001 33609 13035 33643
rect 13645 33609 13679 33643
rect 15117 33609 15151 33643
rect 15577 33609 15611 33643
rect 16221 33609 16255 33643
rect 17969 33609 18003 33643
rect 24501 33609 24535 33643
rect 24961 33609 24995 33643
rect 28457 33609 28491 33643
rect 32413 33609 32447 33643
rect 38945 33609 38979 33643
rect 43269 33609 43303 33643
rect 17417 33541 17451 33575
rect 29745 33541 29779 33575
rect 30941 33541 30975 33575
rect 31125 33541 31159 33575
rect 37473 33541 37507 33575
rect 12265 33473 12299 33507
rect 12725 33473 12759 33507
rect 12909 33473 12943 33507
rect 14105 33473 14139 33507
rect 15761 33473 15795 33507
rect 17141 33473 17175 33507
rect 17877 33473 17911 33507
rect 18061 33473 18095 33507
rect 20361 33473 20395 33507
rect 21097 33473 21131 33507
rect 21281 33473 21315 33507
rect 22569 33473 22603 33507
rect 23397 33473 23431 33507
rect 23581 33473 23615 33507
rect 24317 33473 24351 33507
rect 24501 33473 24535 33507
rect 25145 33473 25179 33507
rect 25237 33473 25271 33507
rect 25329 33473 25363 33507
rect 25513 33473 25547 33507
rect 28181 33473 28215 33507
rect 29648 33473 29682 33507
rect 29837 33473 29871 33507
rect 30020 33473 30054 33507
rect 30113 33473 30147 33507
rect 30849 33473 30883 33507
rect 31585 33473 31619 33507
rect 32781 33473 32815 33507
rect 33241 33473 33275 33507
rect 34069 33473 34103 33507
rect 34529 33473 34563 33507
rect 35357 33473 35391 33507
rect 36001 33473 36035 33507
rect 36737 33473 36771 33507
rect 36921 33473 36955 33507
rect 38209 33473 38243 33507
rect 38669 33473 38703 33507
rect 39405 33473 39439 33507
rect 40049 33473 40083 33507
rect 40877 33473 40911 33507
rect 41705 33473 41739 33507
rect 42073 33473 42107 33507
rect 42809 33473 42843 33507
rect 13185 33405 13219 33439
rect 15853 33405 15887 33439
rect 17417 33405 17451 33439
rect 19165 33405 19199 33439
rect 19257 33405 19291 33439
rect 19625 33405 19659 33439
rect 20269 33405 20303 33439
rect 20453 33405 20487 33439
rect 20545 33405 20579 33439
rect 21189 33405 21223 33439
rect 22293 33405 22327 33439
rect 23857 33405 23891 33439
rect 26617 33405 26651 33439
rect 27813 33405 27847 33439
rect 27905 33405 27939 33439
rect 28273 33405 28307 33439
rect 32689 33405 32723 33439
rect 35265 33405 35299 33439
rect 36553 33405 36587 33439
rect 37841 33405 37875 33439
rect 38945 33405 38979 33439
rect 20085 33337 20119 33371
rect 22385 33337 22419 33371
rect 31677 33337 31711 33371
rect 35817 33337 35851 33371
rect 37933 33337 37967 33371
rect 41061 33337 41095 33371
rect 13829 33269 13863 33303
rect 17233 33269 17267 33303
rect 18981 33269 19015 33303
rect 22477 33269 22511 33303
rect 23765 33269 23799 33303
rect 25973 33269 26007 33303
rect 27261 33269 27295 33303
rect 29009 33269 29043 33303
rect 29469 33269 29503 33303
rect 31125 33269 31159 33303
rect 32781 33269 32815 33303
rect 33425 33269 33459 33303
rect 38071 33269 38105 33303
rect 38761 33269 38795 33303
rect 41521 33269 41555 33303
rect 41889 33269 41923 33303
rect 42717 33269 42751 33303
rect 12633 33065 12667 33099
rect 13093 33065 13127 33099
rect 14381 33065 14415 33099
rect 16497 33065 16531 33099
rect 16773 33065 16807 33099
rect 17877 33065 17911 33099
rect 19901 33065 19935 33099
rect 23489 33065 23523 33099
rect 23857 33065 23891 33099
rect 25881 33065 25915 33099
rect 27077 33065 27111 33099
rect 28825 33065 28859 33099
rect 30757 33065 30791 33099
rect 36553 33065 36587 33099
rect 36737 33065 36771 33099
rect 37381 33065 37415 33099
rect 37749 33065 37783 33099
rect 18705 32997 18739 33031
rect 21097 32997 21131 33031
rect 29745 32997 29779 33031
rect 31769 32997 31803 33031
rect 32965 32997 32999 33031
rect 34161 32997 34195 33031
rect 15853 32929 15887 32963
rect 16497 32929 16531 32963
rect 18429 32929 18463 32963
rect 20453 32929 20487 32963
rect 21649 32929 21683 32963
rect 23949 32929 23983 32963
rect 27629 32929 27663 32963
rect 34069 32929 34103 32963
rect 35633 32929 35667 32963
rect 37473 32929 37507 32963
rect 41337 32929 41371 32963
rect 41613 32929 41647 32963
rect 43361 32929 43395 32963
rect 12449 32861 12483 32895
rect 12633 32861 12667 32895
rect 13369 32861 13403 32895
rect 14749 32861 14783 32895
rect 16405 32861 16439 32895
rect 17509 32861 17543 32895
rect 20269 32861 20303 32895
rect 22477 32861 22511 32895
rect 22569 32861 22603 32895
rect 22661 32861 22695 32895
rect 22845 32861 22879 32895
rect 23673 32861 23707 32895
rect 25053 32861 25087 32895
rect 25421 32861 25455 32895
rect 26525 32861 26559 32895
rect 26893 32861 26927 32895
rect 27721 32861 27755 32895
rect 27905 32861 27939 32895
rect 29745 32861 29779 32895
rect 30021 32861 30055 32895
rect 30481 32861 30515 32895
rect 30573 32861 30607 32895
rect 30757 32861 30791 32895
rect 31953 32861 31987 32895
rect 32045 32861 32079 32895
rect 32321 32861 32355 32895
rect 32781 32861 32815 32895
rect 33977 32861 34011 32895
rect 34253 32861 34287 32895
rect 35541 32861 35575 32895
rect 36093 32861 36127 32895
rect 37381 32861 37415 32895
rect 39221 32861 39255 32895
rect 39405 32861 39439 32895
rect 40049 32861 40083 32895
rect 40233 32861 40267 32895
rect 40693 32861 40727 32895
rect 40877 32861 40911 32895
rect 13093 32793 13127 32827
rect 14565 32793 14599 32827
rect 17693 32793 17727 32827
rect 21465 32793 21499 32827
rect 25145 32793 25179 32827
rect 25237 32793 25271 32827
rect 26709 32793 26743 32827
rect 26801 32793 26835 32827
rect 28457 32793 28491 32827
rect 28641 32793 28675 32827
rect 32137 32793 32171 32827
rect 33793 32793 33827 32827
rect 36921 32793 36955 32827
rect 40141 32793 40175 32827
rect 13277 32725 13311 32759
rect 15209 32725 15243 32759
rect 15577 32725 15611 32759
rect 15669 32725 15703 32759
rect 18889 32725 18923 32759
rect 20361 32725 20395 32759
rect 21557 32725 21591 32759
rect 22293 32725 22327 32759
rect 24869 32725 24903 32759
rect 29929 32725 29963 32759
rect 31217 32725 31251 32759
rect 36721 32725 36755 32759
rect 38209 32725 38243 32759
rect 39313 32725 39347 32759
rect 40785 32725 40819 32759
rect 15945 32521 15979 32555
rect 16313 32521 16347 32555
rect 20177 32521 20211 32555
rect 20821 32521 20855 32555
rect 21465 32521 21499 32555
rect 22201 32521 22235 32555
rect 25789 32521 25823 32555
rect 27169 32521 27203 32555
rect 33615 32521 33649 32555
rect 34345 32521 34379 32555
rect 37473 32521 37507 32555
rect 43269 32521 43303 32555
rect 13093 32453 13127 32487
rect 18061 32453 18095 32487
rect 18705 32453 18739 32487
rect 24133 32453 24167 32487
rect 25145 32453 25179 32487
rect 26157 32453 26191 32487
rect 29193 32453 29227 32487
rect 30941 32453 30975 32487
rect 31125 32453 31159 32487
rect 32697 32453 32731 32487
rect 33517 32453 33551 32487
rect 41521 32453 41555 32487
rect 13277 32385 13311 32419
rect 13737 32385 13771 32419
rect 13921 32385 13955 32419
rect 14105 32385 14139 32419
rect 14197 32385 14231 32419
rect 14933 32385 14967 32419
rect 15117 32385 15151 32419
rect 17785 32385 17819 32419
rect 17877 32385 17911 32419
rect 18981 32385 19015 32419
rect 19073 32385 19107 32419
rect 19165 32385 19199 32419
rect 19349 32385 19383 32419
rect 21281 32385 21315 32419
rect 21465 32385 21499 32419
rect 22753 32385 22787 32419
rect 23949 32385 23983 32419
rect 24041 32385 24075 32419
rect 24317 32385 24351 32419
rect 24961 32385 24995 32419
rect 25053 32385 25087 32419
rect 25329 32385 25363 32419
rect 25973 32385 26007 32419
rect 26065 32385 26099 32419
rect 26341 32385 26375 32419
rect 28181 32385 28215 32419
rect 28365 32385 28399 32419
rect 28917 32385 28951 32419
rect 29010 32385 29044 32419
rect 29285 32385 29319 32419
rect 29423 32385 29457 32419
rect 30021 32385 30055 32419
rect 30205 32385 30239 32419
rect 30849 32385 30883 32419
rect 31585 32385 31619 32419
rect 31769 32385 31803 32419
rect 32573 32385 32607 32419
rect 32781 32385 32815 32419
rect 32965 32385 32999 32419
rect 33701 32385 33735 32419
rect 33793 32385 33827 32419
rect 35081 32385 35115 32419
rect 35173 32385 35207 32419
rect 35265 32385 35299 32419
rect 35449 32385 35483 32419
rect 36001 32385 36035 32419
rect 36093 32385 36127 32419
rect 36277 32385 36311 32419
rect 37749 32385 37783 32419
rect 37841 32385 37875 32419
rect 37933 32385 37967 32419
rect 38117 32385 38151 32419
rect 39129 32385 39163 32419
rect 39497 32385 39531 32419
rect 40233 32385 40267 32419
rect 40325 32385 40359 32419
rect 40601 32385 40635 32419
rect 41429 32385 41463 32419
rect 41613 32385 41647 32419
rect 42809 32385 42843 32419
rect 15761 32317 15795 32351
rect 15853 32317 15887 32351
rect 20361 32317 20395 32351
rect 20453 32317 20487 32351
rect 22477 32317 22511 32351
rect 28273 32317 28307 32351
rect 36737 32317 36771 32351
rect 38761 32317 38795 32351
rect 40141 32317 40175 32351
rect 40969 32317 41003 32351
rect 18061 32249 18095 32283
rect 24777 32249 24811 32283
rect 30205 32249 30239 32283
rect 34897 32249 34931 32283
rect 39497 32249 39531 32283
rect 12909 32181 12943 32215
rect 14933 32181 14967 32215
rect 17233 32181 17267 32215
rect 22569 32181 22603 32215
rect 23305 32181 23339 32215
rect 23765 32181 23799 32215
rect 29561 32181 29595 32215
rect 31125 32181 31159 32215
rect 31585 32181 31619 32215
rect 32413 32181 32447 32215
rect 42625 32181 42659 32215
rect 13093 31977 13127 32011
rect 13277 31977 13311 32011
rect 14289 31977 14323 32011
rect 15853 31977 15887 32011
rect 17049 31977 17083 32011
rect 26709 31977 26743 32011
rect 30205 31977 30239 32011
rect 31861 31977 31895 32011
rect 32321 31977 32355 32011
rect 34897 31977 34931 32011
rect 36553 31977 36587 32011
rect 37657 31977 37691 32011
rect 38209 31977 38243 32011
rect 15393 31909 15427 31943
rect 17601 31909 17635 31943
rect 19441 31909 19475 31943
rect 28733 31909 28767 31943
rect 32965 31909 32999 31943
rect 34161 31909 34195 31943
rect 12541 31841 12575 31875
rect 16497 31841 16531 31875
rect 18245 31841 18279 31875
rect 19993 31841 20027 31875
rect 20729 31841 20763 31875
rect 23121 31841 23155 31875
rect 32137 31841 32171 31875
rect 34253 31841 34287 31875
rect 42901 31841 42935 31875
rect 43177 31841 43211 31875
rect 12449 31773 12483 31807
rect 12633 31773 12667 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 15025 31773 15059 31807
rect 15209 31773 15243 31807
rect 16221 31773 16255 31807
rect 18061 31773 18095 31807
rect 18889 31773 18923 31807
rect 20821 31773 20855 31807
rect 21741 31773 21775 31807
rect 22017 31773 22051 31807
rect 23949 31773 23983 31807
rect 24777 31773 24811 31807
rect 24961 31773 24995 31807
rect 25145 31773 25179 31807
rect 25237 31773 25271 31807
rect 25881 31773 25915 31807
rect 26249 31773 26283 31807
rect 26893 31773 26927 31807
rect 26985 31773 27019 31807
rect 27077 31773 27111 31807
rect 27261 31773 27295 31807
rect 27813 31773 27847 31807
rect 28733 31773 28767 31807
rect 28917 31773 28951 31807
rect 29009 31773 29043 31807
rect 30021 31773 30055 31807
rect 31309 31773 31343 31807
rect 32045 31773 32079 31807
rect 32321 31773 32355 31807
rect 32781 31773 32815 31807
rect 33977 31773 34011 31807
rect 35265 31773 35299 31807
rect 35909 31773 35943 31807
rect 36093 31773 36127 31807
rect 36185 31773 36219 31807
rect 36277 31773 36311 31807
rect 37013 31773 37047 31807
rect 37841 31773 37875 31807
rect 38025 31773 38059 31807
rect 38301 31773 38335 31807
rect 39313 31773 39347 31807
rect 39497 31773 39531 31807
rect 40325 31773 40359 31807
rect 40476 31773 40510 31807
rect 40601 31773 40635 31807
rect 40693 31773 40727 31807
rect 13261 31705 13295 31739
rect 13461 31705 13495 31739
rect 21833 31705 21867 31739
rect 25973 31705 26007 31739
rect 26065 31705 26099 31739
rect 35081 31705 35115 31739
rect 16313 31637 16347 31671
rect 17969 31637 18003 31671
rect 19809 31637 19843 31671
rect 19901 31637 19935 31671
rect 22201 31637 22235 31671
rect 25697 31637 25731 31671
rect 31125 31637 31159 31671
rect 33793 31637 33827 31671
rect 39129 31637 39163 31671
rect 40141 31637 40175 31671
rect 41429 31637 41463 31671
rect 12081 31433 12115 31467
rect 13093 31433 13127 31467
rect 15301 31433 15335 31467
rect 15669 31433 15703 31467
rect 18245 31433 18279 31467
rect 41889 31433 41923 31467
rect 14289 31365 14323 31399
rect 14841 31365 14875 31399
rect 17233 31365 17267 31399
rect 20453 31365 20487 31399
rect 23029 31365 23063 31399
rect 24409 31365 24443 31399
rect 24501 31365 24535 31399
rect 25421 31365 25455 31399
rect 30205 31365 30239 31399
rect 30297 31365 30331 31399
rect 31217 31365 31251 31399
rect 33977 31365 34011 31399
rect 34805 31365 34839 31399
rect 38761 31365 38795 31399
rect 41061 31365 41095 31399
rect 12265 31297 12299 31331
rect 13185 31297 13219 31331
rect 13921 31297 13955 31331
rect 14105 31297 14139 31331
rect 15761 31297 15795 31331
rect 16957 31297 16991 31331
rect 17049 31297 17083 31331
rect 18242 31297 18276 31331
rect 19809 31297 19843 31331
rect 19901 31297 19935 31331
rect 20729 31297 20763 31331
rect 21373 31297 21407 31331
rect 21465 31297 21499 31331
rect 22201 31297 22235 31331
rect 22293 31297 22327 31331
rect 22569 31297 22603 31331
rect 23213 31297 23247 31331
rect 24317 31297 24351 31331
rect 24685 31297 24719 31331
rect 27721 31297 27755 31331
rect 28825 31297 28859 31331
rect 28917 31297 28951 31331
rect 29101 31297 29135 31331
rect 29193 31297 29227 31331
rect 30113 31297 30147 31331
rect 30481 31297 30515 31331
rect 30941 31297 30975 31331
rect 31033 31297 31067 31331
rect 31677 31297 31711 31331
rect 32505 31297 32539 31331
rect 32873 31297 32907 31331
rect 34345 31297 34379 31331
rect 34897 31297 34931 31331
rect 35081 31297 35115 31331
rect 35817 31297 35851 31331
rect 36645 31297 36679 31331
rect 36829 31297 36863 31331
rect 37473 31297 37507 31331
rect 38577 31297 38611 31331
rect 39221 31297 39255 31331
rect 39405 31297 39439 31331
rect 40417 31297 40451 31331
rect 41245 31297 41279 31331
rect 41337 31297 41371 31331
rect 42073 31297 42107 31331
rect 43085 31297 43119 31331
rect 13369 31229 13403 31263
rect 15853 31229 15887 31263
rect 18705 31229 18739 31263
rect 19625 31229 19659 31263
rect 19717 31229 19751 31263
rect 20453 31229 20487 31263
rect 21189 31229 21223 31263
rect 23397 31229 23431 31263
rect 23489 31229 23523 31263
rect 26157 31229 26191 31263
rect 27997 31229 28031 31263
rect 28641 31229 28675 31263
rect 35725 31229 35759 31263
rect 35909 31229 35943 31263
rect 36001 31229 36035 31263
rect 40601 31229 40635 31263
rect 18061 31161 18095 31195
rect 20637 31161 20671 31195
rect 22017 31161 22051 31195
rect 22477 31161 22511 31195
rect 37841 31161 37875 31195
rect 41061 31161 41095 31195
rect 12725 31093 12759 31127
rect 17233 31093 17267 31127
rect 18613 31093 18647 31127
rect 19441 31093 19475 31127
rect 21281 31093 21315 31127
rect 24133 31093 24167 31127
rect 29929 31093 29963 31127
rect 31217 31093 31251 31127
rect 32321 31093 32355 31127
rect 32781 31093 32815 31127
rect 33333 31093 33367 31127
rect 36185 31093 36219 31127
rect 36737 31093 36771 31127
rect 37933 31093 37967 31127
rect 38393 31093 38427 31127
rect 39313 31093 39347 31127
rect 40233 31093 40267 31127
rect 42625 31093 42659 31127
rect 42993 31093 43027 31127
rect 12725 30889 12759 30923
rect 13185 30889 13219 30923
rect 14381 30889 14415 30923
rect 18153 30889 18187 30923
rect 18613 30889 18647 30923
rect 20729 30889 20763 30923
rect 23673 30889 23707 30923
rect 31309 30889 31343 30923
rect 33057 30889 33091 30923
rect 37013 30889 37047 30923
rect 37565 30889 37599 30923
rect 38025 30889 38059 30923
rect 38209 30889 38243 30923
rect 39497 30889 39531 30923
rect 40141 30889 40175 30923
rect 21373 30821 21407 30855
rect 21925 30821 21959 30855
rect 22293 30821 22327 30855
rect 23121 30821 23155 30855
rect 32505 30821 32539 30855
rect 16129 30753 16163 30787
rect 24777 30753 24811 30787
rect 30757 30753 30791 30787
rect 33701 30753 33735 30787
rect 34161 30753 34195 30787
rect 42533 30753 42567 30787
rect 42809 30753 42843 30787
rect 12909 30685 12943 30719
rect 13001 30685 13035 30719
rect 13277 30685 13311 30719
rect 18889 30685 18923 30719
rect 19625 30685 19659 30719
rect 19717 30685 19751 30719
rect 19901 30685 19935 30719
rect 19993 30685 20027 30719
rect 21281 30685 21315 30719
rect 21465 30685 21499 30719
rect 22109 30685 22143 30719
rect 22385 30685 22419 30719
rect 23029 30685 23063 30719
rect 23213 30685 23247 30719
rect 24961 30685 24995 30719
rect 25421 30685 25455 30719
rect 25697 30685 25731 30719
rect 25881 30685 25915 30719
rect 27629 30685 27663 30719
rect 27905 30685 27939 30719
rect 27997 30685 28031 30719
rect 28273 30685 28307 30719
rect 28457 30685 28491 30719
rect 29929 30685 29963 30719
rect 30205 30685 30239 30719
rect 31401 30685 31435 30719
rect 32689 30685 32723 30719
rect 32781 30685 32815 30719
rect 33609 30685 33643 30719
rect 33977 30685 34011 30719
rect 34897 30685 34931 30719
rect 35449 30685 35483 30719
rect 35633 30685 35667 30719
rect 36277 30685 36311 30719
rect 36461 30685 36495 30719
rect 37197 30685 37231 30719
rect 37381 30685 37415 30719
rect 39313 30685 39347 30719
rect 39497 30685 39531 30719
rect 40049 30685 40083 30719
rect 40233 30685 40267 30719
rect 40693 30685 40727 30719
rect 40877 30685 40911 30719
rect 41981 30685 42015 30719
rect 18613 30617 18647 30651
rect 26709 30617 26743 30651
rect 33149 30617 33183 30651
rect 36093 30617 36127 30651
rect 36921 30617 36955 30651
rect 38393 30617 38427 30651
rect 40785 30617 40819 30651
rect 15485 30549 15519 30583
rect 15853 30549 15887 30583
rect 15945 30549 15979 30583
rect 17325 30549 17359 30583
rect 18797 30549 18831 30583
rect 19441 30549 19475 30583
rect 27261 30549 27295 30583
rect 29101 30549 29135 30583
rect 29745 30549 29779 30583
rect 30113 30549 30147 30583
rect 31953 30549 31987 30583
rect 38193 30549 38227 30583
rect 41705 30549 41739 30583
rect 18337 30345 18371 30379
rect 18245 30277 18279 30311
rect 19349 30277 19383 30311
rect 19441 30277 19475 30311
rect 20177 30277 20211 30311
rect 21097 30277 21131 30311
rect 23029 30277 23063 30311
rect 24961 30277 24995 30311
rect 28733 30277 28767 30311
rect 30297 30277 30331 30311
rect 32597 30277 32631 30311
rect 36829 30277 36863 30311
rect 38025 30277 38059 30311
rect 39865 30277 39899 30311
rect 40785 30277 40819 30311
rect 40969 30277 41003 30311
rect 12081 30209 12115 30243
rect 12265 30209 12299 30243
rect 16129 30209 16163 30243
rect 16313 30209 16347 30243
rect 19252 30209 19286 30243
rect 19569 30209 19603 30243
rect 19717 30209 19751 30243
rect 20361 30209 20395 30243
rect 20453 30209 20487 30243
rect 21281 30209 21315 30243
rect 22017 30209 22051 30243
rect 22201 30209 22235 30243
rect 22845 30209 22879 30243
rect 23949 30209 23983 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25421 30209 25455 30243
rect 25881 30209 25915 30243
rect 27445 30209 27479 30243
rect 28641 30209 28675 30243
rect 28825 30209 28859 30243
rect 29561 30209 29595 30243
rect 31401 30209 31435 30243
rect 31677 30209 31711 30243
rect 32873 30209 32907 30243
rect 34069 30209 34103 30243
rect 34529 30209 34563 30243
rect 35449 30209 35483 30243
rect 35725 30209 35759 30243
rect 35817 30209 35851 30243
rect 36737 30209 36771 30243
rect 36921 30209 36955 30243
rect 37473 30209 37507 30243
rect 37565 30209 37599 30243
rect 37749 30209 37783 30243
rect 37850 30209 37884 30243
rect 38945 30209 38979 30243
rect 39773 30209 39807 30243
rect 39957 30209 39991 30243
rect 41153 30209 41187 30243
rect 42073 30209 42107 30243
rect 43085 30209 43119 30243
rect 12173 30141 12207 30175
rect 12725 30141 12759 30175
rect 13829 30141 13863 30175
rect 14105 30141 14139 30175
rect 15485 30141 15519 30175
rect 18521 30141 18555 30175
rect 20177 30141 20211 30175
rect 21465 30141 21499 30175
rect 27353 30141 27387 30175
rect 31033 30141 31067 30175
rect 31217 30141 31251 30175
rect 32597 30141 32631 30175
rect 32781 30141 32815 30175
rect 33885 30141 33919 30175
rect 39037 30141 39071 30175
rect 42625 30141 42659 30175
rect 13093 30073 13127 30107
rect 16313 30073 16347 30107
rect 41889 30073 41923 30107
rect 13185 30005 13219 30039
rect 17877 30005 17911 30039
rect 19073 30005 19107 30039
rect 22017 30005 22051 30039
rect 22661 30005 22695 30039
rect 24409 30005 24443 30039
rect 26525 30005 26559 30039
rect 27721 30005 27755 30039
rect 29745 30005 29779 30039
rect 39037 30005 39071 30039
rect 39313 30005 39347 30039
rect 42809 30005 42843 30039
rect 11989 29801 12023 29835
rect 12633 29801 12667 29835
rect 13737 29801 13771 29835
rect 21925 29801 21959 29835
rect 22385 29801 22419 29835
rect 25697 29801 25731 29835
rect 27537 29801 27571 29835
rect 36093 29801 36127 29835
rect 37013 29801 37047 29835
rect 39221 29801 39255 29835
rect 41245 29801 41279 29835
rect 41429 29801 41463 29835
rect 18889 29733 18923 29767
rect 21465 29733 21499 29767
rect 27997 29733 28031 29767
rect 31125 29733 31159 29767
rect 35081 29733 35115 29767
rect 36461 29733 36495 29767
rect 38025 29733 38059 29767
rect 42901 29733 42935 29767
rect 12173 29665 12207 29699
rect 15485 29665 15519 29699
rect 16497 29665 16531 29699
rect 16681 29665 16715 29699
rect 19717 29665 19751 29699
rect 23305 29665 23339 29699
rect 23949 29665 23983 29699
rect 37197 29665 37231 29699
rect 38853 29665 38887 29699
rect 40049 29665 40083 29699
rect 40233 29665 40267 29699
rect 40325 29665 40359 29699
rect 40417 29665 40451 29699
rect 11437 29597 11471 29631
rect 11897 29597 11931 29631
rect 12817 29597 12851 29631
rect 13001 29597 13035 29631
rect 13093 29597 13127 29631
rect 13553 29597 13587 29631
rect 14289 29597 14323 29631
rect 14473 29597 14507 29631
rect 15393 29597 15427 29631
rect 17233 29597 17267 29631
rect 17417 29597 17451 29631
rect 17877 29597 17911 29631
rect 18153 29597 18187 29631
rect 18705 29597 18739 29631
rect 18889 29597 18923 29631
rect 19993 29597 20027 29631
rect 20085 29597 20119 29631
rect 20177 29597 20211 29631
rect 20361 29597 20395 29631
rect 21189 29597 21223 29631
rect 22109 29597 22143 29631
rect 22201 29597 22235 29631
rect 22477 29597 22511 29631
rect 23121 29597 23155 29631
rect 23397 29597 23431 29631
rect 23857 29597 23891 29631
rect 24041 29597 24075 29631
rect 24777 29597 24811 29631
rect 24869 29597 24903 29631
rect 25145 29597 25179 29631
rect 26157 29597 26191 29631
rect 29101 29597 29135 29631
rect 29745 29597 29779 29631
rect 30001 29597 30035 29631
rect 32689 29597 32723 29631
rect 32873 29597 32907 29631
rect 33333 29597 33367 29631
rect 33517 29597 33551 29631
rect 33977 29597 34011 29631
rect 34161 29597 34195 29631
rect 34897 29597 34931 29631
rect 36277 29597 36311 29631
rect 36553 29597 36587 29631
rect 37289 29597 37323 29631
rect 38025 29597 38059 29631
rect 38209 29597 38243 29631
rect 38945 29597 38979 29631
rect 39313 29597 39347 29631
rect 40509 29597 40543 29631
rect 41521 29597 41555 29631
rect 41613 29597 41647 29631
rect 12173 29529 12207 29563
rect 21281 29529 21315 29563
rect 21465 29529 21499 29563
rect 22937 29529 22971 29563
rect 24961 29529 24995 29563
rect 26424 29529 26458 29563
rect 31677 29529 31711 29563
rect 32505 29529 32539 29563
rect 37013 29529 37047 29563
rect 42257 29529 42291 29563
rect 42441 29529 42475 29563
rect 43085 29529 43119 29563
rect 43269 29529 43303 29563
rect 14289 29461 14323 29495
rect 16037 29461 16071 29495
rect 16405 29461 16439 29495
rect 17325 29461 17359 29495
rect 17975 29461 18009 29495
rect 18061 29461 18095 29495
rect 24593 29461 24627 29495
rect 28549 29461 28583 29495
rect 31953 29461 31987 29495
rect 33425 29461 33459 29495
rect 34345 29461 34379 29495
rect 37473 29461 37507 29495
rect 39497 29461 39531 29495
rect 42073 29461 42107 29495
rect 13553 29257 13587 29291
rect 16957 29257 16991 29291
rect 19533 29257 19567 29291
rect 20085 29257 20119 29291
rect 20545 29257 20579 29291
rect 21465 29257 21499 29291
rect 22845 29257 22879 29291
rect 23213 29257 23247 29291
rect 25145 29257 25179 29291
rect 26617 29257 26651 29291
rect 28549 29257 28583 29291
rect 29377 29257 29411 29291
rect 30021 29257 30055 29291
rect 31217 29257 31251 29291
rect 32321 29257 32355 29291
rect 34805 29257 34839 29291
rect 36645 29257 36679 29291
rect 37565 29257 37599 29291
rect 40233 29257 40267 29291
rect 42625 29257 42659 29291
rect 13921 29189 13955 29223
rect 15025 29189 15059 29223
rect 23857 29189 23891 29223
rect 27414 29189 27448 29223
rect 30205 29189 30239 29223
rect 35265 29189 35299 29223
rect 38485 29189 38519 29223
rect 12633 29121 12667 29155
rect 12909 29121 12943 29155
rect 13001 29121 13035 29155
rect 13737 29121 13771 29155
rect 14841 29121 14875 29155
rect 15117 29121 15151 29155
rect 15669 29121 15703 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 16221 29121 16255 29155
rect 17141 29121 17175 29155
rect 17969 29121 18003 29155
rect 18061 29121 18095 29155
rect 18245 29121 18279 29155
rect 18981 29121 19015 29155
rect 19441 29121 19475 29155
rect 19625 29121 19659 29155
rect 20453 29121 20487 29155
rect 22293 29121 22327 29155
rect 23029 29121 23063 29155
rect 23305 29121 23339 29155
rect 24317 29121 24351 29155
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 25053 29121 25087 29155
rect 25421 29121 25455 29155
rect 26433 29121 26467 29155
rect 29561 29121 29595 29155
rect 30389 29121 30423 29155
rect 30849 29121 30883 29155
rect 31033 29121 31067 29155
rect 32505 29121 32539 29155
rect 32689 29121 32723 29155
rect 33333 29121 33367 29155
rect 34161 29121 34195 29155
rect 34345 29121 34379 29155
rect 34621 29121 34655 29155
rect 35541 29121 35575 29155
rect 36645 29121 36679 29155
rect 36921 29121 36955 29155
rect 37933 29121 37967 29155
rect 39313 29121 39347 29155
rect 39405 29121 39439 29155
rect 39497 29121 39531 29155
rect 39681 29121 39715 29155
rect 41613 29121 41647 29155
rect 42993 29121 43027 29155
rect 18366 29053 18400 29087
rect 20637 29053 20671 29087
rect 25605 29053 25639 29087
rect 27169 29053 27203 29087
rect 31769 29053 31803 29087
rect 35357 29053 35391 29087
rect 37841 29053 37875 29087
rect 39037 29053 39071 29087
rect 40969 29053 41003 29087
rect 41153 29053 41187 29087
rect 41705 29053 41739 29087
rect 42901 29053 42935 29087
rect 12725 28985 12759 29019
rect 14841 28985 14875 29019
rect 22109 28985 22143 29019
rect 24593 28985 24627 29019
rect 33517 28985 33551 29019
rect 34437 28985 34471 29019
rect 34529 28985 34563 29019
rect 35725 28985 35759 29019
rect 36737 28985 36771 29019
rect 13093 28917 13127 28951
rect 18429 28917 18463 28951
rect 35541 28917 35575 28951
rect 37933 28917 37967 28951
rect 41245 28917 41279 28951
rect 42809 28917 42843 28951
rect 15209 28713 15243 28747
rect 15761 28713 15795 28747
rect 16129 28713 16163 28747
rect 16773 28713 16807 28747
rect 19441 28713 19475 28747
rect 20269 28713 20303 28747
rect 30113 28713 30147 28747
rect 34897 28713 34931 28747
rect 35357 28713 35391 28747
rect 35909 28713 35943 28747
rect 36737 28713 36771 28747
rect 38025 28713 38059 28747
rect 13185 28645 13219 28679
rect 13737 28645 13771 28679
rect 18429 28645 18463 28679
rect 21833 28645 21867 28679
rect 36277 28645 36311 28679
rect 41521 28645 41555 28679
rect 42533 28645 42567 28679
rect 16221 28577 16255 28611
rect 17509 28577 17543 28611
rect 17693 28577 17727 28611
rect 17785 28577 17819 28611
rect 18797 28577 18831 28611
rect 20913 28577 20947 28611
rect 26065 28577 26099 28611
rect 26709 28577 26743 28611
rect 27261 28577 27295 28611
rect 28917 28577 28951 28611
rect 30757 28577 30791 28611
rect 32597 28577 32631 28611
rect 34989 28577 35023 28611
rect 38209 28577 38243 28611
rect 41429 28577 41463 28611
rect 42809 28577 42843 28611
rect 13277 28509 13311 28543
rect 13461 28509 13495 28543
rect 15301 28509 15335 28543
rect 15945 28509 15979 28543
rect 16865 28509 16899 28543
rect 17601 28509 17635 28543
rect 19809 28509 19843 28543
rect 20453 28509 20487 28543
rect 20545 28509 20579 28543
rect 21833 28509 21867 28543
rect 22109 28509 22143 28543
rect 22845 28509 22879 28543
rect 23489 28509 23523 28543
rect 26249 28509 26283 28543
rect 26985 28509 27019 28543
rect 27102 28509 27136 28543
rect 30481 28509 30515 28543
rect 32413 28509 32447 28543
rect 33057 28509 33091 28543
rect 33885 28509 33919 28543
rect 33977 28509 34011 28543
rect 34161 28509 34195 28543
rect 35173 28509 35207 28543
rect 35817 28509 35851 28543
rect 36001 28509 36035 28543
rect 36093 28509 36127 28543
rect 37013 28509 37047 28543
rect 37197 28509 37231 28543
rect 38301 28509 38335 28543
rect 40417 28509 40451 28543
rect 40601 28509 40635 28543
rect 41889 28509 41923 28543
rect 41981 28509 42015 28543
rect 42901 28509 42935 28543
rect 12909 28441 12943 28475
rect 19625 28441 19659 28475
rect 22017 28441 22051 28475
rect 23397 28441 23431 28475
rect 25605 28441 25639 28475
rect 31493 28441 31527 28475
rect 31677 28441 31711 28475
rect 34345 28441 34379 28475
rect 34897 28441 34931 28475
rect 38025 28441 38059 28475
rect 39037 28441 39071 28475
rect 39405 28441 39439 28475
rect 40509 28441 40543 28475
rect 14841 28373 14875 28407
rect 17325 28373 17359 28407
rect 18337 28373 18371 28407
rect 22661 28373 22695 28407
rect 24041 28373 24075 28407
rect 25053 28373 25087 28407
rect 27905 28373 27939 28407
rect 28365 28373 28399 28407
rect 28733 28373 28767 28407
rect 28825 28373 28859 28407
rect 30573 28373 30607 28407
rect 31309 28373 31343 28407
rect 36921 28373 36955 28407
rect 38485 28373 38519 28407
rect 41153 28373 41187 28407
rect 14841 28169 14875 28203
rect 16957 28169 16991 28203
rect 18613 28169 18647 28203
rect 22293 28169 22327 28203
rect 23397 28169 23431 28203
rect 25605 28169 25639 28203
rect 27169 28169 27203 28203
rect 27629 28169 27663 28203
rect 28917 28169 28951 28203
rect 32689 28169 32723 28203
rect 32965 28169 32999 28203
rect 33425 28169 33459 28203
rect 35909 28169 35943 28203
rect 36369 28169 36403 28203
rect 41337 28169 41371 28203
rect 41981 28169 42015 28203
rect 20913 28101 20947 28135
rect 21373 28101 21407 28135
rect 27537 28101 27571 28135
rect 32597 28101 32631 28135
rect 12817 28033 12851 28067
rect 15209 28033 15243 28067
rect 17417 28033 17451 28067
rect 17601 28033 17635 28067
rect 18245 28033 18279 28067
rect 23581 28033 23615 28067
rect 24225 28033 24259 28067
rect 24492 28033 24526 28067
rect 28549 28033 28583 28067
rect 29377 28033 29411 28067
rect 29561 28033 29595 28067
rect 30573 28033 30607 28067
rect 30757 28033 30791 28067
rect 31217 28033 31251 28067
rect 32321 28033 32355 28067
rect 34161 28033 34195 28067
rect 34529 28033 34563 28067
rect 34713 28033 34747 28067
rect 35541 28033 35575 28067
rect 35725 28033 35759 28067
rect 38030 28033 38064 28067
rect 38209 28033 38243 28067
rect 39037 28033 39071 28067
rect 40141 28033 40175 28067
rect 43269 28033 43303 28067
rect 12909 27965 12943 27999
rect 15117 27965 15151 27999
rect 17509 27965 17543 27999
rect 18153 27965 18187 27999
rect 20453 27965 20487 27999
rect 23765 27965 23799 27999
rect 27721 27965 27755 27999
rect 28457 27965 28491 27999
rect 32806 27965 32840 27999
rect 34345 27965 34379 27999
rect 34437 27965 34471 27999
rect 39221 27965 39255 27999
rect 40969 27965 41003 27999
rect 41061 27965 41095 27999
rect 41521 27965 41555 27999
rect 20545 27897 20579 27931
rect 29469 27897 29503 27931
rect 30757 27897 30791 27931
rect 33977 27897 34011 27931
rect 37473 27897 37507 27931
rect 13185 27829 13219 27863
rect 22937 27829 22971 27863
rect 26065 27829 26099 27863
rect 30021 27829 30055 27863
rect 31401 27829 31435 27863
rect 35541 27829 35575 27863
rect 38025 27829 38059 27863
rect 38393 27829 38427 27863
rect 38853 27829 38887 27863
rect 40049 27829 40083 27863
rect 43177 27829 43211 27863
rect 26249 27625 26283 27659
rect 27353 27625 27387 27659
rect 29101 27625 29135 27659
rect 29745 27625 29779 27659
rect 35817 27625 35851 27659
rect 39405 27625 39439 27659
rect 41429 27625 41463 27659
rect 42349 27625 42383 27659
rect 20269 27557 20303 27591
rect 23857 27557 23891 27591
rect 25513 27557 25547 27591
rect 27721 27557 27755 27591
rect 31309 27557 31343 27591
rect 31585 27557 31619 27591
rect 32045 27557 32079 27591
rect 34345 27557 34379 27591
rect 37565 27557 37599 27591
rect 40233 27557 40267 27591
rect 43085 27557 43119 27591
rect 14289 27489 14323 27523
rect 21373 27489 21407 27523
rect 26433 27489 26467 27523
rect 30481 27489 30515 27523
rect 31401 27489 31435 27523
rect 33609 27489 33643 27523
rect 36369 27489 36403 27523
rect 38393 27489 38427 27523
rect 42441 27489 42475 27523
rect 14565 27421 14599 27455
rect 21629 27421 21663 27455
rect 23765 27421 23799 27455
rect 23949 27421 23983 27455
rect 25697 27421 25731 27455
rect 26525 27421 26559 27455
rect 27537 27421 27571 27455
rect 27813 27421 27847 27455
rect 29009 27421 29043 27455
rect 29193 27421 29227 27455
rect 30021 27421 30055 27455
rect 31217 27421 31251 27455
rect 32321 27421 32355 27455
rect 32413 27421 32447 27455
rect 33425 27421 33459 27455
rect 33517 27421 33551 27455
rect 34161 27421 34195 27455
rect 34345 27421 34379 27455
rect 34989 27421 35023 27455
rect 35173 27421 35207 27455
rect 35639 27421 35673 27455
rect 35817 27421 35851 27455
rect 36553 27421 36587 27455
rect 36645 27421 36679 27455
rect 37933 27421 37967 27455
rect 38577 27421 38611 27455
rect 38669 27421 38703 27455
rect 39313 27421 39347 27455
rect 39497 27421 39531 27455
rect 40417 27421 40451 27455
rect 40969 27421 41003 27455
rect 41337 27421 41371 27455
rect 41613 27421 41647 27455
rect 42533 27421 42567 27455
rect 42993 27421 43027 27455
rect 43177 27421 43211 27455
rect 15945 27353 15979 27387
rect 24593 27353 24627 27387
rect 24961 27353 24995 27387
rect 26249 27353 26283 27387
rect 29745 27353 29779 27387
rect 31585 27353 31619 27387
rect 32597 27353 32631 27387
rect 37749 27353 37783 27387
rect 20729 27285 20763 27319
rect 22753 27285 22787 27319
rect 26709 27285 26743 27319
rect 28273 27285 28307 27319
rect 29929 27285 29963 27319
rect 32229 27285 32263 27319
rect 35081 27285 35115 27319
rect 36369 27285 36403 27319
rect 38393 27285 38427 27319
rect 41153 27285 41187 27319
rect 42165 27285 42199 27319
rect 16221 27081 16255 27115
rect 22017 27081 22051 27115
rect 24685 27081 24719 27115
rect 25697 27081 25731 27115
rect 26065 27081 26099 27115
rect 29193 27081 29227 27115
rect 30389 27081 30423 27115
rect 31769 27081 31803 27115
rect 32413 27081 32447 27115
rect 35449 27081 35483 27115
rect 36185 27081 36219 27115
rect 42625 27081 42659 27115
rect 17132 27013 17166 27047
rect 20453 27013 20487 27047
rect 23029 27013 23063 27047
rect 29699 27013 29733 27047
rect 31401 27013 31435 27047
rect 39405 27013 39439 27047
rect 39497 27013 39531 27047
rect 41981 27013 42015 27047
rect 16865 26945 16899 26979
rect 19533 26945 19567 26979
rect 22201 26945 22235 26979
rect 23489 26945 23523 26979
rect 23673 26945 23707 26979
rect 24869 26945 24903 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 28089 26945 28123 26979
rect 28181 26945 28215 26979
rect 28365 26945 28399 26979
rect 28457 26945 28491 26979
rect 29377 26945 29411 26979
rect 29469 26945 29503 26979
rect 29561 26945 29595 26979
rect 30297 26945 30331 26979
rect 31585 26945 31619 26979
rect 32321 26945 32355 26979
rect 32505 26945 32539 26979
rect 33149 26945 33183 26979
rect 33333 26945 33367 26979
rect 34253 26945 34287 26979
rect 35081 26945 35115 26979
rect 35173 26945 35207 26979
rect 36369 26945 36403 26979
rect 36737 26945 36771 26979
rect 37749 26945 37783 26979
rect 37841 26945 37875 26979
rect 37933 26945 37967 26979
rect 38117 26945 38151 26979
rect 38945 26945 38979 26979
rect 39773 26945 39807 26979
rect 41153 26945 41187 26979
rect 43085 26945 43119 26979
rect 14657 26877 14691 26911
rect 14933 26877 14967 26911
rect 19625 26877 19659 26911
rect 21373 26877 21407 26911
rect 22385 26877 22419 26911
rect 25053 26877 25087 26911
rect 26157 26877 26191 26911
rect 26249 26877 26283 26911
rect 29837 26877 29871 26911
rect 34069 26877 34103 26911
rect 34161 26877 34195 26911
rect 36829 26877 36863 26911
rect 38853 26877 38887 26911
rect 39865 26877 39899 26911
rect 41061 26877 41095 26911
rect 41613 26877 41647 26911
rect 33885 26809 33919 26843
rect 18245 26741 18279 26775
rect 19809 26741 19843 26775
rect 23489 26741 23523 26775
rect 23857 26741 23891 26775
rect 27169 26741 27203 26775
rect 27905 26741 27939 26775
rect 33149 26741 33183 26775
rect 34069 26741 34103 26775
rect 35081 26741 35115 26775
rect 36369 26741 36403 26775
rect 37473 26741 37507 26775
rect 38577 26741 38611 26775
rect 38853 26741 38887 26775
rect 40049 26741 40083 26775
rect 41521 26741 41555 26775
rect 42809 26741 42843 26775
rect 21649 26537 21683 26571
rect 25789 26537 25823 26571
rect 26709 26537 26743 26571
rect 29837 26537 29871 26571
rect 30573 26537 30607 26571
rect 32781 26537 32815 26571
rect 35725 26537 35759 26571
rect 36829 26537 36863 26571
rect 41337 26537 41371 26571
rect 15669 26469 15703 26503
rect 20085 26469 20119 26503
rect 21005 26469 21039 26503
rect 26249 26469 26283 26503
rect 27905 26469 27939 26503
rect 19809 26401 19843 26435
rect 22569 26401 22603 26435
rect 23581 26401 23615 26435
rect 25973 26401 26007 26435
rect 27169 26401 27203 26435
rect 27353 26401 27387 26435
rect 28457 26401 28491 26435
rect 31125 26401 31159 26435
rect 36921 26401 36955 26435
rect 38945 26401 38979 26435
rect 39313 26401 39347 26435
rect 39405 26401 39439 26435
rect 40049 26401 40083 26435
rect 14289 26333 14323 26367
rect 17417 26333 17451 26367
rect 19717 26333 19751 26367
rect 22477 26333 22511 26367
rect 22661 26333 22695 26367
rect 23673 26333 23707 26367
rect 24961 26333 24995 26367
rect 25145 26333 25179 26367
rect 26065 26333 26099 26367
rect 27077 26333 27111 26367
rect 29929 26333 29963 26367
rect 31769 26333 31803 26367
rect 32965 26333 32999 26367
rect 33609 26333 33643 26367
rect 33793 26333 33827 26367
rect 33885 26333 33919 26367
rect 34897 26333 34931 26367
rect 36645 26333 36679 26367
rect 39037 26333 39071 26367
rect 40325 26333 40359 26367
rect 40417 26333 40451 26367
rect 40509 26333 40543 26367
rect 40693 26333 40727 26367
rect 41429 26333 41463 26367
rect 41797 26333 41831 26367
rect 42073 26333 42107 26367
rect 42901 26333 42935 26367
rect 14534 26265 14568 26299
rect 17684 26265 17718 26299
rect 21617 26265 21651 26299
rect 21833 26265 21867 26299
rect 25789 26265 25823 26299
rect 28273 26265 28307 26299
rect 29193 26265 29227 26299
rect 30941 26265 30975 26299
rect 33149 26265 33183 26299
rect 35081 26265 35115 26299
rect 35265 26265 35299 26299
rect 37381 26265 37415 26299
rect 37565 26265 37599 26299
rect 37749 26265 37783 26299
rect 18797 26197 18831 26231
rect 21465 26197 21499 26231
rect 24041 26197 24075 26231
rect 25053 26197 25087 26231
rect 28365 26197 28399 26231
rect 31033 26197 31067 26231
rect 36461 26197 36495 26231
rect 38209 26197 38243 26231
rect 38761 26197 38795 26231
rect 19625 25993 19659 26027
rect 20545 25993 20579 26027
rect 22017 25993 22051 26027
rect 27353 25993 27387 26027
rect 31033 25993 31067 26027
rect 32413 25993 32447 26027
rect 33333 25993 33367 26027
rect 34069 25993 34103 26027
rect 38301 25993 38335 26027
rect 40325 25993 40359 26027
rect 20453 25925 20487 25959
rect 24685 25925 24719 25959
rect 28365 25925 28399 25959
rect 30113 25925 30147 25959
rect 34621 25925 34655 25959
rect 38761 25925 38795 25959
rect 41061 25925 41095 25959
rect 41705 25925 41739 25959
rect 41910 25925 41944 25959
rect 13728 25857 13762 25891
rect 15853 25857 15887 25891
rect 18521 25857 18555 25891
rect 21281 25857 21315 25891
rect 21465 25857 21499 25891
rect 22477 25857 22511 25891
rect 23305 25857 23339 25891
rect 23581 25857 23615 25891
rect 24593 25857 24627 25891
rect 24869 25857 24903 25891
rect 25697 25857 25731 25891
rect 26157 25857 26191 25891
rect 27537 25857 27571 25891
rect 27629 25857 27663 25891
rect 27905 25857 27939 25891
rect 31401 25857 31435 25891
rect 32413 25857 32447 25891
rect 32505 25857 32539 25891
rect 33149 25857 33183 25891
rect 34161 25857 34195 25891
rect 35725 25857 35759 25891
rect 36185 25857 36219 25891
rect 37657 25857 37691 25891
rect 37749 25857 37783 25891
rect 38945 25857 38979 25891
rect 39129 25857 39163 25891
rect 39221 25857 39255 25891
rect 40509 25857 40543 25891
rect 42809 25857 42843 25891
rect 42901 25857 42935 25891
rect 13461 25789 13495 25823
rect 18613 25789 18647 25823
rect 18889 25789 18923 25823
rect 20729 25789 20763 25823
rect 23397 25789 23431 25823
rect 25053 25789 25087 25823
rect 25881 25789 25915 25823
rect 25973 25789 26007 25823
rect 26065 25789 26099 25823
rect 31493 25789 31527 25823
rect 31585 25789 31619 25823
rect 35817 25789 35851 25823
rect 36001 25789 36035 25823
rect 37473 25789 37507 25823
rect 41245 25789 41279 25823
rect 34621 25721 34655 25755
rect 36645 25721 36679 25755
rect 42073 25721 42107 25755
rect 14841 25653 14875 25687
rect 15669 25653 15703 25687
rect 20085 25653 20119 25687
rect 21465 25653 21499 25687
rect 22385 25653 22419 25687
rect 23765 25653 23799 25687
rect 26341 25653 26375 25687
rect 27813 25653 27847 25687
rect 33885 25653 33919 25687
rect 35449 25653 35483 25687
rect 35909 25653 35943 25687
rect 37749 25653 37783 25687
rect 39681 25653 39715 25687
rect 41889 25653 41923 25687
rect 42625 25653 42659 25687
rect 14289 25449 14323 25483
rect 19625 25449 19659 25483
rect 22937 25449 22971 25483
rect 23121 25449 23155 25483
rect 25237 25449 25271 25483
rect 27537 25449 27571 25483
rect 30389 25449 30423 25483
rect 31217 25449 31251 25483
rect 32321 25449 32355 25483
rect 34253 25449 34287 25483
rect 35725 25449 35759 25483
rect 42993 25449 43027 25483
rect 20177 25381 20211 25415
rect 31585 25381 31619 25415
rect 41337 25381 41371 25415
rect 15301 25313 15335 25347
rect 24961 25313 24995 25347
rect 26341 25313 26375 25347
rect 31493 25313 31527 25347
rect 36369 25313 36403 25347
rect 41245 25313 41279 25347
rect 42349 25313 42383 25347
rect 42834 25313 42868 25347
rect 14473 25245 14507 25279
rect 15568 25245 15602 25279
rect 17693 25245 17727 25279
rect 21097 25245 21131 25279
rect 22293 25245 22327 25279
rect 23673 25245 23707 25279
rect 23857 25245 23891 25279
rect 24593 25245 24627 25279
rect 25053 25245 25087 25279
rect 27721 25245 27755 25279
rect 27997 25245 28031 25279
rect 28181 25245 28215 25279
rect 28641 25245 28675 25279
rect 29745 25245 29779 25279
rect 30021 25245 30055 25279
rect 30205 25245 30239 25279
rect 31401 25245 31435 25279
rect 31677 25245 31711 25279
rect 32413 25245 32447 25279
rect 32873 25245 32907 25279
rect 33057 25245 33091 25279
rect 34069 25245 34103 25279
rect 34989 25245 35023 25279
rect 35173 25245 35207 25279
rect 35633 25245 35667 25279
rect 35817 25245 35851 25279
rect 37289 25245 37323 25279
rect 38209 25245 38243 25279
rect 38393 25245 38427 25279
rect 39129 25245 39163 25279
rect 39221 25245 39255 25279
rect 39405 25245 39439 25279
rect 39497 25245 39531 25279
rect 40049 25245 40083 25279
rect 40233 25245 40267 25279
rect 41705 25245 41739 25279
rect 41797 25245 41831 25279
rect 20913 25177 20947 25211
rect 21741 25177 21775 25211
rect 22753 25177 22787 25211
rect 24041 25177 24075 25211
rect 29883 25177 29917 25211
rect 30113 25177 30147 25211
rect 32965 25177 32999 25211
rect 33885 25177 33919 25211
rect 37105 25177 37139 25211
rect 38301 25177 38335 25211
rect 40877 25177 40911 25211
rect 16681 25109 16715 25143
rect 17509 25109 17543 25143
rect 20729 25109 20763 25143
rect 22953 25109 22987 25143
rect 25697 25109 25731 25143
rect 26893 25109 26927 25143
rect 28825 25109 28859 25143
rect 35081 25109 35115 25143
rect 37473 25109 37507 25143
rect 38945 25109 38979 25143
rect 40141 25109 40175 25143
rect 42625 25109 42659 25143
rect 42717 25109 42751 25143
rect 15577 24905 15611 24939
rect 19441 24905 19475 24939
rect 24777 24905 24811 24939
rect 31401 24905 31435 24939
rect 32321 24905 32355 24939
rect 38485 24905 38519 24939
rect 15945 24837 15979 24871
rect 17500 24837 17534 24871
rect 28926 24837 28960 24871
rect 36001 24837 36035 24871
rect 42763 24837 42797 24871
rect 42993 24837 43027 24871
rect 12909 24769 12943 24803
rect 13809 24769 13843 24803
rect 16037 24769 16071 24803
rect 19993 24769 20027 24803
rect 20177 24769 20211 24803
rect 20637 24769 20671 24803
rect 20913 24769 20947 24803
rect 22017 24769 22051 24803
rect 22109 24769 22143 24803
rect 23029 24769 23063 24803
rect 23213 24769 23247 24803
rect 23949 24769 23983 24803
rect 24961 24769 24995 24803
rect 25145 24769 25179 24803
rect 26525 24769 26559 24803
rect 27261 24769 27295 24803
rect 29193 24769 29227 24803
rect 29929 24769 29963 24803
rect 30021 24769 30055 24803
rect 30297 24769 30331 24803
rect 30941 24769 30975 24803
rect 32505 24769 32539 24803
rect 32781 24769 32815 24803
rect 32965 24769 32999 24803
rect 33701 24769 33735 24803
rect 33885 24769 33919 24803
rect 34529 24769 34563 24803
rect 34713 24769 34747 24803
rect 35725 24769 35759 24803
rect 36461 24769 36495 24803
rect 36645 24769 36679 24803
rect 36737 24769 36771 24803
rect 39313 24769 39347 24803
rect 40141 24769 40175 24803
rect 40325 24769 40359 24803
rect 40785 24769 40819 24803
rect 40877 24769 40911 24803
rect 41705 24769 41739 24803
rect 41981 24769 42015 24803
rect 42625 24769 42659 24803
rect 42901 24769 42935 24803
rect 43085 24769 43119 24803
rect 13553 24701 13587 24735
rect 16221 24701 16255 24735
rect 17233 24701 17267 24735
rect 23857 24701 23891 24735
rect 24225 24701 24259 24735
rect 24317 24701 24351 24735
rect 25053 24701 25087 24735
rect 25237 24701 25271 24735
rect 32689 24701 32723 24735
rect 36001 24701 36035 24735
rect 37473 24701 37507 24735
rect 39405 24701 39439 24735
rect 39497 24701 39531 24735
rect 39589 24701 39623 24735
rect 41797 24701 41831 24735
rect 13093 24633 13127 24667
rect 23121 24633 23155 24667
rect 27813 24633 27847 24667
rect 30849 24633 30883 24667
rect 32597 24633 32631 24667
rect 35173 24633 35207 24667
rect 37749 24633 37783 24667
rect 37933 24633 37967 24667
rect 41521 24633 41555 24667
rect 43269 24633 43303 24667
rect 14933 24565 14967 24599
rect 18613 24565 18647 24599
rect 20085 24565 20119 24599
rect 20729 24565 20763 24599
rect 21097 24565 21131 24599
rect 22017 24565 22051 24599
rect 22385 24565 22419 24599
rect 23673 24565 23707 24599
rect 25789 24565 25823 24599
rect 29745 24565 29779 24599
rect 30205 24565 30239 24599
rect 33885 24565 33919 24599
rect 34713 24565 34747 24599
rect 35817 24565 35851 24599
rect 36461 24565 36495 24599
rect 36921 24565 36955 24599
rect 39129 24565 39163 24599
rect 40325 24565 40359 24599
rect 41889 24565 41923 24599
rect 14289 24361 14323 24395
rect 17693 24361 17727 24395
rect 23765 24361 23799 24395
rect 24777 24361 24811 24395
rect 25697 24361 25731 24395
rect 28457 24361 28491 24395
rect 30941 24361 30975 24395
rect 32965 24361 32999 24395
rect 35081 24361 35115 24395
rect 36737 24361 36771 24395
rect 37381 24361 37415 24395
rect 38117 24361 38151 24395
rect 40049 24361 40083 24395
rect 40417 24361 40451 24395
rect 41245 24361 41279 24395
rect 42073 24361 42107 24395
rect 19809 24293 19843 24327
rect 23121 24293 23155 24327
rect 37197 24293 37231 24327
rect 14933 24225 14967 24259
rect 15485 24225 15519 24259
rect 18337 24225 18371 24259
rect 20269 24225 20303 24259
rect 21557 24225 21591 24259
rect 27813 24225 27847 24259
rect 29101 24225 29135 24259
rect 30297 24225 30331 24259
rect 31125 24225 31159 24259
rect 31585 24225 31619 24259
rect 33885 24225 33919 24259
rect 37565 24225 37599 24259
rect 14749 24157 14783 24191
rect 19533 24157 19567 24191
rect 20637 24157 20671 24191
rect 20729 24157 20763 24191
rect 21649 24157 21683 24191
rect 21741 24157 21775 24191
rect 21833 24157 21867 24191
rect 22385 24157 22419 24191
rect 22569 24157 22603 24191
rect 23765 24157 23799 24191
rect 23949 24157 23983 24191
rect 24041 24157 24075 24191
rect 24593 24157 24627 24191
rect 24961 24157 24995 24191
rect 25881 24157 25915 24191
rect 26617 24157 26651 24191
rect 26710 24157 26744 24191
rect 26893 24157 26927 24191
rect 27123 24157 27157 24191
rect 27721 24157 27755 24191
rect 27905 24157 27939 24191
rect 28825 24157 28859 24191
rect 30113 24157 30147 24191
rect 31217 24157 31251 24191
rect 32413 24157 32447 24191
rect 33609 24157 33643 24191
rect 33793 24157 33827 24191
rect 34069 24157 34103 24191
rect 34253 24157 34287 24191
rect 35081 24157 35115 24191
rect 35449 24157 35483 24191
rect 36369 24157 36403 24191
rect 36553 24157 36587 24191
rect 37381 24157 37415 24191
rect 37657 24157 37691 24191
rect 38117 24157 38151 24191
rect 38301 24157 38335 24191
rect 38945 24157 38979 24191
rect 39129 24157 39163 24191
rect 40049 24157 40083 24191
rect 40141 24157 40175 24191
rect 41429 24157 41463 24191
rect 41889 24157 41923 24191
rect 43269 24157 43303 24191
rect 18061 24089 18095 24123
rect 19809 24089 19843 24123
rect 26985 24089 27019 24123
rect 31493 24089 31527 24123
rect 14657 24021 14691 24055
rect 18153 24021 18187 24055
rect 19625 24021 19659 24055
rect 20913 24021 20947 24055
rect 21373 24021 21407 24055
rect 22477 24021 22511 24055
rect 25145 24021 25179 24055
rect 27261 24021 27295 24055
rect 28917 24021 28951 24055
rect 29745 24021 29779 24055
rect 30205 24021 30239 24055
rect 32229 24021 32263 24055
rect 35265 24021 35299 24055
rect 38485 24021 38519 24055
rect 39037 24021 39071 24055
rect 43177 24021 43211 24055
rect 14105 23817 14139 23851
rect 14565 23817 14599 23851
rect 23673 23817 23707 23851
rect 26617 23817 26651 23851
rect 29101 23817 29135 23851
rect 30297 23817 30331 23851
rect 30757 23817 30791 23851
rect 34345 23817 34379 23851
rect 35265 23817 35299 23851
rect 39681 23817 39715 23851
rect 40693 23817 40727 23851
rect 42993 23817 43027 23851
rect 21005 23749 21039 23783
rect 22293 23749 22327 23783
rect 22385 23749 22419 23783
rect 25482 23749 25516 23783
rect 31769 23749 31803 23783
rect 32321 23749 32355 23783
rect 33609 23749 33643 23783
rect 34897 23749 34931 23783
rect 39037 23749 39071 23783
rect 40785 23749 40819 23783
rect 14473 23681 14507 23715
rect 15301 23681 15335 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 15669 23681 15703 23715
rect 17693 23681 17727 23715
rect 18521 23681 18555 23715
rect 18889 23681 18923 23715
rect 18981 23681 19015 23715
rect 20637 23681 20671 23715
rect 20729 23681 20763 23715
rect 22201 23681 22235 23715
rect 22569 23681 22603 23715
rect 23029 23681 23063 23715
rect 24593 23681 24627 23715
rect 27445 23681 27479 23715
rect 27905 23681 27939 23715
rect 28733 23681 28767 23715
rect 29929 23681 29963 23715
rect 30941 23681 30975 23715
rect 31217 23681 31251 23715
rect 32597 23681 32631 23715
rect 33517 23681 33551 23715
rect 33793 23681 33827 23715
rect 34253 23681 34287 23715
rect 34437 23681 34471 23715
rect 35081 23681 35115 23715
rect 35909 23681 35943 23715
rect 36369 23681 36403 23715
rect 37657 23681 37691 23715
rect 38117 23681 38151 23715
rect 39313 23681 39347 23715
rect 39497 23681 39531 23715
rect 41337 23681 41371 23715
rect 41521 23681 41555 23715
rect 42809 23681 42843 23715
rect 14749 23613 14783 23647
rect 18613 23613 18647 23647
rect 21097 23613 21131 23647
rect 25237 23613 25271 23647
rect 27629 23613 27663 23647
rect 28825 23613 28859 23647
rect 29745 23613 29779 23647
rect 29837 23613 29871 23647
rect 31125 23613 31159 23647
rect 32505 23613 32539 23647
rect 36093 23613 36127 23647
rect 36185 23613 36219 23647
rect 36921 23613 36955 23647
rect 37749 23613 37783 23647
rect 13645 23545 13679 23579
rect 17969 23545 18003 23579
rect 24777 23545 24811 23579
rect 33793 23545 33827 23579
rect 36001 23545 36035 23579
rect 15945 23477 15979 23511
rect 20453 23477 20487 23511
rect 22017 23477 22051 23511
rect 23213 23477 23247 23511
rect 27169 23477 27203 23511
rect 27537 23477 27571 23511
rect 27721 23477 27755 23511
rect 28733 23477 28767 23511
rect 31217 23477 31251 23511
rect 32413 23477 32447 23511
rect 35725 23477 35759 23511
rect 37473 23477 37507 23511
rect 37657 23477 37691 23511
rect 39129 23477 39163 23511
rect 15761 23273 15795 23307
rect 21925 23273 21959 23307
rect 22385 23273 22419 23307
rect 25973 23273 26007 23307
rect 31125 23273 31159 23307
rect 33149 23273 33183 23307
rect 33977 23273 34011 23307
rect 35357 23273 35391 23307
rect 36829 23273 36863 23307
rect 38301 23273 38335 23307
rect 39313 23273 39347 23307
rect 40233 23273 40267 23307
rect 41705 23273 41739 23307
rect 41889 23273 41923 23307
rect 42809 23273 42843 23307
rect 14289 23205 14323 23239
rect 16589 23205 16623 23239
rect 19993 23205 20027 23239
rect 32597 23205 32631 23239
rect 37289 23205 37323 23239
rect 40509 23205 40543 23239
rect 17049 23137 17083 23171
rect 17877 23137 17911 23171
rect 19717 23137 19751 23171
rect 20545 23137 20579 23171
rect 23765 23137 23799 23171
rect 24777 23137 24811 23171
rect 25237 23137 25271 23171
rect 26617 23137 26651 23171
rect 27537 23137 27571 23171
rect 37013 23137 37047 23171
rect 38117 23137 38151 23171
rect 40141 23137 40175 23171
rect 42073 23137 42107 23171
rect 13645 23069 13679 23103
rect 15117 23069 15151 23103
rect 15301 23069 15335 23103
rect 15393 23069 15427 23103
rect 15485 23069 15519 23103
rect 16313 23069 16347 23103
rect 17233 23069 17267 23103
rect 17601 23069 17635 23103
rect 18797 23069 18831 23103
rect 19625 23069 19659 23103
rect 20637 23069 20671 23103
rect 23498 23069 23532 23103
rect 24869 23069 24903 23103
rect 26341 23069 26375 23103
rect 27353 23069 27387 23103
rect 27629 23069 27663 23103
rect 28733 23069 28767 23103
rect 28825 23069 28859 23103
rect 29009 23069 29043 23103
rect 29745 23069 29779 23103
rect 34897 23069 34931 23103
rect 34989 23069 35023 23103
rect 35173 23069 35207 23103
rect 37105 23069 37139 23103
rect 37933 23069 37967 23103
rect 39221 23069 39255 23103
rect 39405 23069 39439 23103
rect 40325 23069 40359 23103
rect 41889 23069 41923 23103
rect 42809 23069 42843 23103
rect 42993 23069 43027 23103
rect 14473 23001 14507 23035
rect 14657 23001 14691 23035
rect 29193 23001 29227 23035
rect 29990 23001 30024 23035
rect 31953 23001 31987 23035
rect 33609 23001 33643 23035
rect 33793 23001 33827 23035
rect 36829 23001 36863 23035
rect 38393 23001 38427 23035
rect 40049 23001 40083 23035
rect 42349 23001 42383 23035
rect 13461 22933 13495 22967
rect 18613 22933 18647 22967
rect 21005 22933 21039 22967
rect 24593 22933 24627 22967
rect 26433 22933 26467 22967
rect 27169 22933 27203 22967
rect 28181 22933 28215 22967
rect 31677 22933 31711 22967
rect 35909 22933 35943 22967
rect 37749 22933 37783 22967
rect 40969 22933 41003 22967
rect 16037 22729 16071 22763
rect 17417 22729 17451 22763
rect 19349 22729 19383 22763
rect 21281 22729 21315 22763
rect 25053 22729 25087 22763
rect 28365 22729 28399 22763
rect 29377 22729 29411 22763
rect 29929 22729 29963 22763
rect 30389 22729 30423 22763
rect 30849 22729 30883 22763
rect 32505 22729 32539 22763
rect 32689 22729 32723 22763
rect 34713 22729 34747 22763
rect 36829 22729 36863 22763
rect 39129 22729 39163 22763
rect 43269 22729 43303 22763
rect 15945 22661 15979 22695
rect 22753 22661 22787 22695
rect 23581 22661 23615 22695
rect 32597 22661 32631 22695
rect 33333 22661 33367 22695
rect 42625 22661 42659 22695
rect 13544 22593 13578 22627
rect 18530 22593 18564 22627
rect 18797 22593 18831 22627
rect 22661 22593 22695 22627
rect 25237 22593 25271 22627
rect 25421 22593 25455 22627
rect 27261 22593 27295 22627
rect 30757 22593 30791 22627
rect 33425 22593 33459 22627
rect 33701 22593 33735 22627
rect 33885 22593 33919 22627
rect 34069 22593 34103 22627
rect 35633 22593 35667 22627
rect 35909 22593 35943 22627
rect 36093 22593 36127 22627
rect 36645 22593 36679 22627
rect 36829 22593 36863 22627
rect 37473 22593 37507 22627
rect 39037 22593 39071 22627
rect 39221 22593 39255 22627
rect 40877 22593 40911 22627
rect 41889 22593 41923 22627
rect 43085 22593 43119 22627
rect 13277 22525 13311 22559
rect 16221 22525 16255 22559
rect 22937 22525 22971 22559
rect 25973 22525 26007 22559
rect 31033 22525 31067 22559
rect 39681 22525 39715 22559
rect 42993 22525 43027 22559
rect 16865 22457 16899 22491
rect 20177 22457 20211 22491
rect 27813 22457 27847 22491
rect 32321 22457 32355 22491
rect 14657 22389 14691 22423
rect 15577 22389 15611 22423
rect 20729 22389 20763 22423
rect 22293 22389 22327 22423
rect 24133 22389 24167 22423
rect 26617 22389 26651 22423
rect 31585 22389 31619 22423
rect 32873 22389 32907 22423
rect 35771 22389 35805 22423
rect 36001 22389 36035 22423
rect 37565 22389 37599 22423
rect 38209 22389 38243 22423
rect 40233 22389 40267 22423
rect 41061 22389 41095 22423
rect 41981 22389 42015 22423
rect 42717 22389 42751 22423
rect 14289 22185 14323 22219
rect 19717 22185 19751 22219
rect 30849 22185 30883 22219
rect 35081 22185 35115 22219
rect 37657 22185 37691 22219
rect 39313 22185 39347 22219
rect 43223 22185 43257 22219
rect 16957 22117 16991 22151
rect 18613 22117 18647 22151
rect 29745 22117 29779 22151
rect 32045 22117 32079 22151
rect 13553 22049 13587 22083
rect 14749 22049 14783 22083
rect 14933 22049 14967 22083
rect 15577 22049 15611 22083
rect 18061 22049 18095 22083
rect 18153 22049 18187 22083
rect 20453 22049 20487 22083
rect 33885 22049 33919 22083
rect 36185 22049 36219 22083
rect 36553 22049 36587 22083
rect 41429 22049 41463 22083
rect 41797 22049 41831 22083
rect 12357 21981 12391 22015
rect 13461 21981 13495 22015
rect 14657 21981 14691 22015
rect 18245 21981 18279 22015
rect 21281 21981 21315 22015
rect 22109 21981 22143 22015
rect 23673 21981 23707 22015
rect 24593 21981 24627 22015
rect 26893 21981 26927 22015
rect 27353 21981 27387 22015
rect 29883 21981 29917 22015
rect 30297 21981 30331 22015
rect 30941 21981 30975 22015
rect 31769 21981 31803 22015
rect 32505 21981 32539 22015
rect 32965 21981 32999 22015
rect 33425 21981 33459 22015
rect 36369 21981 36403 22015
rect 36645 21981 36679 22015
rect 36737 21981 36771 22015
rect 36921 21981 36955 22015
rect 37657 21981 37691 22015
rect 37841 21981 37875 22015
rect 37933 21981 37967 22015
rect 38577 21981 38611 22015
rect 38761 21981 38795 22015
rect 40049 21981 40083 22015
rect 40233 21981 40267 22015
rect 40877 21981 40911 22015
rect 15822 21913 15856 21947
rect 19901 21913 19935 21947
rect 22845 21913 22879 21947
rect 24860 21913 24894 21947
rect 27620 21913 27654 21947
rect 30021 21913 30055 21947
rect 30113 21913 30147 21947
rect 34989 21913 35023 21947
rect 38669 21913 38703 21947
rect 12541 21845 12575 21879
rect 13001 21845 13035 21879
rect 13369 21845 13403 21879
rect 19533 21845 19567 21879
rect 19701 21845 19735 21879
rect 22293 21845 22327 21879
rect 25973 21845 26007 21879
rect 28733 21845 28767 21879
rect 38117 21845 38151 21879
rect 40141 21845 40175 21879
rect 40693 21845 40727 21879
rect 14749 21641 14783 21675
rect 15209 21641 15243 21675
rect 20821 21641 20855 21675
rect 23857 21641 23891 21675
rect 25697 21641 25731 21675
rect 25789 21641 25823 21675
rect 27169 21641 27203 21675
rect 29929 21641 29963 21675
rect 36001 21641 36035 21675
rect 38761 21641 38795 21675
rect 39865 21641 39899 21675
rect 42073 21641 42107 21675
rect 43361 21641 43395 21675
rect 19625 21573 19659 21607
rect 20913 21573 20947 21607
rect 22284 21573 22318 21607
rect 28816 21573 28850 21607
rect 30757 21573 30791 21607
rect 35725 21573 35759 21607
rect 37473 21573 37507 21607
rect 40601 21573 40635 21607
rect 42717 21573 42751 21607
rect 13369 21505 13403 21539
rect 13625 21505 13659 21539
rect 15393 21505 15427 21539
rect 15577 21505 15611 21539
rect 16313 21505 16347 21539
rect 17141 21505 17175 21539
rect 17877 21505 17911 21539
rect 17969 21505 18003 21539
rect 18153 21505 18187 21539
rect 18705 21505 18739 21539
rect 24869 21505 24903 21539
rect 26617 21505 26651 21539
rect 27537 21505 27571 21539
rect 30573 21505 30607 21539
rect 30849 21505 30883 21539
rect 31309 21505 31343 21539
rect 32689 21505 32723 21539
rect 32873 21505 32907 21539
rect 33793 21505 33827 21539
rect 34069 21505 34103 21539
rect 35449 21505 35483 21539
rect 35633 21505 35667 21539
rect 35817 21505 35851 21539
rect 37749 21505 37783 21539
rect 38393 21505 38427 21539
rect 39221 21505 39255 21539
rect 39681 21505 39715 21539
rect 40325 21505 40359 21539
rect 42809 21505 42843 21539
rect 21097 21437 21131 21471
rect 22017 21437 22051 21471
rect 25973 21437 26007 21471
rect 27629 21437 27663 21471
rect 27813 21437 27847 21471
rect 28549 21437 28583 21471
rect 32965 21437 32999 21471
rect 33149 21437 33183 21471
rect 33885 21437 33919 21471
rect 37565 21437 37599 21471
rect 38485 21437 38519 21471
rect 39497 21437 39531 21471
rect 20453 21369 20487 21403
rect 25329 21369 25363 21403
rect 31493 21369 31527 21403
rect 32413 21369 32447 21403
rect 32781 21369 32815 21403
rect 33977 21369 34011 21403
rect 37933 21369 37967 21403
rect 16129 21301 16163 21335
rect 17325 21301 17359 21335
rect 18981 21301 19015 21335
rect 19901 21301 19935 21335
rect 23397 21301 23431 21335
rect 24685 21301 24719 21335
rect 30665 21301 30699 21335
rect 33609 21301 33643 21335
rect 34805 21301 34839 21335
rect 36553 21301 36587 21335
rect 37473 21301 37507 21335
rect 38577 21301 38611 21335
rect 39681 21301 39715 21335
rect 15393 21097 15427 21131
rect 17785 21097 17819 21131
rect 22109 21097 22143 21131
rect 25973 21097 26007 21131
rect 26433 21097 26467 21131
rect 27721 21097 27755 21131
rect 28181 21097 28215 21131
rect 29101 21097 29135 21131
rect 32505 21097 32539 21131
rect 33609 21097 33643 21131
rect 34345 21097 34379 21131
rect 35265 21097 35299 21131
rect 35633 21097 35667 21131
rect 36185 21097 36219 21131
rect 36737 21097 36771 21131
rect 37565 21097 37599 21131
rect 40141 21097 40175 21131
rect 40693 21097 40727 21131
rect 38025 21029 38059 21063
rect 41153 21029 41187 21063
rect 18245 20961 18279 20995
rect 18429 20961 18463 20995
rect 22661 20961 22695 20995
rect 24593 20961 24627 20995
rect 27169 20961 27203 20995
rect 27261 20961 27295 20995
rect 28549 20961 28583 20995
rect 36829 20961 36863 20995
rect 37749 20961 37783 20995
rect 38945 20961 38979 20995
rect 39037 20961 39071 20995
rect 15209 20893 15243 20927
rect 15853 20893 15887 20927
rect 16120 20893 16154 20927
rect 21097 20893 21131 20927
rect 21281 20893 21315 20927
rect 22477 20893 22511 20927
rect 23489 20893 23523 20927
rect 23581 20893 23615 20927
rect 23765 20893 23799 20927
rect 24849 20893 24883 20927
rect 28365 20893 28399 20927
rect 28641 20893 28675 20927
rect 31493 20893 31527 20927
rect 32689 20893 32723 20927
rect 32781 20893 32815 20927
rect 32965 20893 32999 20927
rect 33057 20893 33091 20927
rect 35265 20893 35299 20927
rect 35449 20893 35483 20927
rect 36737 20893 36771 20927
rect 37841 20893 37875 20927
rect 38853 20893 38887 20927
rect 40325 20893 40359 20927
rect 40509 20893 40543 20927
rect 19901 20825 19935 20859
rect 20269 20825 20303 20859
rect 22569 20825 22603 20859
rect 23949 20825 23983 20859
rect 31226 20825 31260 20859
rect 37565 20825 37599 20859
rect 40049 20825 40083 20859
rect 42901 20825 42935 20859
rect 43269 20825 43303 20859
rect 14289 20757 14323 20791
rect 17233 20757 17267 20791
rect 18153 20757 18187 20791
rect 20913 20757 20947 20791
rect 27353 20757 27387 20791
rect 30113 20757 30147 20791
rect 37105 20757 37139 20791
rect 39221 20757 39255 20791
rect 41705 20757 41739 20791
rect 42257 20757 42291 20791
rect 14289 20553 14323 20587
rect 17141 20553 17175 20587
rect 20285 20553 20319 20587
rect 20453 20553 20487 20587
rect 22661 20553 22695 20587
rect 25421 20553 25455 20587
rect 27721 20553 27755 20587
rect 28181 20553 28215 20587
rect 30573 20553 30607 20587
rect 31769 20553 31803 20587
rect 34989 20553 35023 20587
rect 36001 20553 36035 20587
rect 39313 20553 39347 20587
rect 41981 20553 42015 20587
rect 14749 20485 14783 20519
rect 20085 20485 20119 20519
rect 25697 20485 25731 20519
rect 27261 20485 27295 20519
rect 28641 20485 28675 20519
rect 29101 20485 29135 20519
rect 13001 20417 13035 20451
rect 13645 20417 13679 20451
rect 14657 20417 14691 20451
rect 15485 20417 15519 20451
rect 15669 20417 15703 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 18153 20417 18187 20451
rect 19165 20417 19199 20451
rect 19533 20417 19567 20451
rect 21097 20417 21131 20451
rect 23489 20417 23523 20451
rect 25605 20417 25639 20451
rect 25789 20417 25823 20451
rect 25973 20417 26007 20451
rect 27445 20417 27479 20451
rect 27537 20417 27571 20451
rect 28365 20417 28399 20451
rect 29193 20417 29227 20451
rect 31125 20417 31159 20451
rect 32321 20417 32355 20451
rect 32505 20417 32539 20451
rect 32597 20417 32631 20451
rect 32689 20417 32723 20451
rect 33609 20417 33643 20451
rect 33876 20417 33910 20451
rect 35449 20417 35483 20451
rect 36921 20417 36955 20451
rect 37657 20417 37691 20451
rect 37841 20417 37875 20451
rect 38853 20417 38887 20451
rect 39129 20417 39163 20451
rect 40233 20417 40267 20451
rect 42993 20417 43027 20451
rect 14933 20349 14967 20383
rect 17877 20349 17911 20383
rect 18061 20349 18095 20383
rect 22753 20349 22787 20383
rect 22937 20349 22971 20383
rect 23673 20349 23707 20383
rect 28457 20349 28491 20383
rect 30849 20349 30883 20383
rect 35725 20349 35759 20383
rect 36645 20349 36679 20383
rect 38945 20349 38979 20383
rect 40509 20349 40543 20383
rect 36737 20281 36771 20315
rect 13185 20213 13219 20247
rect 13829 20213 13863 20247
rect 15853 20213 15887 20247
rect 20269 20213 20303 20247
rect 20913 20213 20947 20247
rect 22293 20213 22327 20247
rect 27353 20213 27387 20247
rect 28365 20213 28399 20247
rect 30113 20213 30147 20247
rect 31033 20213 31067 20247
rect 32873 20213 32907 20247
rect 35541 20213 35575 20247
rect 36829 20213 36863 20247
rect 37657 20213 37691 20247
rect 38025 20213 38059 20247
rect 38853 20213 38887 20247
rect 42901 20213 42935 20247
rect 13001 20009 13035 20043
rect 15669 20009 15703 20043
rect 16221 20009 16255 20043
rect 18797 20009 18831 20043
rect 19441 20009 19475 20043
rect 21649 20009 21683 20043
rect 22109 20009 22143 20043
rect 28273 20009 28307 20043
rect 28733 20009 28767 20043
rect 29837 20009 29871 20043
rect 30389 20009 30423 20043
rect 33149 20009 33183 20043
rect 33885 20009 33919 20043
rect 36461 20009 36495 20043
rect 38117 20009 38151 20043
rect 40233 20009 40267 20043
rect 43269 20009 43303 20043
rect 12541 19941 12575 19975
rect 37749 19941 37783 19975
rect 40693 19941 40727 19975
rect 13461 19873 13495 19907
rect 13645 19873 13679 19907
rect 16865 19873 16899 19907
rect 22753 19873 22787 19907
rect 23581 19873 23615 19907
rect 35449 19873 35483 19907
rect 41521 19873 41555 19907
rect 14289 19805 14323 19839
rect 17417 19805 17451 19839
rect 17673 19805 17707 19839
rect 19625 19805 19659 19839
rect 19717 19805 19751 19839
rect 20269 19805 20303 19839
rect 22477 19805 22511 19839
rect 23305 19805 23339 19839
rect 23397 19805 23431 19839
rect 24593 19805 24627 19839
rect 24777 19805 24811 19839
rect 27261 19805 27295 19839
rect 27721 19805 27755 19839
rect 28089 19805 28123 19839
rect 30573 19805 30607 19839
rect 30665 19805 30699 19839
rect 30941 19805 30975 19839
rect 31769 19805 31803 19839
rect 34069 19805 34103 19839
rect 35265 19805 35299 19839
rect 36461 19805 36495 19839
rect 36645 19805 36679 19839
rect 37657 19805 37691 19839
rect 37841 19805 37875 19839
rect 37933 19805 37967 19839
rect 38853 19805 38887 19839
rect 38945 19805 38979 19839
rect 39037 19805 39071 19839
rect 40049 19805 40083 19839
rect 14534 19737 14568 19771
rect 20536 19737 20570 19771
rect 24685 19737 24719 19771
rect 27905 19737 27939 19771
rect 27997 19737 28031 19771
rect 30757 19737 30791 19771
rect 32014 19737 32048 19771
rect 39221 19737 39255 19771
rect 41797 19737 41831 19771
rect 13369 19669 13403 19703
rect 16589 19669 16623 19703
rect 16681 19669 16715 19703
rect 22569 19669 22603 19703
rect 23581 19669 23615 19703
rect 27077 19669 27111 19703
rect 34897 19669 34931 19703
rect 35357 19669 35391 19703
rect 14749 19465 14783 19499
rect 15945 19465 15979 19499
rect 18337 19465 18371 19499
rect 19809 19465 19843 19499
rect 22293 19465 22327 19499
rect 22753 19465 22787 19499
rect 23673 19465 23707 19499
rect 24133 19465 24167 19499
rect 26249 19465 26283 19499
rect 27169 19465 27203 19499
rect 31769 19465 31803 19499
rect 35173 19465 35207 19499
rect 36001 19465 36035 19499
rect 37841 19465 37875 19499
rect 39306 19465 39340 19499
rect 41889 19465 41923 19499
rect 13614 19397 13648 19431
rect 22385 19397 22419 19431
rect 28282 19397 28316 19431
rect 29285 19397 29319 19431
rect 29377 19397 29411 19431
rect 30757 19397 30791 19431
rect 31401 19397 31435 19431
rect 31493 19397 31527 19431
rect 13369 19329 13403 19363
rect 15301 19329 15335 19363
rect 15485 19329 15519 19363
rect 15577 19329 15611 19363
rect 15669 19329 15703 19363
rect 17877 19329 17911 19363
rect 18337 19329 18371 19363
rect 19717 19329 19751 19363
rect 21465 19329 21499 19363
rect 23765 19329 23799 19363
rect 24869 19329 24903 19363
rect 25136 19329 25170 19363
rect 29193 19329 29227 19363
rect 29561 19329 29595 19363
rect 31217 19329 31251 19363
rect 31585 19329 31619 19363
rect 32413 19329 32447 19363
rect 33241 19329 33275 19363
rect 33793 19329 33827 19363
rect 34060 19329 34094 19363
rect 35817 19329 35851 19363
rect 37473 19329 37507 19363
rect 38485 19329 38519 19363
rect 38669 19329 38703 19363
rect 39129 19329 39163 19363
rect 39221 19329 39255 19363
rect 39405 19329 39439 19363
rect 39853 19329 39887 19363
rect 40049 19329 40083 19363
rect 40693 19329 40727 19363
rect 40785 19329 40819 19363
rect 40969 19329 41003 19363
rect 41981 19329 42015 19363
rect 19901 19261 19935 19295
rect 20729 19261 20763 19295
rect 22201 19261 22235 19295
rect 23581 19261 23615 19295
rect 28549 19261 28583 19295
rect 30113 19261 30147 19295
rect 36553 19261 36587 19295
rect 37565 19261 37599 19295
rect 42625 19261 42659 19295
rect 43177 19261 43211 19295
rect 38669 19193 38703 19227
rect 40049 19193 40083 19227
rect 19349 19125 19383 19159
rect 29009 19125 29043 19159
rect 37657 19125 37691 19159
rect 40969 19125 41003 19159
rect 15209 18921 15243 18955
rect 21281 18921 21315 18955
rect 22569 18921 22603 18955
rect 24593 18921 24627 18955
rect 31125 18921 31159 18955
rect 34253 18921 34287 18955
rect 34989 18921 35023 18955
rect 35633 18921 35667 18955
rect 36553 18921 36587 18955
rect 36921 18921 36955 18955
rect 37565 18921 37599 18955
rect 38025 18921 38059 18955
rect 39313 18921 39347 18955
rect 40233 18921 40267 18955
rect 43085 18921 43119 18955
rect 28089 18853 28123 18887
rect 18337 18785 18371 18819
rect 21833 18785 21867 18819
rect 41613 18785 41647 18819
rect 16865 18717 16899 18751
rect 17601 18717 17635 18751
rect 18245 18717 18279 18751
rect 19441 18717 19475 18751
rect 21649 18717 21683 18751
rect 21741 18717 21775 18751
rect 23121 18717 23155 18751
rect 23949 18717 23983 18751
rect 26709 18717 26743 18751
rect 26976 18717 27010 18751
rect 28641 18717 28675 18751
rect 28917 18717 28951 18751
rect 29009 18717 29043 18751
rect 29745 18717 29779 18751
rect 32790 18717 32824 18751
rect 33057 18717 33091 18751
rect 33701 18717 33735 18751
rect 33977 18717 34011 18751
rect 34069 18717 34103 18751
rect 35449 18717 35483 18751
rect 35633 18717 35667 18751
rect 36829 18717 36863 18751
rect 36921 18717 36955 18751
rect 37381 18717 37415 18751
rect 37565 18717 37599 18751
rect 40141 18717 40175 18751
rect 40325 18717 40359 18751
rect 42625 18717 42659 18751
rect 19686 18649 19720 18683
rect 28825 18649 28859 18683
rect 29990 18649 30024 18683
rect 33885 18649 33919 18683
rect 38761 18649 38795 18683
rect 40785 18649 40819 18683
rect 40969 18649 41003 18683
rect 17049 18581 17083 18615
rect 20821 18581 20855 18615
rect 29193 18581 29227 18615
rect 31677 18581 31711 18615
rect 38945 18581 38979 18615
rect 39037 18581 39071 18615
rect 39129 18581 39163 18615
rect 41153 18581 41187 18615
rect 42441 18581 42475 18615
rect 19901 18377 19935 18411
rect 22385 18377 22419 18411
rect 25053 18377 25087 18411
rect 32413 18377 32447 18411
rect 35081 18377 35115 18411
rect 36185 18377 36219 18411
rect 37749 18377 37783 18411
rect 38209 18377 38243 18411
rect 40049 18377 40083 18411
rect 42625 18377 42659 18411
rect 14657 18309 14691 18343
rect 23857 18309 23891 18343
rect 29009 18309 29043 18343
rect 31493 18309 31527 18343
rect 33057 18309 33091 18343
rect 37841 18309 37875 18343
rect 37927 18309 37961 18343
rect 39865 18309 39899 18343
rect 40868 18309 40902 18343
rect 14841 18241 14875 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 17417 18241 17451 18275
rect 17877 18241 17911 18275
rect 18245 18241 18279 18275
rect 18613 18241 18647 18275
rect 18705 18241 18739 18275
rect 19809 18241 19843 18275
rect 20085 18241 20119 18275
rect 20729 18241 20763 18275
rect 20913 18241 20947 18275
rect 21005 18241 21039 18275
rect 22753 18241 22787 18275
rect 23581 18241 23615 18275
rect 26177 18241 26211 18275
rect 29920 18241 29954 18275
rect 32321 18241 32355 18275
rect 32505 18241 32539 18275
rect 34437 18241 34471 18275
rect 34621 18241 34655 18275
rect 37473 18241 37507 18275
rect 38669 18241 38703 18275
rect 38761 18241 38795 18275
rect 38945 18241 38979 18275
rect 39037 18241 39071 18275
rect 39681 18241 39715 18275
rect 42993 18241 43027 18275
rect 16129 18173 16163 18207
rect 18153 18173 18187 18207
rect 22845 18173 22879 18207
rect 22937 18173 22971 18207
rect 26433 18173 26467 18207
rect 28181 18173 28215 18207
rect 29653 18173 29687 18207
rect 33793 18173 33827 18207
rect 40601 18173 40635 18207
rect 43085 18173 43119 18207
rect 43177 18173 43211 18207
rect 20085 18105 20119 18139
rect 35817 18105 35851 18139
rect 36369 18105 36403 18139
rect 15025 18037 15059 18071
rect 20545 18037 20579 18071
rect 27629 18037 27663 18071
rect 31033 18037 31067 18071
rect 34529 18037 34563 18071
rect 36185 18037 36219 18071
rect 36921 18037 36955 18071
rect 37565 18037 37599 18071
rect 39221 18037 39255 18071
rect 41981 18037 42015 18071
rect 19901 17833 19935 17867
rect 19993 17833 20027 17867
rect 21097 17833 21131 17867
rect 22293 17833 22327 17867
rect 22937 17833 22971 17867
rect 23581 17833 23615 17867
rect 25973 17833 26007 17867
rect 27445 17833 27479 17867
rect 28457 17833 28491 17867
rect 28641 17833 28675 17867
rect 29837 17833 29871 17867
rect 31493 17833 31527 17867
rect 33517 17833 33551 17867
rect 34345 17833 34379 17867
rect 35081 17833 35115 17867
rect 35817 17833 35851 17867
rect 38945 17833 38979 17867
rect 40141 17833 40175 17867
rect 41337 17833 41371 17867
rect 43361 17833 43395 17867
rect 32137 17765 32171 17799
rect 38209 17765 38243 17799
rect 13737 17697 13771 17731
rect 14933 17697 14967 17731
rect 17325 17697 17359 17731
rect 20085 17697 20119 17731
rect 36277 17697 36311 17731
rect 36369 17697 36403 17731
rect 37841 17697 37875 17731
rect 41981 17697 42015 17731
rect 15485 17629 15519 17663
rect 15669 17629 15703 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 16589 17629 16623 17663
rect 17141 17629 17175 17663
rect 17509 17629 17543 17663
rect 18061 17629 18095 17663
rect 18429 17629 18463 17663
rect 19809 17629 19843 17663
rect 22017 17629 22051 17663
rect 23765 17629 23799 17663
rect 23949 17629 23983 17663
rect 24041 17629 24075 17663
rect 24593 17629 24627 17663
rect 27629 17629 27663 17663
rect 27721 17629 27755 17663
rect 27997 17629 28031 17663
rect 30021 17629 30055 17663
rect 30113 17629 30147 17663
rect 30389 17629 30423 17663
rect 30849 17629 30883 17663
rect 31033 17629 31067 17663
rect 32781 17629 32815 17663
rect 32965 17629 32999 17663
rect 33057 17629 33091 17663
rect 34161 17629 34195 17663
rect 34345 17629 34379 17663
rect 36645 17629 36679 17663
rect 36737 17629 36771 17663
rect 37013 17629 37047 17663
rect 37473 17629 37507 17663
rect 37657 17629 37691 17663
rect 37749 17629 37783 17663
rect 38025 17629 38059 17663
rect 38853 17629 38887 17663
rect 38945 17629 38979 17663
rect 40325 17629 40359 17663
rect 41153 17629 41187 17663
rect 42248 17629 42282 17663
rect 35035 17595 35069 17629
rect 16129 17561 16163 17595
rect 21281 17561 21315 17595
rect 22293 17561 22327 17595
rect 23121 17561 23155 17595
rect 24860 17561 24894 17595
rect 27813 17561 27847 17595
rect 28825 17561 28859 17595
rect 30205 17561 30239 17595
rect 30941 17561 30975 17595
rect 35265 17561 35299 17595
rect 38669 17561 38703 17595
rect 14289 17493 14323 17527
rect 14657 17493 14691 17527
rect 14749 17493 14783 17527
rect 20913 17493 20947 17527
rect 21081 17493 21115 17527
rect 22109 17493 22143 17527
rect 22753 17493 22787 17527
rect 22921 17493 22955 17527
rect 28625 17493 28659 17527
rect 32597 17493 32631 17527
rect 34897 17493 34931 17527
rect 36553 17493 36587 17527
rect 39129 17493 39163 17527
rect 14841 17289 14875 17323
rect 15669 17289 15703 17323
rect 18245 17289 18279 17323
rect 20545 17289 20579 17323
rect 25329 17289 25363 17323
rect 28549 17289 28583 17323
rect 33701 17289 33735 17323
rect 34621 17289 34655 17323
rect 36829 17289 36863 17323
rect 39129 17289 39163 17323
rect 41153 17289 41187 17323
rect 43177 17289 43211 17323
rect 15485 17221 15519 17255
rect 30757 17221 30791 17255
rect 31769 17221 31803 17255
rect 32566 17221 32600 17255
rect 35357 17221 35391 17255
rect 38669 17221 38703 17255
rect 41613 17221 41647 17255
rect 43269 17221 43303 17255
rect 12817 17153 12851 17187
rect 13717 17153 13751 17187
rect 15301 17153 15335 17187
rect 16865 17153 16899 17187
rect 17132 17153 17166 17187
rect 19165 17153 19199 17187
rect 19432 17153 19466 17187
rect 21281 17153 21315 17187
rect 22017 17153 22051 17187
rect 22273 17153 22307 17187
rect 25326 17153 25360 17187
rect 25789 17153 25823 17187
rect 27436 17153 27470 17187
rect 29009 17153 29043 17187
rect 31309 17153 31343 17187
rect 31401 17153 31435 17187
rect 31585 17153 31619 17187
rect 34437 17153 34471 17187
rect 34621 17153 34655 17187
rect 35541 17153 35575 17187
rect 36461 17153 36495 17187
rect 36645 17153 36679 17187
rect 37657 17153 37691 17187
rect 37749 17153 37783 17187
rect 37933 17153 37967 17187
rect 38945 17153 38979 17187
rect 39957 17153 39991 17187
rect 40153 17153 40187 17187
rect 41981 17153 42015 17187
rect 13461 17085 13495 17119
rect 27169 17085 27203 17119
rect 29285 17085 29319 17119
rect 29929 17085 29963 17119
rect 32321 17085 32355 17119
rect 36369 17085 36403 17119
rect 38853 17085 38887 17119
rect 43177 17085 43211 17119
rect 21465 17017 21499 17051
rect 25145 17017 25179 17051
rect 29101 17017 29135 17051
rect 37473 17017 37507 17051
rect 39957 17017 39991 17051
rect 42717 17017 42751 17051
rect 13001 16949 13035 16983
rect 23397 16949 23431 16983
rect 25697 16949 25731 16983
rect 29009 16949 29043 16983
rect 35173 16949 35207 16983
rect 37841 16949 37875 16983
rect 38669 16949 38703 16983
rect 13553 16745 13587 16779
rect 20913 16745 20947 16779
rect 22201 16745 22235 16779
rect 24593 16745 24627 16779
rect 27537 16745 27571 16779
rect 28549 16745 28583 16779
rect 30205 16745 30239 16779
rect 31585 16745 31619 16779
rect 31769 16745 31803 16779
rect 32413 16745 32447 16779
rect 32597 16745 32631 16779
rect 35173 16745 35207 16779
rect 36277 16745 36311 16779
rect 37473 16745 37507 16779
rect 37933 16745 37967 16779
rect 39037 16745 39071 16779
rect 40141 16745 40175 16779
rect 20453 16677 20487 16711
rect 21649 16677 21683 16711
rect 33517 16677 33551 16711
rect 14841 16609 14875 16643
rect 16313 16609 16347 16643
rect 17601 16609 17635 16643
rect 17693 16609 17727 16643
rect 19809 16609 19843 16643
rect 19993 16609 20027 16643
rect 22753 16609 22787 16643
rect 26433 16609 26467 16643
rect 28733 16609 28767 16643
rect 29009 16609 29043 16643
rect 30757 16609 30791 16643
rect 34989 16609 35023 16643
rect 36185 16609 36219 16643
rect 39129 16609 39163 16643
rect 41521 16609 41555 16643
rect 41705 16609 41739 16643
rect 42441 16609 42475 16643
rect 42533 16609 42567 16643
rect 13737 16541 13771 16575
rect 14657 16541 14691 16575
rect 15853 16541 15887 16575
rect 17509 16541 17543 16575
rect 18337 16541 18371 16575
rect 20085 16541 20119 16575
rect 21097 16541 21131 16575
rect 22569 16541 22603 16575
rect 25973 16541 26007 16575
rect 26525 16541 26559 16575
rect 26709 16541 26743 16575
rect 27721 16541 27755 16575
rect 27813 16541 27847 16575
rect 28089 16541 28123 16575
rect 28825 16541 28859 16575
rect 28917 16541 28951 16575
rect 30481 16541 30515 16575
rect 34069 16541 34103 16575
rect 34253 16541 34287 16575
rect 35173 16541 35207 16575
rect 36001 16541 36035 16575
rect 37197 16541 37231 16575
rect 37289 16541 37323 16575
rect 38117 16541 38151 16575
rect 38393 16541 38427 16575
rect 39221 16541 39255 16575
rect 40417 16541 40451 16575
rect 14749 16473 14783 16507
rect 22661 16473 22695 16507
rect 25728 16473 25762 16507
rect 26893 16473 26927 16507
rect 27905 16473 27939 16507
rect 30389 16473 30423 16507
rect 31737 16473 31771 16507
rect 31953 16473 31987 16507
rect 32781 16473 32815 16507
rect 34897 16473 34931 16507
rect 36277 16473 36311 16507
rect 37473 16473 37507 16507
rect 41429 16473 41463 16507
rect 42625 16473 42659 16507
rect 14289 16405 14323 16439
rect 15669 16405 15703 16439
rect 17141 16405 17175 16439
rect 18521 16405 18555 16439
rect 30573 16405 30607 16439
rect 32571 16405 32605 16439
rect 34069 16405 34103 16439
rect 35357 16405 35391 16439
rect 35817 16405 35851 16439
rect 37013 16405 37047 16439
rect 38301 16405 38335 16439
rect 38853 16405 38887 16439
rect 41061 16405 41095 16439
rect 42993 16405 43027 16439
rect 14657 16201 14691 16235
rect 15577 16201 15611 16235
rect 15945 16201 15979 16235
rect 17417 16201 17451 16235
rect 19625 16201 19659 16235
rect 21097 16201 21131 16235
rect 22385 16201 22419 16235
rect 26617 16201 26651 16235
rect 27629 16201 27663 16235
rect 36369 16201 36403 16235
rect 36921 16201 36955 16235
rect 38669 16201 38703 16235
rect 42073 16201 42107 16235
rect 43085 16201 43119 16235
rect 13522 16133 13556 16167
rect 16037 16133 16071 16167
rect 16957 16133 16991 16167
rect 18530 16133 18564 16167
rect 22477 16133 22511 16167
rect 25504 16133 25538 16167
rect 28089 16133 28123 16167
rect 32505 16133 32539 16167
rect 33333 16133 33367 16167
rect 34621 16133 34655 16167
rect 36185 16133 36219 16167
rect 42993 16133 43027 16167
rect 13277 16065 13311 16099
rect 18797 16065 18831 16099
rect 19441 16065 19475 16099
rect 21189 16065 21223 16099
rect 23213 16065 23247 16099
rect 27813 16065 27847 16099
rect 28917 16065 28951 16099
rect 29009 16065 29043 16099
rect 29828 16065 29862 16099
rect 31585 16065 31619 16099
rect 31769 16065 31803 16099
rect 32321 16065 32355 16099
rect 33149 16065 33183 16099
rect 33425 16065 33459 16099
rect 36001 16065 36035 16099
rect 38209 16065 38243 16099
rect 38393 16065 38427 16099
rect 38485 16065 38519 16099
rect 39313 16065 39347 16099
rect 40960 16065 40994 16099
rect 16221 15997 16255 16031
rect 21281 15997 21315 16031
rect 22569 15997 22603 16031
rect 25237 15997 25271 16031
rect 27905 15997 27939 16031
rect 29561 15997 29595 16031
rect 34253 15997 34287 16031
rect 34437 15997 34471 16031
rect 37473 15997 37507 16031
rect 38301 15997 38335 16031
rect 39129 15997 39163 16031
rect 39589 15997 39623 16031
rect 40693 15997 40727 16031
rect 43177 15997 43211 16031
rect 20085 15929 20119 15963
rect 30941 15929 30975 15963
rect 20729 15861 20763 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 28089 15861 28123 15895
rect 31401 15861 31435 15895
rect 32689 15861 32723 15895
rect 33149 15861 33183 15895
rect 34345 15861 34379 15895
rect 34621 15861 34655 15895
rect 35541 15861 35575 15895
rect 39497 15861 39531 15895
rect 40141 15861 40175 15895
rect 42625 15861 42659 15895
rect 16497 15657 16531 15691
rect 18613 15657 18647 15691
rect 22201 15657 22235 15691
rect 23397 15657 23431 15691
rect 27445 15657 27479 15691
rect 28181 15657 28215 15691
rect 30113 15657 30147 15691
rect 31217 15657 31251 15691
rect 31769 15657 31803 15691
rect 35817 15657 35851 15691
rect 36369 15657 36403 15691
rect 38209 15657 38243 15691
rect 43361 15657 43395 15691
rect 26525 15589 26559 15623
rect 38945 15589 38979 15623
rect 17969 15521 18003 15555
rect 20821 15521 20855 15555
rect 22753 15521 22787 15555
rect 23857 15521 23891 15555
rect 25789 15521 25823 15555
rect 25973 15521 26007 15555
rect 30573 15521 30607 15555
rect 32689 15521 32723 15555
rect 32781 15521 32815 15555
rect 32873 15521 32907 15555
rect 33609 15521 33643 15555
rect 36737 15521 36771 15555
rect 40969 15521 41003 15555
rect 41153 15521 41187 15555
rect 41981 15521 42015 15555
rect 14473 15453 14507 15487
rect 15117 15453 15151 15487
rect 15384 15453 15418 15487
rect 16957 15453 16991 15487
rect 18245 15453 18279 15487
rect 19533 15453 19567 15487
rect 20177 15453 20211 15487
rect 23029 15453 23063 15487
rect 28365 15453 28399 15487
rect 30297 15453 30331 15487
rect 30389 15453 30423 15487
rect 30481 15453 30515 15487
rect 32965 15453 32999 15487
rect 33517 15453 33551 15487
rect 33701 15453 33735 15487
rect 34161 15453 34195 15487
rect 34345 15453 34379 15487
rect 35081 15453 35115 15487
rect 35265 15453 35299 15487
rect 36553 15453 36587 15487
rect 36645 15453 36679 15487
rect 36829 15453 36863 15487
rect 37657 15453 37691 15487
rect 37749 15453 37783 15487
rect 37933 15453 37967 15487
rect 38025 15453 38059 15487
rect 39129 15453 39163 15487
rect 39221 15453 39255 15487
rect 21066 15385 21100 15419
rect 22937 15385 22971 15419
rect 34897 15385 34931 15419
rect 40877 15385 40911 15419
rect 42248 15385 42282 15419
rect 14289 15317 14323 15351
rect 17141 15317 17175 15351
rect 18153 15317 18187 15351
rect 19717 15317 19751 15351
rect 20361 15317 20395 15351
rect 25329 15317 25363 15351
rect 25697 15317 25731 15351
rect 28825 15317 28859 15351
rect 32505 15317 32539 15351
rect 34161 15317 34195 15351
rect 40509 15317 40543 15351
rect 14841 15113 14875 15147
rect 15301 15113 15335 15147
rect 15761 15113 15795 15147
rect 18245 15113 18279 15147
rect 19165 15113 19199 15147
rect 21373 15113 21407 15147
rect 22569 15113 22603 15147
rect 26065 15113 26099 15147
rect 28917 15113 28951 15147
rect 29469 15113 29503 15147
rect 32321 15113 32355 15147
rect 35173 15113 35207 15147
rect 36921 15113 36955 15147
rect 38301 15113 38335 15147
rect 41337 15113 41371 15147
rect 41981 15113 42015 15147
rect 42625 15113 42659 15147
rect 43361 15113 43395 15147
rect 23682 15045 23716 15079
rect 27813 15045 27847 15079
rect 27905 15045 27939 15079
rect 33333 15045 33367 15079
rect 34687 15045 34721 15079
rect 38485 15045 38519 15079
rect 38669 15045 38703 15079
rect 39589 15045 39623 15079
rect 13461 14977 13495 15011
rect 13728 14977 13762 15011
rect 15669 14977 15703 15011
rect 16865 14977 16899 15011
rect 17132 14977 17166 15011
rect 19993 14977 20027 15011
rect 20249 14977 20283 15011
rect 24952 14977 24986 15011
rect 27721 14977 27755 15011
rect 28089 14977 28123 15011
rect 28549 14977 28583 15011
rect 28733 14977 28767 15011
rect 29009 14977 29043 15011
rect 29653 14977 29687 15011
rect 29929 14977 29963 15011
rect 33701 14977 33735 15011
rect 34805 14977 34839 15011
rect 34897 14977 34931 15011
rect 34989 14977 35023 15011
rect 35825 14977 35859 15011
rect 36001 14977 36035 15011
rect 36461 14977 36495 15011
rect 36737 14977 36771 15011
rect 37473 14977 37507 15011
rect 37657 14977 37691 15011
rect 39405 14977 39439 15011
rect 39773 14977 39807 15011
rect 40509 14977 40543 15011
rect 41521 14977 41555 15011
rect 42809 14977 42843 15011
rect 15945 14909 15979 14943
rect 18889 14909 18923 14943
rect 19073 14909 19107 14943
rect 23949 14909 23983 14943
rect 24685 14909 24719 14943
rect 29837 14909 29871 14943
rect 34529 14909 34563 14943
rect 35909 14909 35943 14943
rect 36645 14909 36679 14943
rect 40325 14841 40359 14875
rect 19533 14773 19567 14807
rect 27537 14773 27571 14807
rect 29745 14773 29779 14807
rect 33149 14773 33183 14807
rect 33333 14773 33367 14807
rect 36461 14773 36495 14807
rect 37749 14773 37783 14807
rect 17049 14569 17083 14603
rect 20821 14569 20855 14603
rect 22385 14569 22419 14603
rect 25053 14569 25087 14603
rect 27261 14569 27295 14603
rect 29193 14569 29227 14603
rect 29745 14569 29779 14603
rect 34897 14569 34931 14603
rect 35081 14569 35115 14603
rect 36277 14569 36311 14603
rect 38577 14569 38611 14603
rect 39313 14569 39347 14603
rect 41245 14569 41279 14603
rect 41797 14569 41831 14603
rect 14473 14501 14507 14535
rect 16405 14501 16439 14535
rect 33333 14501 33367 14535
rect 39129 14501 39163 14535
rect 15393 14433 15427 14467
rect 15485 14433 15519 14467
rect 17509 14433 17543 14467
rect 17693 14433 17727 14467
rect 19441 14433 19475 14467
rect 25881 14433 25915 14467
rect 30021 14433 30055 14467
rect 31678 14433 31712 14467
rect 31769 14433 31803 14467
rect 31953 14433 31987 14467
rect 36369 14433 36403 14467
rect 40417 14433 40451 14467
rect 15301 14365 15335 14399
rect 17417 14365 17451 14399
rect 18705 14365 18739 14399
rect 25237 14365 25271 14399
rect 28549 14365 28583 14399
rect 28733 14365 28767 14399
rect 28825 14365 28859 14399
rect 28917 14365 28951 14399
rect 29929 14365 29963 14399
rect 30113 14365 30147 14399
rect 30205 14365 30239 14399
rect 31861 14365 31895 14399
rect 32505 14365 32539 14399
rect 32689 14365 32723 14399
rect 33149 14365 33183 14399
rect 33333 14365 33367 14399
rect 33793 14365 33827 14399
rect 33977 14365 34011 14399
rect 36093 14365 36127 14399
rect 36185 14365 36219 14399
rect 37013 14365 37047 14399
rect 37197 14365 37231 14399
rect 37749 14365 37783 14399
rect 38485 14365 38519 14399
rect 38669 14365 38703 14399
rect 40049 14365 40083 14399
rect 40509 14365 40543 14399
rect 43361 14365 43395 14399
rect 19686 14297 19720 14331
rect 26148 14297 26182 14331
rect 33885 14297 33919 14331
rect 35265 14297 35299 14331
rect 36829 14297 36863 14331
rect 39497 14297 39531 14331
rect 42349 14297 42383 14331
rect 43085 14297 43119 14331
rect 14933 14229 14967 14263
rect 18889 14229 18923 14263
rect 30757 14229 30791 14263
rect 31493 14229 31527 14263
rect 32505 14229 32539 14263
rect 35055 14229 35089 14263
rect 37933 14229 37967 14263
rect 39297 14229 39331 14263
rect 15577 14025 15611 14059
rect 16221 14025 16255 14059
rect 17877 14025 17911 14059
rect 19809 14025 19843 14059
rect 20269 14025 20303 14059
rect 20637 14025 20671 14059
rect 22845 14025 22879 14059
rect 24869 14025 24903 14059
rect 25237 14025 25271 14059
rect 25329 14025 25363 14059
rect 27169 14025 27203 14059
rect 30113 14025 30147 14059
rect 30481 14025 30515 14059
rect 31585 14025 31619 14059
rect 34713 14025 34747 14059
rect 37657 14025 37691 14059
rect 38301 14025 38335 14059
rect 41153 14025 41187 14059
rect 42625 14025 42659 14059
rect 42993 14025 43027 14059
rect 20729 13957 20763 13991
rect 22937 13957 22971 13991
rect 28282 13957 28316 13991
rect 31769 13957 31803 13991
rect 33241 13957 33275 13991
rect 33425 13957 33459 13991
rect 38945 13957 38979 13991
rect 41981 13957 42015 13991
rect 14197 13889 14231 13923
rect 14464 13889 14498 13923
rect 18429 13889 18463 13923
rect 18696 13889 18730 13923
rect 24225 13889 24259 13923
rect 26433 13889 26467 13923
rect 26617 13889 26651 13923
rect 29101 13889 29135 13923
rect 29285 13889 29319 13923
rect 29377 13889 29411 13923
rect 29469 13889 29503 13923
rect 30297 13889 30331 13923
rect 30573 13889 30607 13923
rect 31493 13889 31527 13923
rect 32505 13889 32539 13923
rect 33609 13889 33643 13923
rect 34897 13889 34931 13923
rect 35357 13889 35391 13923
rect 35535 13889 35569 13923
rect 36461 13889 36495 13923
rect 36645 13889 36679 13923
rect 37473 13889 37507 13923
rect 38209 13889 38243 13923
rect 38393 13889 38427 13923
rect 38853 13889 38887 13923
rect 39037 13889 39071 13923
rect 39589 13889 39623 13923
rect 39957 13889 39991 13923
rect 40325 13889 40359 13923
rect 20913 13821 20947 13855
rect 23029 13821 23063 13855
rect 25513 13821 25547 13855
rect 28549 13821 28583 13855
rect 32689 13821 32723 13855
rect 35449 13821 35483 13855
rect 36553 13821 36587 13855
rect 41245 13821 41279 13855
rect 41429 13821 41463 13855
rect 43085 13821 43119 13855
rect 43269 13821 43303 13855
rect 24409 13753 24443 13787
rect 40785 13753 40819 13787
rect 22477 13685 22511 13719
rect 26525 13685 26559 13719
rect 29653 13685 29687 13719
rect 31769 13685 31803 13719
rect 32321 13685 32355 13719
rect 14657 13481 14691 13515
rect 15945 13481 15979 13515
rect 19441 13481 19475 13515
rect 23673 13481 23707 13515
rect 25973 13481 26007 13515
rect 26801 13481 26835 13515
rect 29837 13481 29871 13515
rect 31769 13481 31803 13515
rect 33517 13481 33551 13515
rect 35725 13481 35759 13515
rect 37473 13481 37507 13515
rect 38669 13481 38703 13515
rect 43269 13481 43303 13515
rect 20545 13413 20579 13447
rect 29193 13413 29227 13447
rect 33609 13413 33643 13447
rect 34989 13413 35023 13447
rect 36001 13413 36035 13447
rect 21649 13345 21683 13379
rect 26985 13345 27019 13379
rect 27445 13345 27479 13379
rect 30941 13345 30975 13379
rect 31953 13345 31987 13379
rect 32045 13345 32079 13379
rect 33425 13345 33459 13379
rect 36093 13345 36127 13379
rect 14841 13277 14875 13311
rect 19625 13277 19659 13311
rect 21557 13277 21591 13311
rect 22293 13277 22327 13311
rect 24593 13277 24627 13311
rect 27077 13277 27111 13311
rect 28917 13277 28951 13311
rect 29009 13277 29043 13311
rect 30021 13277 30055 13311
rect 30297 13277 30331 13311
rect 31033 13277 31067 13311
rect 31125 13277 31159 13311
rect 31217 13277 31251 13311
rect 32137 13277 32171 13311
rect 32229 13277 32263 13311
rect 33701 13277 33735 13311
rect 33885 13277 33919 13311
rect 35173 13277 35207 13311
rect 35909 13277 35943 13311
rect 36185 13277 36219 13311
rect 37105 13277 37139 13311
rect 37933 13277 37967 13311
rect 38117 13277 38151 13311
rect 38577 13277 38611 13311
rect 38761 13277 38795 13311
rect 39313 13277 39347 13311
rect 40049 13277 40083 13311
rect 41889 13277 41923 13311
rect 21465 13209 21499 13243
rect 22560 13209 22594 13243
rect 24860 13209 24894 13243
rect 27353 13209 27387 13243
rect 27905 13209 27939 13243
rect 37289 13209 37323 13243
rect 40294 13209 40328 13243
rect 42156 13209 42190 13243
rect 21097 13141 21131 13175
rect 30205 13141 30239 13175
rect 30757 13141 30791 13175
rect 33149 13141 33183 13175
rect 38025 13141 38059 13175
rect 39497 13141 39531 13175
rect 41429 13141 41463 13175
rect 20177 12937 20211 12971
rect 21465 12937 21499 12971
rect 23397 12937 23431 12971
rect 25789 12937 25823 12971
rect 26525 12937 26559 12971
rect 28457 12937 28491 12971
rect 31677 12937 31711 12971
rect 32965 12937 32999 12971
rect 33701 12937 33735 12971
rect 37841 12937 37875 12971
rect 39957 12937 39991 12971
rect 40417 12937 40451 12971
rect 41429 12937 41463 12971
rect 42073 12937 42107 12971
rect 42625 12937 42659 12971
rect 42993 12937 43027 12971
rect 43085 12937 43119 12971
rect 22262 12869 22296 12903
rect 34713 12869 34747 12903
rect 35633 12869 35667 12903
rect 21281 12801 21315 12835
rect 22017 12801 22051 12835
rect 27169 12801 27203 12835
rect 29570 12801 29604 12835
rect 30757 12801 30791 12835
rect 30941 12801 30975 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 32505 12801 32539 12835
rect 33609 12801 33643 12835
rect 33793 12801 33827 12835
rect 34437 12801 34471 12835
rect 35817 12801 35851 12835
rect 36277 12801 36311 12835
rect 36461 12801 36495 12835
rect 38025 12801 38059 12835
rect 38209 12801 38243 12835
rect 38761 12801 38795 12835
rect 39037 12801 39071 12835
rect 40325 12801 40359 12835
rect 41889 12801 41923 12835
rect 29837 12733 29871 12767
rect 30665 12733 30699 12767
rect 32597 12733 32631 12767
rect 34621 12733 34655 12767
rect 35449 12733 35483 12767
rect 38669 12733 38703 12767
rect 40601 12733 40635 12767
rect 43177 12733 43211 12767
rect 36277 12665 36311 12699
rect 27353 12597 27387 12631
rect 31125 12597 31159 12631
rect 32321 12597 32355 12631
rect 34253 12597 34287 12631
rect 34621 12597 34655 12631
rect 22661 12393 22695 12427
rect 26433 12393 26467 12427
rect 27353 12393 27387 12427
rect 32229 12393 32263 12427
rect 37105 12393 37139 12427
rect 38669 12393 38703 12427
rect 40601 12393 40635 12427
rect 41521 12393 41555 12427
rect 29929 12325 29963 12359
rect 35817 12325 35851 12359
rect 40049 12325 40083 12359
rect 27997 12257 28031 12291
rect 32321 12257 32355 12291
rect 33977 12257 34011 12291
rect 34069 12257 34103 12291
rect 34897 12257 34931 12291
rect 36277 12257 36311 12291
rect 41981 12257 42015 12291
rect 22477 12189 22511 12223
rect 25605 12189 25639 12223
rect 26157 12189 26191 12223
rect 27813 12189 27847 12223
rect 29745 12189 29779 12223
rect 29929 12189 29963 12223
rect 30573 12189 30607 12223
rect 30665 12189 30699 12223
rect 30849 12189 30883 12223
rect 30941 12189 30975 12223
rect 32229 12189 32263 12223
rect 33793 12189 33827 12223
rect 34161 12189 34195 12223
rect 34345 12189 34379 12223
rect 35265 12189 35299 12223
rect 36369 12189 36403 12223
rect 36553 12189 36587 12223
rect 38393 12189 38427 12223
rect 39221 12189 39255 12223
rect 39405 12189 39439 12223
rect 32689 12121 32723 12155
rect 33609 12121 33643 12155
rect 35081 12121 35115 12155
rect 37289 12121 37323 12155
rect 37473 12121 37507 12155
rect 42226 12121 42260 12155
rect 25421 12053 25455 12087
rect 27721 12053 27755 12087
rect 28641 12053 28675 12087
rect 29193 12053 29227 12087
rect 30389 12053 30423 12087
rect 32045 12053 32079 12087
rect 39221 12053 39255 12087
rect 43361 12053 43395 12087
rect 26525 11849 26559 11883
rect 28549 11849 28583 11883
rect 29469 11849 29503 11883
rect 30849 11849 30883 11883
rect 32597 11849 32631 11883
rect 38301 11849 38335 11883
rect 40509 11849 40543 11883
rect 40877 11849 40911 11883
rect 42073 11849 42107 11883
rect 42625 11849 42659 11883
rect 43085 11849 43119 11883
rect 25412 11781 25446 11815
rect 27436 11781 27470 11815
rect 33885 11781 33919 11815
rect 34713 11781 34747 11815
rect 39681 11781 39715 11815
rect 25145 11713 25179 11747
rect 27169 11713 27203 11747
rect 29377 11713 29411 11747
rect 30757 11713 30791 11747
rect 32781 11713 32815 11747
rect 32873 11713 32907 11747
rect 32965 11713 32999 11747
rect 33149 11713 33183 11747
rect 33977 11713 34011 11747
rect 34621 11713 34655 11747
rect 34805 11713 34839 11747
rect 34989 11713 35023 11747
rect 35633 11713 35667 11747
rect 35817 11713 35851 11747
rect 35909 11713 35943 11747
rect 36645 11713 36679 11747
rect 36829 11713 36863 11747
rect 37473 11713 37507 11747
rect 37657 11713 37691 11747
rect 37749 11713 37783 11747
rect 38485 11713 38519 11747
rect 38669 11713 38703 11747
rect 39773 11713 39807 11747
rect 40969 11713 41003 11747
rect 41889 11713 41923 11747
rect 42993 11713 43027 11747
rect 29653 11645 29687 11679
rect 30941 11645 30975 11679
rect 39957 11645 39991 11679
rect 41061 11645 41095 11679
rect 43177 11645 43211 11679
rect 31585 11577 31619 11611
rect 29009 11509 29043 11543
rect 30389 11509 30423 11543
rect 34437 11509 34471 11543
rect 35449 11509 35483 11543
rect 39313 11509 39347 11543
rect 25605 11305 25639 11339
rect 29193 11305 29227 11339
rect 31125 11305 31159 11339
rect 32229 11305 32263 11339
rect 37013 11305 37047 11339
rect 41797 11305 41831 11339
rect 42349 11305 42383 11339
rect 36553 11237 36587 11271
rect 26065 11169 26099 11203
rect 26249 11169 26283 11203
rect 27813 11169 27847 11203
rect 33609 11169 33643 11203
rect 35173 11169 35207 11203
rect 38945 11169 38979 11203
rect 42809 11169 42843 11203
rect 42901 11169 42935 11203
rect 29745 11101 29779 11135
rect 34161 11101 34195 11135
rect 37013 11101 37047 11135
rect 37197 11101 37231 11135
rect 38117 11101 38151 11135
rect 38301 11101 38335 11135
rect 40417 11101 40451 11135
rect 42717 11101 42751 11135
rect 25973 11033 26007 11067
rect 28080 11033 28114 11067
rect 30012 11033 30046 11067
rect 33342 11033 33376 11067
rect 35418 11033 35452 11067
rect 39037 11033 39071 11067
rect 40684 11033 40718 11067
rect 34345 10965 34379 10999
rect 37933 10965 37967 10999
rect 39129 10965 39163 10999
rect 39497 10965 39531 10999
rect 28365 10761 28399 10795
rect 29929 10761 29963 10795
rect 31769 10761 31803 10795
rect 32413 10761 32447 10795
rect 34437 10761 34471 10795
rect 34897 10761 34931 10795
rect 35725 10761 35759 10795
rect 40141 10761 40175 10795
rect 41061 10761 41095 10795
rect 41153 10761 41187 10795
rect 42625 10761 42659 10795
rect 43361 10761 43395 10795
rect 30634 10693 30668 10727
rect 33977 10693 34011 10727
rect 37841 10693 37875 10727
rect 38025 10693 38059 10727
rect 28549 10625 28583 10659
rect 29745 10625 29779 10659
rect 30389 10625 30423 10659
rect 32597 10625 32631 10659
rect 33057 10625 33091 10659
rect 34805 10625 34839 10659
rect 38761 10625 38795 10659
rect 39028 10625 39062 10659
rect 32781 10557 32815 10591
rect 32873 10557 32907 10591
rect 34989 10557 35023 10591
rect 41245 10557 41279 10591
rect 32689 10489 32723 10523
rect 40693 10421 40727 10455
rect 41981 10421 42015 10455
rect 30573 10217 30607 10251
rect 30941 10217 30975 10251
rect 37841 10217 37875 10251
rect 39221 10217 39255 10251
rect 40049 10217 40083 10251
rect 40693 10217 40727 10251
rect 42073 10217 42107 10251
rect 31033 10081 31067 10115
rect 43085 10081 43119 10115
rect 30757 10013 30791 10047
rect 39405 10013 39439 10047
rect 40877 10013 40911 10047
rect 43361 10013 43395 10047
rect 41429 9877 41463 9911
rect 40141 9673 40175 9707
rect 43269 9673 43303 9707
rect 40877 9605 40911 9639
rect 41613 9605 41647 9639
rect 42809 9605 42843 9639
rect 41429 9129 41463 9163
rect 41889 9129 41923 9163
rect 43361 9129 43395 9163
rect 42809 9061 42843 9095
rect 42809 8585 42843 8619
rect 43269 8585 43303 8619
rect 43361 8041 43395 8075
rect 43085 6341 43119 6375
rect 43361 6273 43395 6307
rect 43361 5865 43395 5899
rect 43361 2805 43395 2839
rect 43085 2465 43119 2499
rect 43361 2397 43395 2431
<< metal1 >>
rect 29454 44072 29460 44124
rect 29512 44112 29518 44124
rect 31754 44112 31760 44124
rect 29512 44084 31760 44112
rect 29512 44072 29518 44084
rect 31754 44072 31760 44084
rect 31812 44072 31818 44124
rect 34146 44072 34152 44124
rect 34204 44112 34210 44124
rect 34606 44112 34612 44124
rect 34204 44084 34612 44112
rect 34204 44072 34210 44084
rect 34606 44072 34612 44084
rect 34664 44072 34670 44124
rect 1104 42458 43884 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 43884 42458
rect 1104 42384 43884 42406
rect 27062 42304 27068 42356
rect 27120 42344 27126 42356
rect 35621 42347 35679 42353
rect 27120 42316 27936 42344
rect 27120 42304 27126 42316
rect 26605 42279 26663 42285
rect 26605 42245 26617 42279
rect 26651 42276 26663 42279
rect 27522 42276 27528 42288
rect 26651 42248 27528 42276
rect 26651 42245 26663 42248
rect 26605 42239 26663 42245
rect 27522 42236 27528 42248
rect 27580 42236 27586 42288
rect 27908 42285 27936 42316
rect 35621 42313 35633 42347
rect 35667 42344 35679 42347
rect 37918 42344 37924 42356
rect 35667 42316 37924 42344
rect 35667 42313 35679 42316
rect 35621 42307 35679 42313
rect 37918 42304 37924 42316
rect 37976 42304 37982 42356
rect 27893 42279 27951 42285
rect 27893 42245 27905 42279
rect 27939 42276 27951 42279
rect 29825 42279 29883 42285
rect 29825 42276 29837 42279
rect 27939 42248 29837 42276
rect 27939 42245 27951 42248
rect 27893 42239 27951 42245
rect 29825 42245 29837 42248
rect 29871 42276 29883 42279
rect 29871 42248 35894 42276
rect 29871 42245 29883 42248
rect 29825 42239 29883 42245
rect 13814 42168 13820 42220
rect 13872 42208 13878 42220
rect 14277 42211 14335 42217
rect 14277 42208 14289 42211
rect 13872 42180 14289 42208
rect 13872 42168 13878 42180
rect 14277 42177 14289 42180
rect 14323 42177 14335 42211
rect 14277 42171 14335 42177
rect 15378 42168 15384 42220
rect 15436 42208 15442 42220
rect 15473 42211 15531 42217
rect 15473 42208 15485 42211
rect 15436 42180 15485 42208
rect 15436 42168 15442 42180
rect 15473 42177 15485 42180
rect 15519 42177 15531 42211
rect 15473 42171 15531 42177
rect 20625 42211 20683 42217
rect 20625 42177 20637 42211
rect 20671 42208 20683 42211
rect 20714 42208 20720 42220
rect 20671 42180 20720 42208
rect 20671 42177 20683 42180
rect 20625 42171 20683 42177
rect 20714 42168 20720 42180
rect 20772 42168 20778 42220
rect 22738 42168 22744 42220
rect 22796 42168 22802 42220
rect 25406 42168 25412 42220
rect 25464 42168 25470 42220
rect 27338 42168 27344 42220
rect 27396 42168 27402 42220
rect 27430 42168 27436 42220
rect 27488 42208 27494 42220
rect 28353 42211 28411 42217
rect 28353 42208 28365 42211
rect 27488 42180 28365 42208
rect 27488 42168 27494 42180
rect 28353 42177 28365 42180
rect 28399 42177 28411 42211
rect 28353 42171 28411 42177
rect 30650 42168 30656 42220
rect 30708 42168 30714 42220
rect 32306 42168 32312 42220
rect 32364 42168 32370 42220
rect 34790 42168 34796 42220
rect 34848 42208 34854 42220
rect 34885 42211 34943 42217
rect 34885 42208 34897 42211
rect 34848 42180 34897 42208
rect 34848 42168 34854 42180
rect 34885 42177 34897 42180
rect 34931 42177 34943 42211
rect 35866 42208 35894 42248
rect 37550 42236 37556 42288
rect 37608 42276 37614 42288
rect 41693 42279 41751 42285
rect 41693 42276 41705 42279
rect 37608 42248 41705 42276
rect 37608 42236 37614 42248
rect 41693 42245 41705 42248
rect 41739 42245 41751 42279
rect 41693 42239 41751 42245
rect 38378 42208 38384 42220
rect 35866 42180 38384 42208
rect 34885 42171 34943 42177
rect 38378 42168 38384 42180
rect 38436 42168 38442 42220
rect 43349 42211 43407 42217
rect 43349 42208 43361 42211
rect 39224 42180 43361 42208
rect 19981 42143 20039 42149
rect 19981 42109 19993 42143
rect 20027 42140 20039 42143
rect 33781 42143 33839 42149
rect 20027 42112 31708 42140
rect 20027 42109 20039 42112
rect 19981 42103 20039 42109
rect 21450 42032 21456 42084
rect 21508 42072 21514 42084
rect 29638 42072 29644 42084
rect 21508 42044 29644 42072
rect 21508 42032 21514 42044
rect 29638 42032 29644 42044
rect 29696 42072 29702 42084
rect 31389 42075 31447 42081
rect 31389 42072 31401 42075
rect 29696 42044 31401 42072
rect 29696 42032 29702 42044
rect 31389 42041 31401 42044
rect 31435 42072 31447 42075
rect 31570 42072 31576 42084
rect 31435 42044 31576 42072
rect 31435 42041 31447 42044
rect 31389 42035 31447 42041
rect 31570 42032 31576 42044
rect 31628 42032 31634 42084
rect 31680 42072 31708 42112
rect 33781 42109 33793 42143
rect 33827 42140 33839 42143
rect 34330 42140 34336 42152
rect 33827 42112 34336 42140
rect 33827 42109 33839 42112
rect 33781 42103 33839 42109
rect 34330 42100 34336 42112
rect 34388 42100 34394 42152
rect 37553 42143 37611 42149
rect 37553 42109 37565 42143
rect 37599 42140 37611 42143
rect 38194 42140 38200 42152
rect 37599 42112 38200 42140
rect 37599 42109 37611 42112
rect 37553 42103 37611 42109
rect 38194 42100 38200 42112
rect 38252 42140 38258 42152
rect 39117 42143 39175 42149
rect 39117 42140 39129 42143
rect 38252 42112 39129 42140
rect 38252 42100 38258 42112
rect 39117 42109 39129 42112
rect 39163 42109 39175 42143
rect 39117 42103 39175 42109
rect 39224 42072 39252 42180
rect 43349 42177 43361 42180
rect 43395 42208 43407 42211
rect 43990 42208 43996 42220
rect 43395 42180 43996 42208
rect 43395 42177 43407 42180
rect 43349 42171 43407 42177
rect 43990 42168 43996 42180
rect 44048 42168 44054 42220
rect 42794 42100 42800 42152
rect 42852 42140 42858 42152
rect 43073 42143 43131 42149
rect 43073 42140 43085 42143
rect 42852 42112 43085 42140
rect 42852 42100 42858 42112
rect 43073 42109 43085 42112
rect 43119 42109 43131 42143
rect 43073 42103 43131 42109
rect 31680 42044 39252 42072
rect 39298 42032 39304 42084
rect 39356 42072 39362 42084
rect 41141 42075 41199 42081
rect 41141 42072 41153 42075
rect 39356 42044 41153 42072
rect 39356 42032 39362 42044
rect 41141 42041 41153 42044
rect 41187 42041 41199 42075
rect 41141 42035 41199 42041
rect 20438 41964 20444 42016
rect 20496 41964 20502 42016
rect 22094 41964 22100 42016
rect 22152 41964 22158 42016
rect 22554 41964 22560 42016
rect 22612 41964 22618 42016
rect 23382 41964 23388 42016
rect 23440 42004 23446 42016
rect 23937 42007 23995 42013
rect 23937 42004 23949 42007
rect 23440 41976 23949 42004
rect 23440 41964 23446 41976
rect 23937 41973 23949 41976
rect 23983 41973 23995 42007
rect 23937 41967 23995 41973
rect 24765 42007 24823 42013
rect 24765 41973 24777 42007
rect 24811 42004 24823 42007
rect 25038 42004 25044 42016
rect 24811 41976 25044 42004
rect 24811 41973 24823 41976
rect 24765 41967 24823 41973
rect 25038 41964 25044 41976
rect 25096 41964 25102 42016
rect 25222 41964 25228 42016
rect 25280 41964 25286 42016
rect 26053 42007 26111 42013
rect 26053 41973 26065 42007
rect 26099 42004 26111 42007
rect 26602 42004 26608 42016
rect 26099 41976 26608 42004
rect 26099 41973 26111 41976
rect 26053 41967 26111 41973
rect 26602 41964 26608 41976
rect 26660 42004 26666 42016
rect 27062 42004 27068 42016
rect 26660 41976 27068 42004
rect 26660 41964 26666 41976
rect 27062 41964 27068 41976
rect 27120 41964 27126 42016
rect 27154 41964 27160 42016
rect 27212 41964 27218 42016
rect 28994 41964 29000 42016
rect 29052 42004 29058 42016
rect 29089 42007 29147 42013
rect 29089 42004 29101 42007
rect 29052 41976 29101 42004
rect 29052 41964 29058 41976
rect 29089 41973 29101 41976
rect 29135 41973 29147 42007
rect 29089 41967 29147 41973
rect 30834 41964 30840 42016
rect 30892 41964 30898 42016
rect 32493 42007 32551 42013
rect 32493 41973 32505 42007
rect 32539 42004 32551 42007
rect 32582 42004 32588 42016
rect 32539 41976 32588 42004
rect 32539 41973 32551 41976
rect 32493 41967 32551 41973
rect 32582 41964 32588 41976
rect 32640 41964 32646 42016
rect 33229 42007 33287 42013
rect 33229 41973 33241 42007
rect 33275 42004 33287 42007
rect 33594 42004 33600 42016
rect 33275 41976 33600 42004
rect 33275 41973 33287 41976
rect 33229 41967 33287 41973
rect 33594 41964 33600 41976
rect 33652 41964 33658 42016
rect 34238 41964 34244 42016
rect 34296 41964 34302 42016
rect 35069 42007 35127 42013
rect 35069 41973 35081 42007
rect 35115 42004 35127 42007
rect 35434 42004 35440 42016
rect 35115 41976 35440 42004
rect 35115 41973 35127 41976
rect 35069 41967 35127 41973
rect 35434 41964 35440 41976
rect 35492 41964 35498 42016
rect 36078 41964 36084 42016
rect 36136 41964 36142 42016
rect 36170 41964 36176 42016
rect 36228 42004 36234 42016
rect 36633 42007 36691 42013
rect 36633 42004 36645 42007
rect 36228 41976 36645 42004
rect 36228 41964 36234 41976
rect 36633 41973 36645 41976
rect 36679 41973 36691 42007
rect 36633 41967 36691 41973
rect 38105 42007 38163 42013
rect 38105 41973 38117 42007
rect 38151 42004 38163 42007
rect 38378 42004 38384 42016
rect 38151 41976 38384 42004
rect 38151 41973 38163 41976
rect 38105 41967 38163 41973
rect 38378 41964 38384 41976
rect 38436 41964 38442 42016
rect 38657 42007 38715 42013
rect 38657 41973 38669 42007
rect 38703 42004 38715 42007
rect 38930 42004 38936 42016
rect 38703 41976 38936 42004
rect 38703 41973 38715 41976
rect 38657 41967 38715 41973
rect 38930 41964 38936 41976
rect 38988 41964 38994 42016
rect 40129 42007 40187 42013
rect 40129 41973 40141 42007
rect 40175 42004 40187 42007
rect 40494 42004 40500 42016
rect 40175 41976 40500 42004
rect 40175 41973 40187 41976
rect 40129 41967 40187 41973
rect 40494 41964 40500 41976
rect 40552 41964 40558 42016
rect 40586 41964 40592 42016
rect 40644 41964 40650 42016
rect 1104 41914 43884 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 43884 41914
rect 1104 41840 43884 41862
rect 31478 41760 31484 41812
rect 31536 41800 31542 41812
rect 37550 41800 37556 41812
rect 31536 41772 37556 41800
rect 31536 41760 31542 41772
rect 37550 41760 37556 41772
rect 37608 41760 37614 41812
rect 41966 41760 41972 41812
rect 42024 41800 42030 41812
rect 42061 41803 42119 41809
rect 42061 41800 42073 41803
rect 42024 41772 42073 41800
rect 42024 41760 42030 41772
rect 42061 41769 42073 41772
rect 42107 41769 42119 41803
rect 42061 41763 42119 41769
rect 38841 41735 38899 41741
rect 38841 41701 38853 41735
rect 38887 41732 38899 41735
rect 39390 41732 39396 41744
rect 38887 41704 39396 41732
rect 38887 41701 38899 41704
rect 38841 41695 38899 41701
rect 39390 41692 39396 41704
rect 39448 41692 39454 41744
rect 29638 41624 29644 41676
rect 29696 41664 29702 41676
rect 29733 41667 29791 41673
rect 29733 41664 29745 41667
rect 29696 41636 29745 41664
rect 29696 41624 29702 41636
rect 29733 41633 29745 41636
rect 29779 41633 29791 41667
rect 29733 41627 29791 41633
rect 31570 41624 31576 41676
rect 31628 41624 31634 41676
rect 40126 41624 40132 41676
rect 40184 41624 40190 41676
rect 19981 41599 20039 41605
rect 19981 41565 19993 41599
rect 20027 41596 20039 41599
rect 20070 41596 20076 41608
rect 20027 41568 20076 41596
rect 20027 41565 20039 41568
rect 19981 41559 20039 41565
rect 20070 41556 20076 41568
rect 20128 41596 20134 41608
rect 22554 41605 22560 41608
rect 22281 41599 22339 41605
rect 22281 41596 22293 41599
rect 20128 41568 22293 41596
rect 20128 41556 20134 41568
rect 22281 41565 22293 41568
rect 22327 41565 22339 41599
rect 22548 41596 22560 41605
rect 22515 41568 22560 41596
rect 22281 41559 22339 41565
rect 22548 41559 22560 41568
rect 22554 41556 22560 41559
rect 22612 41556 22618 41608
rect 24946 41556 24952 41608
rect 25004 41596 25010 41608
rect 25041 41599 25099 41605
rect 25041 41596 25053 41599
rect 25004 41568 25053 41596
rect 25004 41556 25010 41568
rect 25041 41565 25053 41568
rect 25087 41565 25099 41599
rect 25041 41559 25099 41565
rect 25308 41599 25366 41605
rect 25308 41565 25320 41599
rect 25354 41565 25366 41599
rect 26878 41596 26884 41608
rect 25308 41559 25366 41565
rect 26206 41568 26884 41596
rect 20248 41531 20306 41537
rect 20248 41497 20260 41531
rect 20294 41528 20306 41531
rect 20438 41528 20444 41540
rect 20294 41500 20444 41528
rect 20294 41497 20306 41500
rect 20248 41491 20306 41497
rect 20438 41488 20444 41500
rect 20496 41488 20502 41540
rect 21358 41420 21364 41472
rect 21416 41420 21422 41472
rect 23661 41463 23719 41469
rect 23661 41429 23673 41463
rect 23707 41460 23719 41463
rect 24118 41460 24124 41472
rect 23707 41432 24124 41460
rect 23707 41429 23719 41432
rect 23661 41423 23719 41429
rect 24118 41420 24124 41432
rect 24176 41420 24182 41472
rect 25056 41460 25084 41559
rect 25222 41488 25228 41540
rect 25280 41528 25286 41540
rect 25332 41528 25360 41559
rect 25280 41500 25360 41528
rect 25280 41488 25286 41500
rect 26206 41460 26234 41568
rect 26878 41556 26884 41568
rect 26936 41556 26942 41608
rect 27154 41605 27160 41608
rect 27148 41596 27160 41605
rect 27115 41568 27160 41596
rect 27148 41559 27160 41568
rect 27154 41556 27160 41559
rect 27212 41556 27218 41608
rect 28721 41599 28779 41605
rect 28721 41565 28733 41599
rect 28767 41596 28779 41599
rect 29086 41596 29092 41608
rect 28767 41568 29092 41596
rect 28767 41565 28779 41568
rect 28721 41559 28779 41565
rect 29086 41556 29092 41568
rect 29144 41556 29150 41608
rect 30834 41556 30840 41608
rect 30892 41596 30898 41608
rect 31829 41599 31887 41605
rect 31829 41596 31841 41599
rect 30892 41568 31841 41596
rect 30892 41556 30898 41568
rect 31829 41565 31841 41568
rect 31875 41565 31887 41599
rect 31829 41559 31887 41565
rect 35434 41556 35440 41608
rect 35492 41596 35498 41608
rect 35998 41599 36056 41605
rect 35998 41596 36010 41599
rect 35492 41568 36010 41596
rect 35492 41556 35498 41568
rect 35998 41565 36010 41568
rect 36044 41565 36056 41599
rect 35998 41559 36056 41565
rect 36265 41599 36323 41605
rect 36265 41565 36277 41599
rect 36311 41596 36323 41599
rect 36722 41596 36728 41608
rect 36311 41568 36728 41596
rect 36311 41565 36323 41568
rect 36265 41559 36323 41565
rect 36722 41556 36728 41568
rect 36780 41556 36786 41608
rect 36906 41556 36912 41608
rect 36964 41556 36970 41608
rect 37458 41556 37464 41608
rect 37516 41556 37522 41608
rect 38654 41556 38660 41608
rect 38712 41556 38718 41608
rect 42150 41556 42156 41608
rect 42208 41596 42214 41608
rect 43530 41596 43536 41608
rect 42208 41568 43536 41596
rect 42208 41556 42214 41568
rect 43530 41556 43536 41568
rect 43588 41556 43594 41608
rect 29978 41531 30036 41537
rect 29978 41528 29990 41531
rect 28920 41500 29990 41528
rect 25056 41432 26234 41460
rect 26421 41463 26479 41469
rect 26421 41429 26433 41463
rect 26467 41460 26479 41463
rect 26694 41460 26700 41472
rect 26467 41432 26700 41460
rect 26467 41429 26479 41432
rect 26421 41423 26479 41429
rect 26694 41420 26700 41432
rect 26752 41420 26758 41472
rect 28258 41420 28264 41472
rect 28316 41420 28322 41472
rect 28920 41469 28948 41500
rect 29978 41497 29990 41500
rect 30024 41497 30036 41531
rect 29978 41491 30036 41497
rect 33502 41488 33508 41540
rect 33560 41488 33566 41540
rect 33870 41488 33876 41540
rect 33928 41528 33934 41540
rect 40586 41528 40592 41540
rect 33928 41500 40592 41528
rect 33928 41488 33934 41500
rect 40586 41488 40592 41500
rect 40644 41528 40650 41540
rect 43070 41528 43076 41540
rect 40644 41500 43076 41528
rect 40644 41488 40650 41500
rect 43070 41488 43076 41500
rect 43128 41488 43134 41540
rect 28905 41463 28963 41469
rect 28905 41429 28917 41463
rect 28951 41429 28963 41463
rect 28905 41423 28963 41429
rect 30926 41420 30932 41472
rect 30984 41460 30990 41472
rect 31113 41463 31171 41469
rect 31113 41460 31125 41463
rect 30984 41432 31125 41460
rect 30984 41420 30990 41432
rect 31113 41429 31125 41432
rect 31159 41429 31171 41463
rect 31113 41423 31171 41429
rect 31846 41420 31852 41472
rect 31904 41460 31910 41472
rect 32490 41460 32496 41472
rect 31904 41432 32496 41460
rect 31904 41420 31910 41432
rect 32490 41420 32496 41432
rect 32548 41460 32554 41472
rect 32953 41463 33011 41469
rect 32953 41460 32965 41463
rect 32548 41432 32965 41460
rect 32548 41420 32554 41432
rect 32953 41429 32965 41432
rect 32999 41429 33011 41463
rect 32953 41423 33011 41429
rect 34698 41420 34704 41472
rect 34756 41460 34762 41472
rect 34885 41463 34943 41469
rect 34885 41460 34897 41463
rect 34756 41432 34897 41460
rect 34756 41420 34762 41432
rect 34885 41429 34897 41432
rect 34931 41429 34943 41463
rect 34885 41423 34943 41429
rect 36262 41420 36268 41472
rect 36320 41460 36326 41472
rect 36725 41463 36783 41469
rect 36725 41460 36737 41463
rect 36320 41432 36737 41460
rect 36320 41420 36326 41432
rect 36725 41429 36737 41432
rect 36771 41429 36783 41463
rect 36725 41423 36783 41429
rect 37645 41463 37703 41469
rect 37645 41429 37657 41463
rect 37691 41460 37703 41463
rect 37734 41460 37740 41472
rect 37691 41432 37740 41460
rect 37691 41429 37703 41432
rect 37645 41423 37703 41429
rect 37734 41420 37740 41432
rect 37792 41420 37798 41472
rect 38197 41463 38255 41469
rect 38197 41429 38209 41463
rect 38243 41460 38255 41463
rect 38378 41460 38384 41472
rect 38243 41432 38384 41460
rect 38243 41429 38255 41432
rect 38197 41423 38255 41429
rect 38378 41420 38384 41432
rect 38436 41420 38442 41472
rect 39298 41420 39304 41472
rect 39356 41420 39362 41472
rect 39666 41420 39672 41472
rect 39724 41460 39730 41472
rect 40310 41460 40316 41472
rect 39724 41432 40316 41460
rect 39724 41420 39730 41432
rect 40310 41420 40316 41432
rect 40368 41420 40374 41472
rect 40402 41420 40408 41472
rect 40460 41420 40466 41472
rect 40773 41463 40831 41469
rect 40773 41429 40785 41463
rect 40819 41460 40831 41463
rect 41138 41460 41144 41472
rect 40819 41432 41144 41460
rect 40819 41429 40831 41432
rect 40773 41423 40831 41429
rect 41138 41420 41144 41432
rect 41196 41420 41202 41472
rect 41230 41420 41236 41472
rect 41288 41420 41294 41472
rect 42610 41420 42616 41472
rect 42668 41420 42674 41472
rect 42886 41420 42892 41472
rect 42944 41460 42950 41472
rect 43165 41463 43223 41469
rect 43165 41460 43177 41463
rect 42944 41432 43177 41460
rect 42944 41420 42950 41432
rect 43165 41429 43177 41432
rect 43211 41429 43223 41463
rect 43165 41423 43223 41429
rect 1104 41370 43884 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 43884 41370
rect 1104 41296 43884 41318
rect 19705 41259 19763 41265
rect 19705 41225 19717 41259
rect 19751 41256 19763 41259
rect 21450 41256 21456 41268
rect 19751 41228 21456 41256
rect 19751 41225 19763 41228
rect 19705 41219 19763 41225
rect 21450 41216 21456 41228
rect 21508 41216 21514 41268
rect 22738 41216 22744 41268
rect 22796 41256 22802 41268
rect 22833 41259 22891 41265
rect 22833 41256 22845 41259
rect 22796 41228 22845 41256
rect 22796 41216 22802 41228
rect 22833 41225 22845 41228
rect 22879 41225 22891 41259
rect 22833 41219 22891 41225
rect 25317 41259 25375 41265
rect 25317 41225 25329 41259
rect 25363 41256 25375 41259
rect 25406 41256 25412 41268
rect 25363 41228 25412 41256
rect 25363 41225 25375 41228
rect 25317 41219 25375 41225
rect 25406 41216 25412 41228
rect 25464 41216 25470 41268
rect 27157 41259 27215 41265
rect 27157 41225 27169 41259
rect 27203 41256 27215 41259
rect 27338 41256 27344 41268
rect 27203 41228 27344 41256
rect 27203 41225 27215 41228
rect 27157 41219 27215 41225
rect 27338 41216 27344 41228
rect 27396 41216 27402 41268
rect 27525 41259 27583 41265
rect 27525 41225 27537 41259
rect 27571 41256 27583 41259
rect 28258 41256 28264 41268
rect 27571 41228 28264 41256
rect 27571 41225 27583 41228
rect 27525 41219 27583 41225
rect 28258 41216 28264 41228
rect 28316 41216 28322 41268
rect 29086 41216 29092 41268
rect 29144 41216 29150 41268
rect 30650 41216 30656 41268
rect 30708 41216 30714 41268
rect 32858 41216 32864 41268
rect 32916 41256 32922 41268
rect 33689 41259 33747 41265
rect 33689 41256 33701 41259
rect 32916 41228 33701 41256
rect 32916 41216 32922 41228
rect 33689 41225 33701 41228
rect 33735 41225 33747 41259
rect 33689 41219 33747 41225
rect 34790 41216 34796 41268
rect 34848 41256 34854 41268
rect 35069 41259 35127 41265
rect 35069 41256 35081 41259
rect 34848 41228 35081 41256
rect 34848 41216 34854 41228
rect 35069 41225 35081 41228
rect 35115 41225 35127 41259
rect 35069 41219 35127 41225
rect 39942 41216 39948 41268
rect 40000 41256 40006 41268
rect 40681 41259 40739 41265
rect 40681 41256 40693 41259
rect 40000 41228 40693 41256
rect 40000 41216 40006 41228
rect 40681 41225 40693 41228
rect 40727 41256 40739 41259
rect 42886 41256 42892 41268
rect 40727 41228 42892 41256
rect 40727 41225 40739 41228
rect 40681 41219 40739 41225
rect 42886 41216 42892 41228
rect 42944 41216 42950 41268
rect 43070 41216 43076 41268
rect 43128 41256 43134 41268
rect 43165 41259 43223 41265
rect 43165 41256 43177 41259
rect 43128 41228 43177 41256
rect 43128 41216 43134 41228
rect 43165 41225 43177 41228
rect 43211 41225 43223 41259
rect 43165 41219 43223 41225
rect 21085 41191 21143 41197
rect 21085 41157 21097 41191
rect 21131 41188 21143 41191
rect 21358 41188 21364 41200
rect 21131 41160 21364 41188
rect 21131 41157 21143 41160
rect 21085 41151 21143 41157
rect 21358 41148 21364 41160
rect 21416 41188 21422 41200
rect 21542 41188 21548 41200
rect 21416 41160 21548 41188
rect 21416 41148 21422 41160
rect 21542 41148 21548 41160
rect 21600 41148 21606 41200
rect 31021 41191 31079 41197
rect 31021 41157 31033 41191
rect 31067 41188 31079 41191
rect 31846 41188 31852 41200
rect 31067 41160 31852 41188
rect 31067 41157 31079 41160
rect 31021 41151 31079 41157
rect 31846 41148 31852 41160
rect 31904 41148 31910 41200
rect 39298 41188 39304 41200
rect 32324 41160 39304 41188
rect 21177 41123 21235 41129
rect 21177 41089 21189 41123
rect 21223 41120 21235 41123
rect 21634 41120 21640 41132
rect 21223 41092 21640 41120
rect 21223 41089 21235 41092
rect 21177 41083 21235 41089
rect 21634 41080 21640 41092
rect 21692 41120 21698 41132
rect 21818 41120 21824 41132
rect 21692 41092 21824 41120
rect 21692 41080 21698 41092
rect 21818 41080 21824 41092
rect 21876 41080 21882 41132
rect 23201 41123 23259 41129
rect 23201 41089 23213 41123
rect 23247 41120 23259 41123
rect 24118 41120 24124 41132
rect 23247 41092 24124 41120
rect 23247 41089 23259 41092
rect 23201 41083 23259 41089
rect 24118 41080 24124 41092
rect 24176 41080 24182 41132
rect 25685 41123 25743 41129
rect 25685 41089 25697 41123
rect 25731 41120 25743 41123
rect 26694 41120 26700 41132
rect 25731 41092 26700 41120
rect 25731 41089 25743 41092
rect 25685 41083 25743 41089
rect 26694 41080 26700 41092
rect 26752 41080 26758 41132
rect 27890 41080 27896 41132
rect 27948 41120 27954 41132
rect 28721 41123 28779 41129
rect 27948 41092 28580 41120
rect 27948 41080 27954 41092
rect 28552 41064 28580 41092
rect 28721 41089 28733 41123
rect 28767 41120 28779 41123
rect 30466 41120 30472 41132
rect 28767 41092 30472 41120
rect 28767 41089 28779 41092
rect 28721 41083 28779 41089
rect 30466 41080 30472 41092
rect 30524 41120 30530 41132
rect 30926 41120 30932 41132
rect 30524 41092 30932 41120
rect 30524 41080 30530 41092
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 31662 41080 31668 41132
rect 31720 41120 31726 41132
rect 32324 41129 32352 41160
rect 39298 41148 39304 41160
rect 39356 41148 39362 41200
rect 39390 41148 39396 41200
rect 39448 41188 39454 41200
rect 39546 41191 39604 41197
rect 39546 41188 39558 41191
rect 39448 41160 39558 41188
rect 39448 41148 39454 41160
rect 39546 41157 39558 41160
rect 39592 41157 39604 41191
rect 39546 41151 39604 41157
rect 32582 41129 32588 41132
rect 32309 41123 32367 41129
rect 32309 41120 32321 41123
rect 31720 41092 32321 41120
rect 31720 41080 31726 41092
rect 32309 41089 32321 41092
rect 32355 41089 32367 41123
rect 32576 41120 32588 41129
rect 32543 41092 32588 41120
rect 32309 41083 32367 41089
rect 32576 41083 32588 41092
rect 32582 41080 32588 41083
rect 32640 41080 32646 41132
rect 34698 41080 34704 41132
rect 34756 41080 34762 41132
rect 35796 41123 35854 41129
rect 35796 41089 35808 41123
rect 35842 41120 35854 41123
rect 36262 41120 36268 41132
rect 35842 41092 36268 41120
rect 35842 41089 35854 41092
rect 35796 41083 35854 41089
rect 36262 41080 36268 41092
rect 36320 41080 36326 41132
rect 37734 41129 37740 41132
rect 37728 41120 37740 41129
rect 37695 41092 37740 41120
rect 37728 41083 37740 41092
rect 37734 41080 37740 41083
rect 37792 41080 37798 41132
rect 41138 41080 41144 41132
rect 41196 41080 41202 41132
rect 18874 41012 18880 41064
rect 18932 41052 18938 41064
rect 20257 41055 20315 41061
rect 20257 41052 20269 41055
rect 18932 41024 20269 41052
rect 18932 41012 18938 41024
rect 20257 41021 20269 41024
rect 20303 41052 20315 41055
rect 21361 41055 21419 41061
rect 21361 41052 21373 41055
rect 20303 41024 21373 41052
rect 20303 41021 20315 41024
rect 20257 41015 20315 41021
rect 21361 41021 21373 41024
rect 21407 41052 21419 41055
rect 21407 41024 22094 41052
rect 21407 41021 21419 41024
rect 21361 41015 21419 41021
rect 22066 40996 22094 41024
rect 23290 41012 23296 41064
rect 23348 41012 23354 41064
rect 23382 41012 23388 41064
rect 23440 41052 23446 41064
rect 23477 41055 23535 41061
rect 23477 41052 23489 41055
rect 23440 41024 23489 41052
rect 23440 41012 23446 41024
rect 23477 41021 23489 41024
rect 23523 41021 23535 41055
rect 23477 41015 23535 41021
rect 20714 40944 20720 40996
rect 20772 40944 20778 40996
rect 22066 40956 22100 40996
rect 22094 40944 22100 40956
rect 22152 40984 22158 40996
rect 23492 40984 23520 41015
rect 24854 41012 24860 41064
rect 24912 41052 24918 41064
rect 25774 41052 25780 41064
rect 24912 41024 25780 41052
rect 24912 41012 24918 41024
rect 25774 41012 25780 41024
rect 25832 41012 25838 41064
rect 25961 41055 26019 41061
rect 25961 41021 25973 41055
rect 26007 41021 26019 41055
rect 25961 41015 26019 41021
rect 24121 40987 24179 40993
rect 24121 40984 24133 40987
rect 22152 40956 24133 40984
rect 22152 40944 22158 40956
rect 24121 40953 24133 40956
rect 24167 40984 24179 40987
rect 25976 40984 26004 41015
rect 26326 41012 26332 41064
rect 26384 41052 26390 41064
rect 27614 41052 27620 41064
rect 26384 41024 27620 41052
rect 26384 41012 26390 41024
rect 27614 41012 27620 41024
rect 27672 41012 27678 41064
rect 27801 41055 27859 41061
rect 27801 41021 27813 41055
rect 27847 41052 27859 41055
rect 28445 41055 28503 41061
rect 28445 41052 28457 41055
rect 27847 41024 28457 41052
rect 27847 41021 27859 41024
rect 27801 41015 27859 41021
rect 28445 41021 28457 41024
rect 28491 41021 28503 41055
rect 28445 41015 28503 41021
rect 27816 40984 27844 41015
rect 24167 40956 27844 40984
rect 28460 40984 28488 41015
rect 28534 41012 28540 41064
rect 28592 41052 28598 41064
rect 28629 41055 28687 41061
rect 28629 41052 28641 41055
rect 28592 41024 28641 41052
rect 28592 41012 28598 41024
rect 28629 41021 28641 41024
rect 28675 41021 28687 41055
rect 28629 41015 28687 41021
rect 29641 41055 29699 41061
rect 29641 41021 29653 41055
rect 29687 41052 29699 41055
rect 30282 41052 30288 41064
rect 29687 41024 30288 41052
rect 29687 41021 29699 41024
rect 29641 41015 29699 41021
rect 30282 41012 30288 41024
rect 30340 41012 30346 41064
rect 31110 41012 31116 41064
rect 31168 41012 31174 41064
rect 31297 41055 31355 41061
rect 31297 41021 31309 41055
rect 31343 41052 31355 41055
rect 31343 41024 31616 41052
rect 31343 41021 31355 41024
rect 31297 41015 31355 41021
rect 31312 40984 31340 41015
rect 28460 40956 31340 40984
rect 24167 40953 24179 40956
rect 24121 40947 24179 40953
rect 31588 40928 31616 41024
rect 33502 41012 33508 41064
rect 33560 41052 33566 41064
rect 34422 41052 34428 41064
rect 33560 41024 34428 41052
rect 33560 41012 33566 41024
rect 34422 41012 34428 41024
rect 34480 41012 34486 41064
rect 34606 41012 34612 41064
rect 34664 41052 34670 41064
rect 34790 41052 34796 41064
rect 34664 41024 34796 41052
rect 34664 41012 34670 41024
rect 34790 41012 34796 41024
rect 34848 41012 34854 41064
rect 35529 41055 35587 41061
rect 35529 41021 35541 41055
rect 35575 41021 35587 41055
rect 37461 41055 37519 41061
rect 37461 41052 37473 41055
rect 35529 41015 35587 41021
rect 36556 41024 37473 41052
rect 33870 40984 33876 40996
rect 33244 40956 33876 40984
rect 22373 40919 22431 40925
rect 22373 40885 22385 40919
rect 22419 40916 22431 40919
rect 22646 40916 22652 40928
rect 22419 40888 22652 40916
rect 22419 40885 22431 40888
rect 22373 40879 22431 40885
rect 22646 40876 22652 40888
rect 22704 40876 22710 40928
rect 24857 40919 24915 40925
rect 24857 40885 24869 40919
rect 24903 40916 24915 40919
rect 25222 40916 25228 40928
rect 24903 40888 25228 40916
rect 24903 40885 24915 40888
rect 24857 40879 24915 40885
rect 25222 40876 25228 40888
rect 25280 40876 25286 40928
rect 26602 40876 26608 40928
rect 26660 40916 26666 40928
rect 26970 40916 26976 40928
rect 26660 40888 26976 40916
rect 26660 40876 26666 40888
rect 26970 40876 26976 40888
rect 27028 40876 27034 40928
rect 30098 40876 30104 40928
rect 30156 40876 30162 40928
rect 31570 40876 31576 40928
rect 31628 40916 31634 40928
rect 33244 40916 33272 40956
rect 33870 40944 33876 40956
rect 33928 40944 33934 40996
rect 34054 40944 34060 40996
rect 34112 40984 34118 40996
rect 35544 40984 35572 41015
rect 34112 40956 35572 40984
rect 34112 40944 34118 40956
rect 31628 40888 33272 40916
rect 35544 40916 35572 40956
rect 36556 40916 36584 41024
rect 37461 41021 37473 41024
rect 37507 41021 37519 41055
rect 37461 41015 37519 41021
rect 35544 40888 36584 40916
rect 36909 40919 36967 40925
rect 31628 40876 31634 40888
rect 36909 40885 36921 40919
rect 36955 40916 36967 40919
rect 36998 40916 37004 40928
rect 36955 40888 37004 40916
rect 36955 40885 36967 40888
rect 36909 40879 36967 40885
rect 36998 40876 37004 40888
rect 37056 40876 37062 40928
rect 37476 40916 37504 41015
rect 38838 41012 38844 41064
rect 38896 41052 38902 41064
rect 39301 41055 39359 41061
rect 39301 41052 39313 41055
rect 38896 41024 39313 41052
rect 38896 41012 38902 41024
rect 39301 41021 39313 41024
rect 39347 41021 39359 41055
rect 39301 41015 39359 41021
rect 41414 40984 41420 40996
rect 38396 40956 39344 40984
rect 38396 40916 38424 40956
rect 37476 40888 38424 40916
rect 38746 40876 38752 40928
rect 38804 40916 38810 40928
rect 38841 40919 38899 40925
rect 38841 40916 38853 40919
rect 38804 40888 38853 40916
rect 38804 40876 38810 40888
rect 38841 40885 38853 40888
rect 38887 40885 38899 40919
rect 39316 40916 39344 40956
rect 40236 40956 41420 40984
rect 40236 40916 40264 40956
rect 41414 40944 41420 40956
rect 41472 40944 41478 40996
rect 39316 40888 40264 40916
rect 38841 40879 38899 40885
rect 41322 40876 41328 40928
rect 41380 40876 41386 40928
rect 41782 40876 41788 40928
rect 41840 40876 41846 40928
rect 42610 40876 42616 40928
rect 42668 40876 42674 40928
rect 1104 40826 43884 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 43884 40826
rect 1104 40752 43884 40774
rect 19981 40715 20039 40721
rect 19981 40681 19993 40715
rect 20027 40712 20039 40715
rect 24302 40712 24308 40724
rect 20027 40684 24308 40712
rect 20027 40681 20039 40684
rect 19981 40675 20039 40681
rect 24302 40672 24308 40684
rect 24360 40672 24366 40724
rect 32217 40715 32275 40721
rect 32217 40681 32229 40715
rect 32263 40712 32275 40715
rect 32306 40712 32312 40724
rect 32263 40684 32312 40712
rect 32263 40681 32275 40684
rect 32217 40675 32275 40681
rect 32306 40672 32312 40684
rect 32364 40672 32370 40724
rect 34238 40712 34244 40724
rect 32968 40684 34244 40712
rect 30282 40604 30288 40656
rect 30340 40644 30346 40656
rect 32968 40644 32996 40684
rect 34238 40672 34244 40684
rect 34296 40672 34302 40724
rect 34422 40672 34428 40724
rect 34480 40712 34486 40724
rect 35529 40715 35587 40721
rect 35529 40712 35541 40715
rect 34480 40684 35541 40712
rect 34480 40672 34486 40684
rect 35529 40681 35541 40684
rect 35575 40681 35587 40715
rect 35529 40675 35587 40681
rect 30340 40616 32996 40644
rect 30340 40604 30346 40616
rect 20717 40579 20775 40585
rect 20717 40545 20729 40579
rect 20763 40576 20775 40579
rect 22922 40576 22928 40588
rect 20763 40548 22928 40576
rect 20763 40545 20775 40548
rect 20717 40539 20775 40545
rect 22922 40536 22928 40548
rect 22980 40536 22986 40588
rect 24029 40579 24087 40585
rect 24029 40545 24041 40579
rect 24075 40576 24087 40579
rect 24946 40576 24952 40588
rect 24075 40548 24952 40576
rect 24075 40545 24087 40548
rect 24029 40539 24087 40545
rect 24946 40536 24952 40548
rect 25004 40536 25010 40588
rect 31570 40536 31576 40588
rect 31628 40536 31634 40588
rect 35544 40576 35572 40675
rect 36906 40672 36912 40724
rect 36964 40672 36970 40724
rect 37369 40715 37427 40721
rect 37369 40681 37381 40715
rect 37415 40712 37427 40715
rect 37458 40712 37464 40724
rect 37415 40684 37464 40712
rect 37415 40681 37427 40684
rect 37369 40675 37427 40681
rect 37458 40672 37464 40684
rect 37516 40672 37522 40724
rect 38565 40715 38623 40721
rect 38565 40681 38577 40715
rect 38611 40712 38623 40715
rect 38654 40712 38660 40724
rect 38611 40684 38660 40712
rect 38611 40681 38623 40684
rect 38565 40675 38623 40681
rect 38654 40672 38660 40684
rect 38712 40672 38718 40724
rect 40037 40715 40095 40721
rect 40037 40681 40049 40715
rect 40083 40712 40095 40715
rect 40402 40712 40408 40724
rect 40083 40684 40408 40712
rect 40083 40681 40095 40684
rect 40037 40675 40095 40681
rect 38028 40616 38332 40644
rect 38028 40585 38056 40616
rect 36265 40579 36323 40585
rect 36265 40576 36277 40579
rect 35544 40548 36277 40576
rect 36265 40545 36277 40548
rect 36311 40576 36323 40579
rect 38013 40579 38071 40585
rect 38013 40576 38025 40579
rect 36311 40548 38025 40576
rect 36311 40545 36323 40548
rect 36265 40539 36323 40545
rect 38013 40545 38025 40548
rect 38059 40545 38071 40579
rect 38304 40576 38332 40616
rect 38378 40604 38384 40656
rect 38436 40644 38442 40656
rect 40052 40644 40080 40675
rect 40402 40672 40408 40684
rect 40460 40672 40466 40724
rect 38436 40616 40080 40644
rect 38436 40604 38442 40616
rect 39209 40579 39267 40585
rect 39209 40576 39221 40579
rect 38304 40548 39221 40576
rect 38013 40539 38071 40545
rect 39209 40545 39221 40548
rect 39255 40576 39267 40579
rect 40126 40576 40132 40588
rect 39255 40548 40132 40576
rect 39255 40545 39267 40548
rect 39209 40539 39267 40545
rect 40126 40536 40132 40548
rect 40184 40536 40190 40588
rect 20622 40468 20628 40520
rect 20680 40468 20686 40520
rect 25038 40468 25044 40520
rect 25096 40508 25102 40520
rect 25096 40480 26004 40508
rect 25096 40468 25102 40480
rect 25976 40452 26004 40480
rect 27706 40468 27712 40520
rect 27764 40508 27770 40520
rect 30837 40511 30895 40517
rect 30837 40508 30849 40511
rect 27764 40480 30849 40508
rect 27764 40468 27770 40480
rect 30837 40477 30849 40480
rect 30883 40508 30895 40511
rect 31478 40508 31484 40520
rect 30883 40480 31484 40508
rect 30883 40477 30895 40480
rect 30837 40471 30895 40477
rect 31478 40468 31484 40480
rect 31536 40468 31542 40520
rect 31849 40511 31907 40517
rect 31849 40477 31861 40511
rect 31895 40508 31907 40511
rect 32858 40508 32864 40520
rect 31895 40480 32864 40508
rect 31895 40477 31907 40480
rect 31849 40471 31907 40477
rect 32858 40468 32864 40480
rect 32916 40468 32922 40520
rect 34054 40468 34060 40520
rect 34112 40468 34118 40520
rect 35710 40468 35716 40520
rect 35768 40468 35774 40520
rect 36541 40511 36599 40517
rect 36541 40477 36553 40511
rect 36587 40508 36599 40511
rect 36998 40508 37004 40520
rect 36587 40480 37004 40508
rect 36587 40477 36599 40480
rect 36541 40471 36599 40477
rect 36998 40468 37004 40480
rect 37056 40508 37062 40520
rect 37734 40508 37740 40520
rect 37056 40480 37740 40508
rect 37056 40468 37062 40480
rect 37734 40468 37740 40480
rect 37792 40468 37798 40520
rect 37918 40468 37924 40520
rect 37976 40508 37982 40520
rect 41161 40511 41219 40517
rect 37976 40480 40080 40508
rect 37976 40468 37982 40480
rect 23566 40400 23572 40452
rect 23624 40440 23630 40452
rect 23762 40443 23820 40449
rect 23762 40440 23774 40443
rect 23624 40412 23774 40440
rect 23624 40400 23630 40412
rect 23762 40409 23774 40412
rect 23808 40409 23820 40443
rect 23762 40403 23820 40409
rect 24854 40400 24860 40452
rect 24912 40440 24918 40452
rect 25286 40443 25344 40449
rect 25286 40440 25298 40443
rect 24912 40412 25298 40440
rect 24912 40400 24918 40412
rect 25286 40409 25298 40412
rect 25332 40409 25344 40443
rect 25286 40403 25344 40409
rect 25958 40400 25964 40452
rect 26016 40400 26022 40452
rect 26234 40400 26240 40452
rect 26292 40440 26298 40452
rect 26881 40443 26939 40449
rect 26881 40440 26893 40443
rect 26292 40412 26893 40440
rect 26292 40400 26298 40412
rect 26881 40409 26893 40412
rect 26927 40409 26939 40443
rect 26881 40403 26939 40409
rect 28350 40400 28356 40452
rect 28408 40440 28414 40452
rect 28721 40443 28779 40449
rect 28721 40440 28733 40443
rect 28408 40412 28733 40440
rect 28408 40400 28414 40412
rect 28721 40409 28733 40412
rect 28767 40409 28779 40443
rect 28721 40403 28779 40409
rect 28902 40400 28908 40452
rect 28960 40400 28966 40452
rect 29089 40443 29147 40449
rect 29089 40409 29101 40443
rect 29135 40440 29147 40443
rect 30650 40440 30656 40452
rect 29135 40412 30656 40440
rect 29135 40409 29147 40412
rect 29089 40403 29147 40409
rect 30650 40400 30656 40412
rect 30708 40400 30714 40452
rect 31754 40400 31760 40452
rect 31812 40440 31818 40452
rect 32766 40440 32772 40452
rect 31812 40412 32772 40440
rect 31812 40400 31818 40412
rect 32766 40400 32772 40412
rect 32824 40400 32830 40452
rect 33134 40400 33140 40452
rect 33192 40440 33198 40452
rect 33812 40443 33870 40449
rect 33192 40412 33364 40440
rect 33192 40400 33198 40412
rect 18782 40332 18788 40384
rect 18840 40332 18846 40384
rect 20993 40375 21051 40381
rect 20993 40341 21005 40375
rect 21039 40372 21051 40375
rect 21082 40372 21088 40384
rect 21039 40344 21088 40372
rect 21039 40341 21051 40344
rect 20993 40335 21051 40341
rect 21082 40332 21088 40344
rect 21140 40332 21146 40384
rect 21266 40332 21272 40384
rect 21324 40372 21330 40384
rect 21453 40375 21511 40381
rect 21453 40372 21465 40375
rect 21324 40344 21465 40372
rect 21324 40332 21330 40344
rect 21453 40341 21465 40344
rect 21499 40341 21511 40375
rect 21453 40335 21511 40341
rect 22189 40375 22247 40381
rect 22189 40341 22201 40375
rect 22235 40372 22247 40375
rect 22554 40372 22560 40384
rect 22235 40344 22560 40372
rect 22235 40341 22247 40344
rect 22189 40335 22247 40341
rect 22554 40332 22560 40344
rect 22612 40332 22618 40384
rect 22649 40375 22707 40381
rect 22649 40341 22661 40375
rect 22695 40372 22707 40375
rect 22738 40372 22744 40384
rect 22695 40344 22744 40372
rect 22695 40341 22707 40344
rect 22649 40335 22707 40341
rect 22738 40332 22744 40344
rect 22796 40332 22802 40384
rect 26326 40332 26332 40384
rect 26384 40372 26390 40384
rect 26421 40375 26479 40381
rect 26421 40372 26433 40375
rect 26384 40344 26433 40372
rect 26384 40332 26390 40344
rect 26421 40341 26433 40344
rect 26467 40341 26479 40375
rect 26421 40335 26479 40341
rect 27801 40375 27859 40381
rect 27801 40341 27813 40375
rect 27847 40372 27859 40375
rect 27890 40372 27896 40384
rect 27847 40344 27896 40372
rect 27847 40341 27859 40344
rect 27801 40335 27859 40341
rect 27890 40332 27896 40344
rect 27948 40332 27954 40384
rect 29822 40332 29828 40384
rect 29880 40332 29886 40384
rect 30374 40332 30380 40384
rect 30432 40332 30438 40384
rect 32677 40375 32735 40381
rect 32677 40341 32689 40375
rect 32723 40372 32735 40375
rect 33226 40372 33232 40384
rect 32723 40344 33232 40372
rect 32723 40341 32735 40344
rect 32677 40335 32735 40341
rect 33226 40332 33232 40344
rect 33284 40332 33290 40384
rect 33336 40372 33364 40412
rect 33812 40409 33824 40443
rect 33858 40440 33870 40443
rect 33962 40440 33968 40452
rect 33858 40412 33968 40440
rect 33858 40409 33870 40412
rect 33812 40403 33870 40409
rect 33962 40400 33968 40412
rect 34020 40400 34026 40452
rect 34330 40400 34336 40452
rect 34388 40440 34394 40452
rect 34977 40443 35035 40449
rect 34977 40440 34989 40443
rect 34388 40412 34989 40440
rect 34388 40400 34394 40412
rect 34977 40409 34989 40412
rect 35023 40440 35035 40443
rect 37182 40440 37188 40452
rect 35023 40412 37188 40440
rect 35023 40409 35035 40412
rect 34977 40403 35035 40409
rect 37182 40400 37188 40412
rect 37240 40400 37246 40452
rect 37458 40400 37464 40452
rect 37516 40440 37522 40452
rect 37829 40443 37887 40449
rect 37829 40440 37841 40443
rect 37516 40412 37841 40440
rect 37516 40400 37522 40412
rect 37829 40409 37841 40412
rect 37875 40409 37887 40443
rect 39942 40440 39948 40452
rect 37829 40403 37887 40409
rect 38948 40412 39948 40440
rect 34348 40372 34376 40400
rect 38948 40384 38976 40412
rect 39942 40400 39948 40412
rect 40000 40400 40006 40452
rect 33336 40344 34376 40372
rect 35894 40332 35900 40384
rect 35952 40372 35958 40384
rect 36446 40372 36452 40384
rect 35952 40344 36452 40372
rect 35952 40332 35958 40344
rect 36446 40332 36452 40344
rect 36504 40332 36510 40384
rect 37737 40375 37795 40381
rect 37737 40341 37749 40375
rect 37783 40372 37795 40375
rect 38746 40372 38752 40384
rect 37783 40344 38752 40372
rect 37783 40341 37795 40344
rect 37737 40335 37795 40341
rect 38746 40332 38752 40344
rect 38804 40332 38810 40384
rect 38930 40332 38936 40384
rect 38988 40332 38994 40384
rect 39022 40332 39028 40384
rect 39080 40372 39086 40384
rect 39482 40372 39488 40384
rect 39080 40344 39488 40372
rect 39080 40332 39086 40344
rect 39482 40332 39488 40344
rect 39540 40332 39546 40384
rect 40052 40372 40080 40480
rect 41161 40477 41173 40511
rect 41207 40508 41219 40511
rect 41322 40508 41328 40520
rect 41207 40480 41328 40508
rect 41207 40477 41219 40480
rect 41161 40471 41219 40477
rect 41322 40468 41328 40480
rect 41380 40468 41386 40520
rect 41414 40468 41420 40520
rect 41472 40508 41478 40520
rect 41874 40508 41880 40520
rect 41472 40480 41880 40508
rect 41472 40468 41478 40480
rect 41874 40468 41880 40480
rect 41932 40468 41938 40520
rect 42610 40440 42616 40452
rect 41386 40412 42616 40440
rect 41386 40372 41414 40412
rect 42610 40400 42616 40412
rect 42668 40400 42674 40452
rect 40052 40344 41414 40372
rect 41598 40332 41604 40384
rect 41656 40372 41662 40384
rect 41877 40375 41935 40381
rect 41877 40372 41889 40375
rect 41656 40344 41889 40372
rect 41656 40332 41662 40344
rect 41877 40341 41889 40344
rect 41923 40341 41935 40375
rect 41877 40335 41935 40341
rect 42334 40332 42340 40384
rect 42392 40372 42398 40384
rect 42429 40375 42487 40381
rect 42429 40372 42441 40375
rect 42392 40344 42441 40372
rect 42392 40332 42398 40344
rect 42429 40341 42441 40344
rect 42475 40341 42487 40375
rect 42429 40335 42487 40341
rect 42886 40332 42892 40384
rect 42944 40372 42950 40384
rect 42981 40375 43039 40381
rect 42981 40372 42993 40375
rect 42944 40344 42993 40372
rect 42944 40332 42950 40344
rect 42981 40341 42993 40344
rect 43027 40341 43039 40375
rect 42981 40335 43039 40341
rect 1104 40282 43884 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 43884 40282
rect 1104 40208 43884 40230
rect 21453 40171 21511 40177
rect 19352 40140 20760 40168
rect 9122 40060 9128 40112
rect 9180 40100 9186 40112
rect 9674 40100 9680 40112
rect 9180 40072 9680 40100
rect 9180 40060 9186 40072
rect 9674 40060 9680 40072
rect 9732 40060 9738 40112
rect 16942 40060 16948 40112
rect 17000 40100 17006 40112
rect 19150 40100 19156 40112
rect 17000 40072 19156 40100
rect 17000 40060 17006 40072
rect 19150 40060 19156 40072
rect 19208 40060 19214 40112
rect 18322 39992 18328 40044
rect 18380 40032 18386 40044
rect 18969 40035 19027 40041
rect 18969 40032 18981 40035
rect 18380 40004 18981 40032
rect 18380 39992 18386 40004
rect 18969 40001 18981 40004
rect 19015 40032 19027 40035
rect 19352 40032 19380 40140
rect 20622 40100 20628 40112
rect 19444 40072 20628 40100
rect 19444 40041 19472 40072
rect 20622 40060 20628 40072
rect 20680 40060 20686 40112
rect 19015 40004 19380 40032
rect 19429 40035 19487 40041
rect 19015 40001 19027 40004
rect 18969 39995 19027 40001
rect 19429 40001 19441 40035
rect 19475 40001 19487 40035
rect 19429 39995 19487 40001
rect 19613 40035 19671 40041
rect 19613 40001 19625 40035
rect 19659 40032 19671 40035
rect 19886 40032 19892 40044
rect 19659 40004 19892 40032
rect 19659 40001 19671 40004
rect 19613 39995 19671 40001
rect 19886 39992 19892 40004
rect 19944 39992 19950 40044
rect 20329 40035 20387 40041
rect 20329 40032 20341 40035
rect 19996 40004 20341 40032
rect 19521 39967 19579 39973
rect 19521 39933 19533 39967
rect 19567 39964 19579 39967
rect 19996 39964 20024 40004
rect 20329 40001 20341 40004
rect 20375 40001 20387 40035
rect 20732 40032 20760 40140
rect 21453 40137 21465 40171
rect 21499 40168 21511 40171
rect 22370 40168 22376 40180
rect 21499 40140 22376 40168
rect 21499 40137 21511 40140
rect 21453 40131 21511 40137
rect 22370 40128 22376 40140
rect 22428 40128 22434 40180
rect 23106 40168 23112 40180
rect 22940 40140 23112 40168
rect 22646 40032 22652 40044
rect 20732 40004 22652 40032
rect 20329 39995 20387 40001
rect 22646 39992 22652 40004
rect 22704 39992 22710 40044
rect 22940 40041 22968 40140
rect 23106 40128 23112 40140
rect 23164 40168 23170 40180
rect 23164 40140 25544 40168
rect 23164 40128 23170 40140
rect 25038 40100 25044 40112
rect 24504 40072 25044 40100
rect 24504 40041 24532 40072
rect 25038 40060 25044 40072
rect 25096 40060 25102 40112
rect 25516 40109 25544 40140
rect 29178 40128 29184 40180
rect 29236 40168 29242 40180
rect 30098 40168 30104 40180
rect 29236 40140 30104 40168
rect 29236 40128 29242 40140
rect 30098 40128 30104 40140
rect 30156 40168 30162 40180
rect 30285 40171 30343 40177
rect 30285 40168 30297 40171
rect 30156 40140 30297 40168
rect 30156 40128 30162 40140
rect 30285 40137 30297 40140
rect 30331 40137 30343 40171
rect 30285 40131 30343 40137
rect 33597 40171 33655 40177
rect 33597 40137 33609 40171
rect 33643 40137 33655 40171
rect 33597 40131 33655 40137
rect 25317 40103 25375 40109
rect 25317 40100 25329 40103
rect 25148 40072 25329 40100
rect 22925 40035 22983 40041
rect 22925 40001 22937 40035
rect 22971 40001 22983 40035
rect 22925 39995 22983 40001
rect 24489 40035 24547 40041
rect 24489 40001 24501 40035
rect 24535 40001 24547 40035
rect 25148 40032 25176 40072
rect 25317 40069 25329 40072
rect 25363 40069 25375 40103
rect 25317 40063 25375 40069
rect 25501 40103 25559 40109
rect 25501 40069 25513 40103
rect 25547 40069 25559 40103
rect 25501 40063 25559 40069
rect 28644 40072 28856 40100
rect 27798 40032 27804 40044
rect 24489 39995 24547 40001
rect 24780 40004 25176 40032
rect 26804 40004 27804 40032
rect 19567 39936 20024 39964
rect 19567 39933 19579 39936
rect 19521 39927 19579 39933
rect 20070 39924 20076 39976
rect 20128 39924 20134 39976
rect 23017 39967 23075 39973
rect 23017 39933 23029 39967
rect 23063 39933 23075 39967
rect 23017 39927 23075 39933
rect 23293 39967 23351 39973
rect 23293 39933 23305 39967
rect 23339 39964 23351 39967
rect 23566 39964 23572 39976
rect 23339 39936 23572 39964
rect 23339 39933 23351 39936
rect 23293 39927 23351 39933
rect 20088 39828 20116 39924
rect 21174 39856 21180 39908
rect 21232 39896 21238 39908
rect 23032 39896 23060 39927
rect 23566 39924 23572 39936
rect 23624 39924 23630 39976
rect 23750 39924 23756 39976
rect 23808 39924 23814 39976
rect 24578 39924 24584 39976
rect 24636 39924 24642 39976
rect 24210 39896 24216 39908
rect 21232 39868 22968 39896
rect 23032 39868 24216 39896
rect 21232 39856 21238 39868
rect 20714 39828 20720 39840
rect 20088 39800 20720 39828
rect 20714 39788 20720 39800
rect 20772 39788 20778 39840
rect 22281 39831 22339 39837
rect 22281 39797 22293 39831
rect 22327 39828 22339 39831
rect 22646 39828 22652 39840
rect 22327 39800 22652 39828
rect 22327 39797 22339 39800
rect 22281 39791 22339 39797
rect 22646 39788 22652 39800
rect 22704 39788 22710 39840
rect 22940 39828 22968 39868
rect 24210 39856 24216 39868
rect 24268 39896 24274 39908
rect 24780 39896 24808 40004
rect 24854 39924 24860 39976
rect 24912 39924 24918 39976
rect 26804 39964 26832 40004
rect 27798 39992 27804 40004
rect 27856 40032 27862 40044
rect 28644 40032 28672 40072
rect 28718 40041 28724 40044
rect 27856 40004 28672 40032
rect 27856 39992 27862 40004
rect 28712 39995 28724 40041
rect 28718 39992 28724 39995
rect 28776 39992 28782 40044
rect 28828 40032 28856 40072
rect 30190 40060 30196 40112
rect 30248 40100 30254 40112
rect 30929 40103 30987 40109
rect 30929 40100 30941 40103
rect 30248 40072 30941 40100
rect 30248 40060 30254 40072
rect 30929 40069 30941 40072
rect 30975 40069 30987 40103
rect 30929 40063 30987 40069
rect 31113 40103 31171 40109
rect 31113 40069 31125 40103
rect 31159 40100 31171 40103
rect 31846 40100 31852 40112
rect 31159 40072 31852 40100
rect 31159 40069 31171 40072
rect 31113 40063 31171 40069
rect 31846 40060 31852 40072
rect 31904 40060 31910 40112
rect 33612 40100 33640 40131
rect 33962 40128 33968 40180
rect 34020 40168 34026 40180
rect 34057 40171 34115 40177
rect 34057 40168 34069 40171
rect 34020 40140 34069 40168
rect 34020 40128 34026 40140
rect 34057 40137 34069 40140
rect 34103 40137 34115 40171
rect 34057 40131 34115 40137
rect 34146 40128 34152 40180
rect 34204 40168 34210 40180
rect 35345 40171 35403 40177
rect 35345 40168 35357 40171
rect 34204 40140 35357 40168
rect 34204 40128 34210 40140
rect 35345 40137 35357 40140
rect 35391 40137 35403 40171
rect 35345 40131 35403 40137
rect 37090 40128 37096 40180
rect 37148 40168 37154 40180
rect 37918 40168 37924 40180
rect 37148 40140 37924 40168
rect 37148 40128 37154 40140
rect 37918 40128 37924 40140
rect 37976 40128 37982 40180
rect 41322 40128 41328 40180
rect 41380 40128 41386 40180
rect 33612 40072 34284 40100
rect 30374 40032 30380 40044
rect 28828 40004 30380 40032
rect 30374 39992 30380 40004
rect 30432 39992 30438 40044
rect 30837 40035 30895 40041
rect 30837 40001 30849 40035
rect 30883 40001 30895 40035
rect 30837 39995 30895 40001
rect 24964 39936 26832 39964
rect 24268 39868 24808 39896
rect 24268 39856 24274 39868
rect 24964 39828 24992 39936
rect 26878 39924 26884 39976
rect 26936 39964 26942 39976
rect 27154 39964 27160 39976
rect 26936 39936 27160 39964
rect 26936 39924 26942 39936
rect 27154 39924 27160 39936
rect 27212 39964 27218 39976
rect 28445 39967 28503 39973
rect 28445 39964 28457 39967
rect 27212 39936 28457 39964
rect 27212 39924 27218 39936
rect 28445 39933 28457 39936
rect 28491 39933 28503 39967
rect 30852 39964 30880 39995
rect 31018 39992 31024 40044
rect 31076 40032 31082 40044
rect 31573 40035 31631 40041
rect 31573 40032 31585 40035
rect 31076 40004 31585 40032
rect 31076 39992 31082 40004
rect 31573 40001 31585 40004
rect 31619 40001 31631 40035
rect 31573 39995 31631 40001
rect 31754 39992 31760 40044
rect 31812 39992 31818 40044
rect 32674 39992 32680 40044
rect 32732 40032 32738 40044
rect 33137 40035 33195 40041
rect 33137 40032 33149 40035
rect 32732 40004 33149 40032
rect 32732 39992 32738 40004
rect 33137 40001 33149 40004
rect 33183 40001 33195 40035
rect 33137 39995 33195 40001
rect 33226 39992 33232 40044
rect 33284 40032 33290 40044
rect 33778 40032 33784 40044
rect 33284 40004 33784 40032
rect 33284 39992 33290 40004
rect 33778 39992 33784 40004
rect 33836 39992 33842 40044
rect 34256 40041 34284 40072
rect 34241 40035 34299 40041
rect 34241 40001 34253 40035
rect 34287 40001 34299 40035
rect 34241 39995 34299 40001
rect 35434 39992 35440 40044
rect 35492 40032 35498 40044
rect 36458 40035 36516 40041
rect 36458 40032 36470 40035
rect 35492 40004 36470 40032
rect 35492 39992 35498 40004
rect 36458 40001 36470 40004
rect 36504 40001 36516 40035
rect 36458 39995 36516 40001
rect 36630 39992 36636 40044
rect 36688 40032 36694 40044
rect 38470 40032 38476 40044
rect 36688 40004 38476 40032
rect 36688 39992 36694 40004
rect 38470 39992 38476 40004
rect 38528 40032 38534 40044
rect 40865 40035 40923 40041
rect 40865 40032 40877 40035
rect 38528 40004 40877 40032
rect 38528 39992 38534 40004
rect 40865 40001 40877 40004
rect 40911 40032 40923 40035
rect 41877 40035 41935 40041
rect 41877 40032 41889 40035
rect 40911 40004 41889 40032
rect 40911 40001 40923 40004
rect 40865 39995 40923 40001
rect 41877 40001 41889 40004
rect 41923 40001 41935 40035
rect 41877 39995 41935 40001
rect 31386 39964 31392 39976
rect 30852 39936 31392 39964
rect 28445 39927 28503 39933
rect 31386 39924 31392 39936
rect 31444 39924 31450 39976
rect 33045 39967 33103 39973
rect 33045 39933 33057 39967
rect 33091 39964 33103 39967
rect 33502 39964 33508 39976
rect 33091 39936 33508 39964
rect 33091 39933 33103 39936
rect 33045 39927 33103 39933
rect 33502 39924 33508 39936
rect 33560 39924 33566 39976
rect 36722 39924 36728 39976
rect 36780 39964 36786 39976
rect 38838 39964 38844 39976
rect 36780 39936 38844 39964
rect 36780 39924 36786 39936
rect 38838 39924 38844 39936
rect 38896 39924 38902 39976
rect 41230 39964 41236 39976
rect 38948 39936 41236 39964
rect 32398 39856 32404 39908
rect 32456 39896 32462 39908
rect 38948 39896 38976 39936
rect 41230 39924 41236 39936
rect 41288 39924 41294 39976
rect 39669 39899 39727 39905
rect 39669 39896 39681 39899
rect 32456 39868 35112 39896
rect 32456 39856 32462 39868
rect 22940 39800 24992 39828
rect 25038 39788 25044 39840
rect 25096 39828 25102 39840
rect 25685 39831 25743 39837
rect 25685 39828 25697 39831
rect 25096 39800 25697 39828
rect 25096 39788 25102 39800
rect 25685 39797 25697 39800
rect 25731 39797 25743 39831
rect 25685 39791 25743 39797
rect 26237 39831 26295 39837
rect 26237 39797 26249 39831
rect 26283 39828 26295 39831
rect 27062 39828 27068 39840
rect 26283 39800 27068 39828
rect 26283 39797 26295 39800
rect 26237 39791 26295 39797
rect 27062 39788 27068 39800
rect 27120 39788 27126 39840
rect 27249 39831 27307 39837
rect 27249 39797 27261 39831
rect 27295 39828 27307 39831
rect 27522 39828 27528 39840
rect 27295 39800 27528 39828
rect 27295 39797 27307 39800
rect 27249 39791 27307 39797
rect 27522 39788 27528 39800
rect 27580 39788 27586 39840
rect 27706 39788 27712 39840
rect 27764 39788 27770 39840
rect 29086 39788 29092 39840
rect 29144 39828 29150 39840
rect 29825 39831 29883 39837
rect 29825 39828 29837 39831
rect 29144 39800 29837 39828
rect 29144 39788 29150 39800
rect 29825 39797 29837 39800
rect 29871 39797 29883 39831
rect 29825 39791 29883 39797
rect 30834 39788 30840 39840
rect 30892 39828 30898 39840
rect 31113 39831 31171 39837
rect 31113 39828 31125 39831
rect 30892 39800 31125 39828
rect 30892 39788 30898 39800
rect 31113 39797 31125 39800
rect 31159 39797 31171 39831
rect 31113 39791 31171 39797
rect 31570 39788 31576 39840
rect 31628 39788 31634 39840
rect 34606 39788 34612 39840
rect 34664 39828 34670 39840
rect 34701 39831 34759 39837
rect 34701 39828 34713 39831
rect 34664 39800 34713 39828
rect 34664 39788 34670 39800
rect 34701 39797 34713 39800
rect 34747 39797 34759 39831
rect 35084 39828 35112 39868
rect 36740 39868 38976 39896
rect 39040 39868 39681 39896
rect 36740 39828 36768 39868
rect 35084 39800 36768 39828
rect 34701 39791 34759 39797
rect 37550 39788 37556 39840
rect 37608 39828 37614 39840
rect 38013 39831 38071 39837
rect 38013 39828 38025 39831
rect 37608 39800 38025 39828
rect 37608 39788 37614 39800
rect 38013 39797 38025 39800
rect 38059 39797 38071 39831
rect 38013 39791 38071 39797
rect 38102 39788 38108 39840
rect 38160 39828 38166 39840
rect 38657 39831 38715 39837
rect 38657 39828 38669 39831
rect 38160 39800 38669 39828
rect 38160 39788 38166 39800
rect 38657 39797 38669 39800
rect 38703 39828 38715 39831
rect 39040 39828 39068 39868
rect 39669 39865 39681 39868
rect 39715 39865 39727 39899
rect 39669 39859 39727 39865
rect 40313 39899 40371 39905
rect 40313 39865 40325 39899
rect 40359 39896 40371 39899
rect 42702 39896 42708 39908
rect 40359 39868 42708 39896
rect 40359 39865 40371 39868
rect 40313 39859 40371 39865
rect 42702 39856 42708 39868
rect 42760 39856 42766 39908
rect 38703 39800 39068 39828
rect 39209 39831 39267 39837
rect 38703 39797 38715 39800
rect 38657 39791 38715 39797
rect 39209 39797 39221 39831
rect 39255 39828 39267 39831
rect 39298 39828 39304 39840
rect 39255 39800 39304 39828
rect 39255 39797 39267 39800
rect 39209 39791 39267 39797
rect 39298 39788 39304 39800
rect 39356 39788 39362 39840
rect 39390 39788 39396 39840
rect 39448 39828 39454 39840
rect 42610 39828 42616 39840
rect 39448 39800 42616 39828
rect 39448 39788 39454 39800
rect 42610 39788 42616 39800
rect 42668 39788 42674 39840
rect 43349 39831 43407 39837
rect 43349 39797 43361 39831
rect 43395 39828 43407 39831
rect 43438 39828 43444 39840
rect 43395 39800 43444 39828
rect 43395 39797 43407 39800
rect 43349 39791 43407 39797
rect 43438 39788 43444 39800
rect 43496 39788 43502 39840
rect 1104 39738 43884 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 43884 39738
rect 1104 39664 43884 39686
rect 16114 39584 16120 39636
rect 16172 39624 16178 39636
rect 17773 39627 17831 39633
rect 17773 39624 17785 39627
rect 16172 39596 17785 39624
rect 16172 39584 16178 39596
rect 17773 39593 17785 39596
rect 17819 39624 17831 39627
rect 18322 39624 18328 39636
rect 17819 39596 18328 39624
rect 17819 39593 17831 39596
rect 17773 39587 17831 39593
rect 18322 39584 18328 39596
rect 18380 39584 18386 39636
rect 18874 39584 18880 39636
rect 18932 39584 18938 39636
rect 20073 39627 20131 39633
rect 20073 39593 20085 39627
rect 20119 39624 20131 39627
rect 20622 39624 20628 39636
rect 20119 39596 20628 39624
rect 20119 39593 20131 39596
rect 20073 39587 20131 39593
rect 20622 39584 20628 39596
rect 20680 39584 20686 39636
rect 23106 39584 23112 39636
rect 23164 39584 23170 39636
rect 23569 39627 23627 39633
rect 23569 39593 23581 39627
rect 23615 39593 23627 39627
rect 23569 39587 23627 39593
rect 28629 39627 28687 39633
rect 28629 39593 28641 39627
rect 28675 39624 28687 39627
rect 28718 39624 28724 39636
rect 28675 39596 28724 39624
rect 28675 39593 28687 39596
rect 28629 39587 28687 39593
rect 20257 39559 20315 39565
rect 20257 39525 20269 39559
rect 20303 39556 20315 39559
rect 20806 39556 20812 39568
rect 20303 39528 20812 39556
rect 20303 39525 20315 39528
rect 20257 39519 20315 39525
rect 20806 39516 20812 39528
rect 20864 39516 20870 39568
rect 22186 39516 22192 39568
rect 22244 39556 22250 39568
rect 23584 39556 23612 39587
rect 28718 39584 28724 39596
rect 28776 39584 28782 39636
rect 36078 39633 36084 39636
rect 36072 39587 36084 39633
rect 36136 39624 36142 39636
rect 41322 39624 41328 39636
rect 36136 39596 36172 39624
rect 38212 39596 41328 39624
rect 36078 39584 36084 39587
rect 36136 39584 36142 39596
rect 29730 39556 29736 39568
rect 22244 39528 29736 39556
rect 22244 39516 22250 39528
rect 29730 39516 29736 39528
rect 29788 39516 29794 39568
rect 32217 39559 32275 39565
rect 32217 39525 32229 39559
rect 32263 39556 32275 39559
rect 33686 39556 33692 39568
rect 32263 39528 33692 39556
rect 32263 39525 32275 39528
rect 32217 39519 32275 39525
rect 33686 39516 33692 39528
rect 33744 39516 33750 39568
rect 35434 39516 35440 39568
rect 35492 39516 35498 39568
rect 36725 39559 36783 39565
rect 36725 39525 36737 39559
rect 36771 39556 36783 39559
rect 36906 39556 36912 39568
rect 36771 39528 36912 39556
rect 36771 39525 36783 39528
rect 36725 39519 36783 39525
rect 36906 39516 36912 39528
rect 36964 39516 36970 39568
rect 37182 39516 37188 39568
rect 37240 39556 37246 39568
rect 38212 39556 38240 39596
rect 41322 39584 41328 39596
rect 41380 39584 41386 39636
rect 43257 39627 43315 39633
rect 43257 39624 43269 39627
rect 41800 39596 43269 39624
rect 40034 39556 40040 39568
rect 37240 39528 38240 39556
rect 39408 39528 40040 39556
rect 37240 39516 37246 39528
rect 24946 39488 24952 39500
rect 23308 39460 24952 39488
rect 18782 39380 18788 39432
rect 18840 39380 18846 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 19613 39423 19671 39429
rect 19613 39420 19625 39423
rect 19484 39392 19625 39420
rect 19484 39380 19490 39392
rect 19613 39389 19625 39392
rect 19659 39389 19671 39423
rect 19613 39383 19671 39389
rect 20714 39380 20720 39432
rect 20772 39420 20778 39432
rect 20993 39423 21051 39429
rect 20993 39420 21005 39423
rect 20772 39392 21005 39420
rect 20772 39380 20778 39392
rect 20993 39389 21005 39392
rect 21039 39389 21051 39423
rect 20993 39383 21051 39389
rect 21082 39380 21088 39432
rect 21140 39420 21146 39432
rect 21249 39423 21307 39429
rect 21249 39420 21261 39423
rect 21140 39392 21261 39420
rect 21140 39380 21146 39392
rect 21249 39389 21261 39392
rect 21295 39389 21307 39423
rect 21249 39383 21307 39389
rect 22922 39380 22928 39432
rect 22980 39420 22986 39432
rect 23308 39429 23336 39460
rect 24946 39448 24952 39460
rect 25004 39448 25010 39500
rect 26510 39448 26516 39500
rect 26568 39448 26574 39500
rect 26786 39448 26792 39500
rect 26844 39448 26850 39500
rect 28350 39448 28356 39500
rect 28408 39448 28414 39500
rect 29825 39491 29883 39497
rect 29825 39457 29837 39491
rect 29871 39488 29883 39491
rect 30282 39488 30288 39500
rect 29871 39460 30288 39488
rect 29871 39457 29883 39460
rect 29825 39451 29883 39457
rect 30282 39448 30288 39460
rect 30340 39448 30346 39500
rect 31754 39448 31760 39500
rect 31812 39488 31818 39500
rect 35161 39491 35219 39497
rect 31812 39460 35112 39488
rect 31812 39448 31818 39460
rect 23293 39423 23351 39429
rect 23293 39420 23305 39423
rect 22980 39392 23305 39420
rect 22980 39380 22986 39392
rect 23293 39389 23305 39392
rect 23339 39389 23351 39423
rect 23293 39383 23351 39389
rect 23658 39380 23664 39432
rect 23716 39380 23722 39432
rect 24578 39380 24584 39432
rect 24636 39420 24642 39432
rect 24857 39423 24915 39429
rect 24857 39420 24869 39423
rect 24636 39392 24869 39420
rect 24636 39380 24642 39392
rect 24857 39389 24869 39392
rect 24903 39389 24915 39423
rect 24857 39383 24915 39389
rect 25038 39380 25044 39432
rect 25096 39380 25102 39432
rect 25225 39423 25283 39429
rect 25225 39389 25237 39423
rect 25271 39420 25283 39423
rect 26421 39423 26479 39429
rect 26421 39420 26433 39423
rect 25271 39392 26433 39420
rect 25271 39389 25283 39392
rect 25225 39383 25283 39389
rect 26421 39389 26433 39392
rect 26467 39420 26479 39423
rect 27433 39423 27491 39429
rect 27433 39420 27445 39423
rect 26467 39392 27445 39420
rect 26467 39389 26479 39392
rect 26421 39383 26479 39389
rect 27433 39389 27445 39392
rect 27479 39389 27491 39423
rect 27433 39383 27491 39389
rect 27617 39423 27675 39429
rect 27617 39389 27629 39423
rect 27663 39420 27675 39423
rect 28261 39423 28319 39429
rect 28261 39420 28273 39423
rect 27663 39392 28273 39420
rect 27663 39389 27675 39392
rect 27617 39383 27675 39389
rect 28261 39389 28273 39392
rect 28307 39420 28319 39423
rect 28902 39420 28908 39432
rect 28307 39392 28908 39420
rect 28307 39389 28319 39392
rect 28261 39383 28319 39389
rect 28902 39380 28908 39392
rect 28960 39380 28966 39432
rect 31409 39423 31467 39429
rect 31409 39389 31421 39423
rect 31455 39420 31467 39423
rect 31570 39420 31576 39432
rect 31455 39392 31576 39420
rect 31455 39389 31467 39392
rect 31409 39383 31467 39389
rect 31570 39380 31576 39392
rect 31628 39380 31634 39432
rect 31662 39380 31668 39432
rect 31720 39380 31726 39432
rect 32858 39380 32864 39432
rect 32916 39380 32922 39432
rect 33229 39423 33287 39429
rect 33229 39389 33241 39423
rect 33275 39420 33287 39423
rect 34514 39420 34520 39432
rect 33275 39392 34520 39420
rect 33275 39389 33287 39392
rect 33229 39383 33287 39389
rect 34514 39380 34520 39392
rect 34572 39380 34578 39432
rect 35084 39429 35112 39460
rect 35161 39457 35173 39491
rect 35207 39488 35219 39491
rect 35342 39488 35348 39500
rect 35207 39460 35348 39488
rect 35207 39457 35219 39460
rect 35161 39451 35219 39457
rect 35342 39448 35348 39460
rect 35400 39488 35406 39500
rect 36078 39488 36084 39500
rect 35400 39460 36084 39488
rect 35400 39448 35406 39460
rect 36078 39448 36084 39460
rect 36136 39488 36142 39500
rect 39209 39491 39267 39497
rect 36136 39460 37044 39488
rect 36136 39448 36142 39460
rect 37016 39429 37044 39460
rect 39209 39457 39221 39491
rect 39255 39488 39267 39491
rect 39408 39488 39436 39528
rect 40034 39516 40040 39528
rect 40092 39516 40098 39568
rect 39255 39460 39436 39488
rect 39485 39491 39543 39497
rect 39255 39457 39267 39460
rect 39209 39451 39267 39457
rect 39485 39457 39497 39491
rect 39531 39488 39543 39491
rect 39531 39460 40172 39488
rect 39531 39457 39543 39460
rect 39485 39451 39543 39457
rect 35069 39423 35127 39429
rect 35069 39389 35081 39423
rect 35115 39389 35127 39423
rect 36909 39423 36967 39429
rect 36909 39420 36921 39423
rect 35069 39383 35127 39389
rect 35912 39392 36921 39420
rect 18800 39352 18828 39380
rect 18800 39324 19564 39352
rect 18874 39244 18880 39296
rect 18932 39284 18938 39296
rect 19429 39287 19487 39293
rect 19429 39284 19441 39287
rect 18932 39256 19441 39284
rect 18932 39244 18938 39256
rect 19429 39253 19441 39256
rect 19475 39253 19487 39287
rect 19536 39284 19564 39324
rect 20530 39312 20536 39364
rect 20588 39352 20594 39364
rect 22186 39352 22192 39364
rect 20588 39324 22192 39352
rect 20588 39312 20594 39324
rect 22186 39312 22192 39324
rect 22244 39312 22250 39364
rect 22296 39324 26464 39352
rect 22296 39284 22324 39324
rect 19536 39256 22324 39284
rect 22373 39287 22431 39293
rect 19429 39247 19487 39253
rect 22373 39253 22385 39287
rect 22419 39284 22431 39287
rect 22922 39284 22928 39296
rect 22419 39256 22928 39284
rect 22419 39253 22431 39256
rect 22373 39247 22431 39253
rect 22922 39244 22928 39256
rect 22980 39244 22986 39296
rect 25038 39244 25044 39296
rect 25096 39284 25102 39296
rect 25685 39287 25743 39293
rect 25685 39284 25697 39287
rect 25096 39256 25697 39284
rect 25096 39244 25102 39256
rect 25685 39253 25697 39256
rect 25731 39253 25743 39287
rect 26436 39284 26464 39324
rect 26510 39312 26516 39364
rect 26568 39352 26574 39364
rect 27249 39355 27307 39361
rect 27249 39352 27261 39355
rect 26568 39324 27261 39352
rect 26568 39312 26574 39324
rect 27249 39321 27261 39324
rect 27295 39321 27307 39355
rect 29638 39352 29644 39364
rect 27249 39315 27307 39321
rect 28920 39324 29644 39352
rect 28920 39284 28948 39324
rect 29638 39312 29644 39324
rect 29696 39312 29702 39364
rect 32582 39312 32588 39364
rect 32640 39352 32646 39364
rect 33045 39355 33103 39361
rect 33045 39352 33057 39355
rect 32640 39324 33057 39352
rect 32640 39312 32646 39324
rect 33045 39321 33057 39324
rect 33091 39321 33103 39355
rect 33045 39315 33103 39321
rect 33137 39355 33195 39361
rect 33137 39321 33149 39355
rect 33183 39321 33195 39355
rect 35084 39352 35112 39383
rect 35912 39361 35940 39392
rect 36909 39389 36921 39392
rect 36955 39389 36967 39423
rect 36909 39383 36967 39389
rect 37001 39423 37059 39429
rect 37001 39389 37013 39423
rect 37047 39389 37059 39423
rect 37001 39383 37059 39389
rect 38010 39380 38016 39432
rect 38068 39380 38074 39432
rect 39114 39420 39120 39432
rect 38488 39392 39120 39420
rect 35897 39355 35955 39361
rect 35897 39352 35909 39355
rect 35084 39324 35909 39352
rect 33137 39315 33195 39321
rect 35897 39321 35909 39324
rect 35943 39321 35955 39355
rect 36725 39355 36783 39361
rect 36725 39352 36737 39355
rect 35897 39315 35955 39321
rect 36188 39324 36737 39352
rect 26436 39256 28948 39284
rect 25685 39247 25743 39253
rect 28994 39244 29000 39296
rect 29052 39284 29058 39296
rect 29089 39287 29147 39293
rect 29089 39284 29101 39287
rect 29052 39256 29101 39284
rect 29052 39244 29058 39256
rect 29089 39253 29101 39256
rect 29135 39253 29147 39287
rect 29089 39247 29147 39253
rect 29454 39244 29460 39296
rect 29512 39284 29518 39296
rect 30190 39284 30196 39296
rect 29512 39256 30196 39284
rect 29512 39244 29518 39256
rect 30190 39244 30196 39256
rect 30248 39284 30254 39296
rect 30285 39287 30343 39293
rect 30285 39284 30297 39287
rect 30248 39256 30297 39284
rect 30248 39244 30254 39256
rect 30285 39253 30297 39256
rect 30331 39253 30343 39287
rect 33152 39284 33180 39315
rect 33226 39284 33232 39296
rect 33152 39256 33232 39284
rect 30285 39247 30343 39253
rect 33226 39244 33232 39256
rect 33284 39244 33290 39296
rect 33318 39244 33324 39296
rect 33376 39284 33382 39296
rect 33413 39287 33471 39293
rect 33413 39284 33425 39287
rect 33376 39256 33425 39284
rect 33376 39244 33382 39256
rect 33413 39253 33425 39256
rect 33459 39253 33471 39287
rect 33413 39247 33471 39253
rect 33594 39244 33600 39296
rect 33652 39284 33658 39296
rect 33870 39284 33876 39296
rect 33652 39256 33876 39284
rect 33652 39244 33658 39256
rect 33870 39244 33876 39256
rect 33928 39284 33934 39296
rect 33965 39287 34023 39293
rect 33965 39284 33977 39287
rect 33928 39256 33977 39284
rect 33928 39244 33934 39256
rect 33965 39253 33977 39256
rect 34011 39284 34023 39287
rect 35986 39284 35992 39296
rect 34011 39256 35992 39284
rect 34011 39253 34023 39256
rect 33965 39247 34023 39253
rect 35986 39244 35992 39256
rect 36044 39244 36050 39296
rect 36078 39244 36084 39296
rect 36136 39293 36142 39296
rect 36136 39287 36155 39293
rect 36143 39284 36155 39287
rect 36188 39284 36216 39324
rect 36725 39321 36737 39324
rect 36771 39321 36783 39355
rect 38488 39352 38516 39392
rect 39114 39380 39120 39392
rect 39172 39380 39178 39432
rect 40037 39423 40095 39429
rect 40037 39389 40049 39423
rect 40083 39389 40095 39423
rect 40144 39420 40172 39460
rect 40293 39423 40351 39429
rect 40293 39420 40305 39423
rect 40144 39392 40305 39420
rect 40037 39383 40095 39389
rect 40293 39389 40305 39392
rect 40339 39389 40351 39423
rect 41800 39420 41828 39596
rect 43257 39593 43269 39596
rect 43303 39593 43315 39627
rect 43257 39587 43315 39593
rect 40293 39383 40351 39389
rect 40420 39392 41828 39420
rect 36725 39315 36783 39321
rect 36832 39324 38516 39352
rect 36143 39256 36216 39284
rect 36143 39253 36155 39256
rect 36136 39247 36155 39253
rect 36136 39244 36142 39247
rect 36262 39244 36268 39296
rect 36320 39284 36326 39296
rect 36832 39284 36860 39324
rect 38838 39312 38844 39364
rect 38896 39352 38902 39364
rect 40052 39352 40080 39383
rect 40420 39364 40448 39392
rect 41874 39380 41880 39432
rect 41932 39380 41938 39432
rect 38896 39324 40080 39352
rect 38896 39312 38902 39324
rect 40402 39312 40408 39364
rect 40460 39312 40466 39364
rect 41138 39312 41144 39364
rect 41196 39352 41202 39364
rect 42122 39355 42180 39361
rect 42122 39352 42134 39355
rect 41196 39324 42134 39352
rect 41196 39312 41202 39324
rect 42122 39321 42134 39324
rect 42168 39321 42180 39355
rect 42122 39315 42180 39321
rect 36320 39256 36860 39284
rect 37553 39287 37611 39293
rect 36320 39244 36326 39256
rect 37553 39253 37565 39287
rect 37599 39284 37611 39287
rect 38562 39284 38568 39296
rect 37599 39256 38568 39284
rect 37599 39253 37611 39256
rect 37553 39247 37611 39253
rect 38562 39244 38568 39256
rect 38620 39284 38626 39296
rect 39298 39284 39304 39296
rect 38620 39256 39304 39284
rect 38620 39244 38626 39256
rect 39298 39244 39304 39256
rect 39356 39244 39362 39296
rect 40310 39244 40316 39296
rect 40368 39284 40374 39296
rect 41417 39287 41475 39293
rect 41417 39284 41429 39287
rect 40368 39256 41429 39284
rect 40368 39244 40374 39256
rect 41417 39253 41429 39256
rect 41463 39253 41475 39287
rect 41417 39247 41475 39253
rect 1104 39194 43884 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 43884 39194
rect 1104 39120 43884 39142
rect 19978 39040 19984 39092
rect 20036 39080 20042 39092
rect 20349 39083 20407 39089
rect 20349 39080 20361 39083
rect 20036 39052 20361 39080
rect 20036 39040 20042 39052
rect 20349 39049 20361 39052
rect 20395 39049 20407 39083
rect 23658 39080 23664 39092
rect 20349 39043 20407 39049
rect 20824 39052 23664 39080
rect 20824 39024 20852 39052
rect 23658 39040 23664 39052
rect 23716 39040 23722 39092
rect 24213 39083 24271 39089
rect 24213 39080 24225 39083
rect 24044 39052 24225 39080
rect 18776 39015 18834 39021
rect 18776 38981 18788 39015
rect 18822 39012 18834 39015
rect 18874 39012 18880 39024
rect 18822 38984 18880 39012
rect 18822 38981 18834 38984
rect 18776 38975 18834 38981
rect 18874 38972 18880 38984
rect 18932 38972 18938 39024
rect 20806 38972 20812 39024
rect 20864 38972 20870 39024
rect 22373 39015 22431 39021
rect 22373 38981 22385 39015
rect 22419 39012 22431 39015
rect 22462 39012 22468 39024
rect 22419 38984 22468 39012
rect 22419 38981 22431 38984
rect 22373 38975 22431 38981
rect 22462 38972 22468 38984
rect 22520 38972 22526 39024
rect 22738 38972 22744 39024
rect 22796 39012 22802 39024
rect 24044 39012 24072 39052
rect 24213 39049 24225 39052
rect 24259 39080 24271 39083
rect 24486 39080 24492 39092
rect 24259 39052 24492 39080
rect 24259 39049 24271 39052
rect 24213 39043 24271 39049
rect 24486 39040 24492 39052
rect 24544 39040 24550 39092
rect 24578 39040 24584 39092
rect 24636 39080 24642 39092
rect 25034 39083 25092 39089
rect 25034 39080 25046 39083
rect 24636 39052 25046 39080
rect 24636 39040 24642 39052
rect 25034 39049 25046 39052
rect 25080 39049 25092 39083
rect 25034 39043 25092 39049
rect 29638 39040 29644 39092
rect 29696 39080 29702 39092
rect 29733 39083 29791 39089
rect 29733 39080 29745 39083
rect 29696 39052 29745 39080
rect 29696 39040 29702 39052
rect 29733 39049 29745 39052
rect 29779 39049 29791 39083
rect 29733 39043 29791 39049
rect 31018 39040 31024 39092
rect 31076 39040 31082 39092
rect 31573 39083 31631 39089
rect 31573 39049 31585 39083
rect 31619 39080 31631 39083
rect 31754 39080 31760 39092
rect 31619 39052 31760 39080
rect 31619 39049 31631 39052
rect 31573 39043 31631 39049
rect 31754 39040 31760 39052
rect 31812 39040 31818 39092
rect 32582 39040 32588 39092
rect 32640 39080 32646 39092
rect 37642 39080 37648 39092
rect 32640 39052 37648 39080
rect 32640 39040 32646 39052
rect 22796 38984 24072 39012
rect 24136 38984 25084 39012
rect 22796 38972 22802 38984
rect 16574 38904 16580 38956
rect 16632 38944 16638 38956
rect 17497 38947 17555 38953
rect 17497 38944 17509 38947
rect 16632 38916 17509 38944
rect 16632 38904 16638 38916
rect 17497 38913 17509 38916
rect 17543 38944 17555 38947
rect 21174 38944 21180 38956
rect 17543 38916 21180 38944
rect 17543 38913 17555 38916
rect 17497 38907 17555 38913
rect 21174 38904 21180 38916
rect 21232 38904 21238 38956
rect 22094 38904 22100 38956
rect 22152 38953 22158 38956
rect 22152 38947 22201 38953
rect 22152 38913 22155 38947
rect 22189 38913 22201 38947
rect 22152 38907 22201 38913
rect 22281 38947 22339 38953
rect 22281 38913 22293 38947
rect 22327 38913 22339 38947
rect 22554 38944 22560 38956
rect 22515 38916 22560 38944
rect 22281 38907 22339 38913
rect 22152 38904 22158 38907
rect 18046 38836 18052 38888
rect 18104 38876 18110 38888
rect 18509 38879 18567 38885
rect 18509 38876 18521 38879
rect 18104 38848 18521 38876
rect 18104 38836 18110 38848
rect 18509 38845 18521 38848
rect 18555 38845 18567 38879
rect 22296 38876 22324 38907
rect 22554 38904 22560 38916
rect 22612 38904 22618 38956
rect 22646 38904 22652 38956
rect 22704 38904 22710 38956
rect 24136 38953 24164 38984
rect 24121 38947 24179 38953
rect 24121 38913 24133 38947
rect 24167 38913 24179 38947
rect 24121 38907 24179 38913
rect 24394 38904 24400 38956
rect 24452 38904 24458 38956
rect 24872 38953 24900 38984
rect 24857 38947 24915 38953
rect 24857 38913 24869 38947
rect 24903 38913 24915 38947
rect 24857 38907 24915 38913
rect 24949 38947 25007 38953
rect 24949 38913 24961 38947
rect 24995 38913 25007 38947
rect 24949 38907 25007 38913
rect 18509 38839 18567 38845
rect 19904 38848 24900 38876
rect 16942 38768 16948 38820
rect 17000 38768 17006 38820
rect 19794 38768 19800 38820
rect 19852 38808 19858 38820
rect 19904 38817 19932 38848
rect 24872 38820 24900 38848
rect 19889 38811 19947 38817
rect 19889 38808 19901 38811
rect 19852 38780 19901 38808
rect 19852 38768 19858 38780
rect 19889 38777 19901 38780
rect 19935 38777 19947 38811
rect 19889 38771 19947 38777
rect 20530 38768 20536 38820
rect 20588 38768 20594 38820
rect 20990 38768 20996 38820
rect 21048 38808 21054 38820
rect 22005 38811 22063 38817
rect 22005 38808 22017 38811
rect 21048 38780 22017 38808
rect 21048 38768 21054 38780
rect 22005 38777 22017 38780
rect 22051 38777 22063 38811
rect 22005 38771 22063 38777
rect 24210 38768 24216 38820
rect 24268 38808 24274 38820
rect 24397 38811 24455 38817
rect 24397 38808 24409 38811
rect 24268 38780 24409 38808
rect 24268 38768 24274 38780
rect 24397 38777 24409 38780
rect 24443 38777 24455 38811
rect 24397 38771 24455 38777
rect 24854 38768 24860 38820
rect 24912 38768 24918 38820
rect 24964 38808 24992 38907
rect 25056 38876 25084 38984
rect 26786 38972 26792 39024
rect 26844 39012 26850 39024
rect 27402 39015 27460 39021
rect 27402 39012 27414 39015
rect 26844 38984 27414 39012
rect 26844 38972 26850 38984
rect 27402 38981 27414 38984
rect 27448 38981 27460 39015
rect 27402 38975 27460 38981
rect 27522 38972 27528 39024
rect 27580 39012 27586 39024
rect 29822 39012 29828 39024
rect 27580 38984 29828 39012
rect 27580 38972 27586 38984
rect 29822 38972 29828 38984
rect 29880 39012 29886 39024
rect 30558 39012 30564 39024
rect 29880 38984 30564 39012
rect 29880 38972 29886 38984
rect 30558 38972 30564 38984
rect 30616 38972 30622 39024
rect 30668 38984 31524 39012
rect 30668 38956 30696 38984
rect 25130 38904 25136 38956
rect 25188 38904 25194 38956
rect 28626 38904 28632 38956
rect 28684 38944 28690 38956
rect 28997 38947 29055 38953
rect 28997 38944 29009 38947
rect 28684 38916 29009 38944
rect 28684 38904 28690 38916
rect 28997 38913 29009 38916
rect 29043 38913 29055 38947
rect 28997 38907 29055 38913
rect 29086 38904 29092 38956
rect 29144 38944 29150 38956
rect 29181 38947 29239 38953
rect 29181 38944 29193 38947
rect 29144 38916 29193 38944
rect 29144 38904 29150 38916
rect 29181 38913 29193 38916
rect 29227 38913 29239 38947
rect 29181 38907 29239 38913
rect 29273 38947 29331 38953
rect 29273 38913 29285 38947
rect 29319 38913 29331 38947
rect 29273 38907 29331 38913
rect 26786 38876 26792 38888
rect 25056 38848 26792 38876
rect 26786 38836 26792 38848
rect 26844 38836 26850 38888
rect 27154 38836 27160 38888
rect 27212 38836 27218 38888
rect 29288 38820 29316 38907
rect 30650 38904 30656 38956
rect 30708 38904 30714 38956
rect 30834 38904 30840 38956
rect 30892 38904 30898 38956
rect 31496 38953 31524 38984
rect 32674 38972 32680 39024
rect 32732 39012 32738 39024
rect 32861 39015 32919 39021
rect 32861 39012 32873 39015
rect 32732 38984 32873 39012
rect 32732 38972 32738 38984
rect 32861 38981 32873 38984
rect 32907 38981 32919 39015
rect 32861 38975 32919 38981
rect 33612 38984 33824 39012
rect 33612 38956 33640 38984
rect 31481 38947 31539 38953
rect 31481 38913 31493 38947
rect 31527 38913 31539 38947
rect 31481 38907 31539 38913
rect 31665 38947 31723 38953
rect 31665 38913 31677 38947
rect 31711 38913 31723 38947
rect 33321 38947 33379 38953
rect 33321 38944 33333 38947
rect 31665 38907 31723 38913
rect 33244 38916 33333 38944
rect 30852 38876 30880 38904
rect 31680 38876 31708 38907
rect 33244 38888 33272 38916
rect 33321 38913 33333 38916
rect 33367 38913 33379 38947
rect 33321 38907 33379 38913
rect 33594 38904 33600 38956
rect 33652 38904 33658 38956
rect 33689 38947 33747 38953
rect 33689 38913 33701 38947
rect 33735 38913 33747 38947
rect 33689 38907 33747 38913
rect 30852 38848 31708 38876
rect 33226 38836 33232 38888
rect 33284 38836 33290 38888
rect 25314 38808 25320 38820
rect 24964 38780 25320 38808
rect 25314 38768 25320 38780
rect 25372 38808 25378 38820
rect 26326 38808 26332 38820
rect 25372 38780 26332 38808
rect 25372 38768 25378 38780
rect 26326 38768 26332 38780
rect 26384 38768 26390 38820
rect 28350 38768 28356 38820
rect 28408 38808 28414 38820
rect 28997 38811 29055 38817
rect 28997 38808 29009 38811
rect 28408 38780 29009 38808
rect 28408 38768 28414 38780
rect 28997 38777 29009 38780
rect 29043 38777 29055 38811
rect 28997 38771 29055 38777
rect 29270 38768 29276 38820
rect 29328 38808 29334 38820
rect 31386 38808 31392 38820
rect 29328 38780 31392 38808
rect 29328 38768 29334 38780
rect 31386 38768 31392 38780
rect 31444 38768 31450 38820
rect 31754 38768 31760 38820
rect 31812 38808 31818 38820
rect 31812 38780 32444 38808
rect 31812 38768 31818 38780
rect 18049 38743 18107 38749
rect 18049 38709 18061 38743
rect 18095 38740 18107 38743
rect 20254 38740 20260 38752
rect 18095 38712 20260 38740
rect 18095 38709 18107 38712
rect 18049 38703 18107 38709
rect 20254 38700 20260 38712
rect 20312 38700 20318 38752
rect 21358 38700 21364 38752
rect 21416 38700 21422 38752
rect 23201 38743 23259 38749
rect 23201 38709 23213 38743
rect 23247 38740 23259 38743
rect 23382 38740 23388 38752
rect 23247 38712 23388 38740
rect 23247 38709 23259 38712
rect 23201 38703 23259 38709
rect 23382 38700 23388 38712
rect 23440 38700 23446 38752
rect 25590 38700 25596 38752
rect 25648 38700 25654 38752
rect 26418 38700 26424 38752
rect 26476 38700 26482 38752
rect 28442 38700 28448 38752
rect 28500 38740 28506 38752
rect 28537 38743 28595 38749
rect 28537 38740 28549 38743
rect 28500 38712 28549 38740
rect 28500 38700 28506 38712
rect 28537 38709 28549 38712
rect 28583 38709 28595 38743
rect 28537 38703 28595 38709
rect 28902 38700 28908 38752
rect 28960 38740 28966 38752
rect 32309 38743 32367 38749
rect 32309 38740 32321 38743
rect 28960 38712 32321 38740
rect 28960 38700 28966 38712
rect 32309 38709 32321 38712
rect 32355 38709 32367 38743
rect 32416 38740 32444 38780
rect 32858 38768 32864 38820
rect 32916 38808 32922 38820
rect 33134 38808 33140 38820
rect 32916 38780 33140 38808
rect 32916 38768 32922 38780
rect 33134 38768 33140 38780
rect 33192 38768 33198 38820
rect 33704 38740 33732 38907
rect 33796 38808 33824 38984
rect 33980 38953 34008 39052
rect 34790 38972 34796 39024
rect 34848 38972 34854 39024
rect 33965 38947 34023 38953
rect 33965 38913 33977 38947
rect 34011 38913 34023 38947
rect 33965 38907 34023 38913
rect 34238 38904 34244 38956
rect 34296 38904 34302 38956
rect 34422 38904 34428 38956
rect 34480 38944 34486 38956
rect 35253 38947 35311 38953
rect 35253 38944 35265 38947
rect 34480 38916 35265 38944
rect 34480 38904 34486 38916
rect 35253 38913 35265 38916
rect 35299 38913 35311 38947
rect 35253 38907 35311 38913
rect 35526 38904 35532 38956
rect 35584 38904 35590 38956
rect 35618 38904 35624 38956
rect 35676 38904 35682 38956
rect 35912 38953 35940 39052
rect 37642 39040 37648 39052
rect 37700 39040 37706 39092
rect 39298 39040 39304 39092
rect 39356 39040 39362 39092
rect 41138 39040 41144 39092
rect 41196 39040 41202 39092
rect 41785 39083 41843 39089
rect 41785 39049 41797 39083
rect 41831 39080 41843 39083
rect 42610 39080 42616 39092
rect 41831 39052 42616 39080
rect 41831 39049 41843 39052
rect 41785 39043 41843 39049
rect 42610 39040 42616 39052
rect 42668 39080 42674 39092
rect 43165 39083 43223 39089
rect 43165 39080 43177 39083
rect 42668 39052 43177 39080
rect 42668 39040 42674 39052
rect 43165 39049 43177 39052
rect 43211 39049 43223 39083
rect 43165 39043 43223 39049
rect 35986 38972 35992 39024
rect 36044 39012 36050 39024
rect 36817 39015 36875 39021
rect 36044 38984 36216 39012
rect 36044 38972 36050 38984
rect 35897 38947 35955 38953
rect 35897 38913 35909 38947
rect 35943 38913 35955 38947
rect 35897 38907 35955 38913
rect 36081 38947 36139 38953
rect 36081 38913 36093 38947
rect 36127 38913 36139 38947
rect 36081 38907 36139 38913
rect 34698 38836 34704 38888
rect 34756 38876 34762 38888
rect 35434 38876 35440 38888
rect 34756 38848 35440 38876
rect 34756 38836 34762 38848
rect 35434 38836 35440 38848
rect 35492 38876 35498 38888
rect 36096 38876 36124 38907
rect 35492 38848 36124 38876
rect 36188 38876 36216 38984
rect 36817 38981 36829 39015
rect 36863 39012 36875 39015
rect 38574 39015 38632 39021
rect 38574 39012 38586 39015
rect 36863 38984 38586 39012
rect 36863 38981 36875 38984
rect 36817 38975 36875 38981
rect 38574 38981 38586 38984
rect 38620 38981 38632 39015
rect 38574 38975 38632 38981
rect 39114 38972 39120 39024
rect 39172 39012 39178 39024
rect 40037 39015 40095 39021
rect 40037 39012 40049 39015
rect 39172 38984 40049 39012
rect 39172 38972 39178 38984
rect 40037 38981 40049 38984
rect 40083 39012 40095 39015
rect 40126 39012 40132 39024
rect 40083 38984 40132 39012
rect 40083 38981 40095 38984
rect 40037 38975 40095 38981
rect 40126 38972 40132 38984
rect 40184 38972 40190 39024
rect 40253 39015 40311 39021
rect 40253 38981 40265 39015
rect 40299 39012 40311 39015
rect 40678 39012 40684 39024
rect 40299 38984 40684 39012
rect 40299 38981 40311 38984
rect 40253 38975 40311 38981
rect 40678 38972 40684 38984
rect 40736 38972 40742 39024
rect 36262 38904 36268 38956
rect 36320 38944 36326 38956
rect 36725 38947 36783 38953
rect 36725 38944 36737 38947
rect 36320 38916 36737 38944
rect 36320 38904 36326 38916
rect 36725 38913 36737 38916
rect 36771 38913 36783 38947
rect 36725 38907 36783 38913
rect 36906 38904 36912 38956
rect 36964 38904 36970 38956
rect 40862 38944 40868 38956
rect 37016 38916 40868 38944
rect 37016 38876 37044 38916
rect 40862 38904 40868 38916
rect 40920 38904 40926 38956
rect 41046 38904 41052 38956
rect 41104 38904 41110 38956
rect 41233 38947 41291 38953
rect 41233 38913 41245 38947
rect 41279 38913 41291 38947
rect 41233 38907 41291 38913
rect 36188 38848 37044 38876
rect 35492 38836 35498 38848
rect 38838 38836 38844 38888
rect 38896 38836 38902 38888
rect 41138 38876 41144 38888
rect 40420 38848 41144 38876
rect 40310 38808 40316 38820
rect 33796 38780 37596 38808
rect 32416 38712 33732 38740
rect 32309 38703 32367 38709
rect 33778 38700 33784 38752
rect 33836 38740 33842 38752
rect 34238 38740 34244 38752
rect 33836 38712 34244 38740
rect 33836 38700 33842 38712
rect 34238 38700 34244 38712
rect 34296 38700 34302 38752
rect 37274 38700 37280 38752
rect 37332 38740 37338 38752
rect 37461 38743 37519 38749
rect 37461 38740 37473 38743
rect 37332 38712 37473 38740
rect 37332 38700 37338 38712
rect 37461 38709 37473 38712
rect 37507 38709 37519 38743
rect 37568 38740 37596 38780
rect 39960 38780 40316 38808
rect 39960 38740 39988 38780
rect 40310 38768 40316 38780
rect 40368 38768 40374 38820
rect 40420 38817 40448 38848
rect 41138 38836 41144 38848
rect 41196 38876 41202 38888
rect 41248 38876 41276 38907
rect 41196 38848 41276 38876
rect 41196 38836 41202 38848
rect 40405 38811 40463 38817
rect 40405 38777 40417 38811
rect 40451 38777 40463 38811
rect 40405 38771 40463 38777
rect 40862 38768 40868 38820
rect 40920 38808 40926 38820
rect 42613 38811 42671 38817
rect 42613 38808 42625 38811
rect 40920 38780 42625 38808
rect 40920 38768 40926 38780
rect 42613 38777 42625 38780
rect 42659 38777 42671 38811
rect 42613 38771 42671 38777
rect 37568 38712 39988 38740
rect 37461 38703 37519 38709
rect 40034 38700 40040 38752
rect 40092 38740 40098 38752
rect 40221 38743 40279 38749
rect 40221 38740 40233 38743
rect 40092 38712 40233 38740
rect 40092 38700 40098 38712
rect 40221 38709 40233 38712
rect 40267 38709 40279 38743
rect 40221 38703 40279 38709
rect 1104 38650 43884 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 43884 38650
rect 1104 38576 43884 38598
rect 16485 38539 16543 38545
rect 16485 38505 16497 38539
rect 16531 38536 16543 38539
rect 18782 38536 18788 38548
rect 16531 38508 18788 38536
rect 16531 38505 16543 38508
rect 16485 38499 16543 38505
rect 18782 38496 18788 38508
rect 18840 38496 18846 38548
rect 19426 38496 19432 38548
rect 19484 38496 19490 38548
rect 21361 38539 21419 38545
rect 21361 38505 21373 38539
rect 21407 38536 21419 38539
rect 21450 38536 21456 38548
rect 21407 38508 21456 38536
rect 21407 38505 21419 38508
rect 21361 38499 21419 38505
rect 21450 38496 21456 38508
rect 21508 38496 21514 38548
rect 21634 38496 21640 38548
rect 21692 38536 21698 38548
rect 22094 38536 22100 38548
rect 21692 38508 22100 38536
rect 21692 38496 21698 38508
rect 22094 38496 22100 38508
rect 22152 38496 22158 38548
rect 22462 38496 22468 38548
rect 22520 38536 22526 38548
rect 23106 38536 23112 38548
rect 22520 38508 23112 38536
rect 22520 38496 22526 38508
rect 23106 38496 23112 38508
rect 23164 38496 23170 38548
rect 24394 38496 24400 38548
rect 24452 38536 24458 38548
rect 24581 38539 24639 38545
rect 24581 38536 24593 38539
rect 24452 38508 24593 38536
rect 24452 38496 24458 38508
rect 24581 38505 24593 38508
rect 24627 38505 24639 38539
rect 24581 38499 24639 38505
rect 24670 38496 24676 38548
rect 24728 38536 24734 38548
rect 24728 38508 26740 38536
rect 24728 38496 24734 38508
rect 22480 38468 22508 38496
rect 21008 38440 22508 38468
rect 18966 38360 18972 38412
rect 19024 38400 19030 38412
rect 19426 38400 19432 38412
rect 19024 38372 19432 38400
rect 19024 38360 19030 38372
rect 19426 38360 19432 38372
rect 19484 38400 19490 38412
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 19484 38372 19993 38400
rect 19484 38360 19490 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 19981 38363 20039 38369
rect 20263 38372 20852 38400
rect 17494 38292 17500 38344
rect 17552 38332 17558 38344
rect 18046 38332 18052 38344
rect 17552 38304 18052 38332
rect 17552 38292 17558 38304
rect 18046 38292 18052 38304
rect 18104 38292 18110 38344
rect 19794 38292 19800 38344
rect 19852 38292 19858 38344
rect 19889 38335 19947 38341
rect 19889 38301 19901 38335
rect 19935 38332 19947 38335
rect 20162 38332 20168 38344
rect 19935 38304 20168 38332
rect 19935 38301 19947 38304
rect 19889 38295 19947 38301
rect 20162 38292 20168 38304
rect 20220 38292 20226 38344
rect 17764 38267 17822 38273
rect 17764 38233 17776 38267
rect 17810 38264 17822 38267
rect 18230 38264 18236 38276
rect 17810 38236 18236 38264
rect 17810 38233 17822 38236
rect 17764 38227 17822 38233
rect 18230 38224 18236 38236
rect 18288 38224 18294 38276
rect 20263 38264 20291 38372
rect 20824 38344 20852 38372
rect 20717 38335 20775 38341
rect 20717 38301 20729 38335
rect 20763 38301 20775 38335
rect 20717 38295 20775 38301
rect 18800 38236 20291 38264
rect 14458 38156 14464 38208
rect 14516 38196 14522 38208
rect 17037 38199 17095 38205
rect 17037 38196 17049 38199
rect 14516 38168 17049 38196
rect 14516 38156 14522 38168
rect 17037 38165 17049 38168
rect 17083 38196 17095 38199
rect 18800 38196 18828 38236
rect 17083 38168 18828 38196
rect 18877 38199 18935 38205
rect 17083 38165 17095 38168
rect 17037 38159 17095 38165
rect 18877 38165 18889 38199
rect 18923 38196 18935 38199
rect 19242 38196 19248 38208
rect 18923 38168 19248 38196
rect 18923 38165 18935 38168
rect 18877 38159 18935 38165
rect 19242 38156 19248 38168
rect 19300 38156 19306 38208
rect 20732 38196 20760 38295
rect 20806 38292 20812 38344
rect 20864 38332 20870 38344
rect 21008 38341 21036 38440
rect 22646 38428 22652 38480
rect 22704 38468 22710 38480
rect 26712 38468 26740 38508
rect 26786 38496 26792 38548
rect 26844 38536 26850 38548
rect 26844 38508 28580 38536
rect 26844 38496 26850 38508
rect 27341 38471 27399 38477
rect 27341 38468 27353 38471
rect 22704 38440 26646 38468
rect 26712 38440 27353 38468
rect 22704 38428 22710 38440
rect 21542 38400 21548 38412
rect 21100 38372 21548 38400
rect 21100 38341 21128 38372
rect 21542 38360 21548 38372
rect 21600 38360 21606 38412
rect 22281 38403 22339 38409
rect 22281 38400 22293 38403
rect 21744 38372 22293 38400
rect 20993 38335 21051 38341
rect 20864 38304 20909 38332
rect 20864 38292 20870 38304
rect 20993 38301 21005 38335
rect 21039 38301 21051 38335
rect 20993 38295 21051 38301
rect 21085 38335 21143 38341
rect 21085 38301 21097 38335
rect 21131 38301 21143 38335
rect 21085 38295 21143 38301
rect 21223 38335 21281 38341
rect 21223 38301 21235 38335
rect 21269 38332 21281 38335
rect 21634 38332 21640 38344
rect 21269 38304 21640 38332
rect 21269 38301 21281 38304
rect 21223 38295 21281 38301
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 21450 38224 21456 38276
rect 21508 38264 21514 38276
rect 21744 38264 21772 38372
rect 22281 38369 22293 38372
rect 22327 38369 22339 38403
rect 22281 38363 22339 38369
rect 22738 38360 22744 38412
rect 22796 38360 22802 38412
rect 23768 38409 23796 38440
rect 23753 38403 23811 38409
rect 23753 38369 23765 38403
rect 23799 38369 23811 38403
rect 23753 38363 23811 38369
rect 24578 38360 24584 38412
rect 24636 38400 24642 38412
rect 26618 38400 26646 38440
rect 27341 38437 27353 38440
rect 27387 38468 27399 38471
rect 28350 38468 28356 38480
rect 27387 38440 28356 38468
rect 27387 38437 27399 38440
rect 27341 38431 27399 38437
rect 28350 38428 28356 38440
rect 28408 38428 28414 38480
rect 28552 38468 28580 38508
rect 28626 38496 28632 38548
rect 28684 38496 28690 38548
rect 29178 38496 29184 38548
rect 29236 38536 29242 38548
rect 29546 38536 29552 38548
rect 29236 38508 29552 38536
rect 29236 38496 29242 38508
rect 29546 38496 29552 38508
rect 29604 38496 29610 38548
rect 29730 38496 29736 38548
rect 29788 38496 29794 38548
rect 30558 38496 30564 38548
rect 30616 38496 30622 38548
rect 31110 38496 31116 38548
rect 31168 38536 31174 38548
rect 31297 38539 31355 38545
rect 31297 38536 31309 38539
rect 31168 38508 31309 38536
rect 31168 38496 31174 38508
rect 31297 38505 31309 38508
rect 31343 38505 31355 38539
rect 31297 38499 31355 38505
rect 32766 38496 32772 38548
rect 32824 38496 32830 38548
rect 35437 38539 35495 38545
rect 35437 38505 35449 38539
rect 35483 38536 35495 38539
rect 35618 38536 35624 38548
rect 35483 38508 35624 38536
rect 35483 38505 35495 38508
rect 35437 38499 35495 38505
rect 35618 38496 35624 38508
rect 35676 38496 35682 38548
rect 36446 38496 36452 38548
rect 36504 38536 36510 38548
rect 36633 38539 36691 38545
rect 36633 38536 36645 38539
rect 36504 38508 36645 38536
rect 36504 38496 36510 38508
rect 36633 38505 36645 38508
rect 36679 38505 36691 38539
rect 36633 38499 36691 38505
rect 38565 38539 38623 38545
rect 38565 38505 38577 38539
rect 38611 38536 38623 38539
rect 39206 38536 39212 38548
rect 38611 38508 39212 38536
rect 38611 38505 38623 38508
rect 38565 38499 38623 38505
rect 39206 38496 39212 38508
rect 39264 38496 39270 38548
rect 40313 38539 40371 38545
rect 40313 38505 40325 38539
rect 40359 38536 40371 38539
rect 41046 38536 41052 38548
rect 40359 38508 41052 38536
rect 40359 38505 40371 38508
rect 40313 38499 40371 38505
rect 41046 38496 41052 38508
rect 41104 38496 41110 38548
rect 29270 38468 29276 38480
rect 28552 38440 29276 38468
rect 29270 38428 29276 38440
rect 29328 38428 29334 38480
rect 33226 38468 33232 38480
rect 29564 38440 33232 38468
rect 29564 38400 29592 38440
rect 32784 38412 32812 38440
rect 33226 38428 33232 38440
rect 33284 38428 33290 38480
rect 34882 38428 34888 38480
rect 34940 38468 34946 38480
rect 40494 38468 40500 38480
rect 34940 38440 40500 38468
rect 34940 38428 34946 38440
rect 40494 38428 40500 38440
rect 40552 38428 40558 38480
rect 24636 38372 26556 38400
rect 26618 38372 29592 38400
rect 24636 38360 24642 38372
rect 21818 38292 21824 38344
rect 21876 38292 21882 38344
rect 22462 38292 22468 38344
rect 22520 38292 22526 38344
rect 24762 38341 24768 38344
rect 22833 38335 22891 38341
rect 22833 38301 22845 38335
rect 22879 38301 22891 38335
rect 23937 38335 23995 38341
rect 23937 38332 23949 38335
rect 22833 38295 22891 38301
rect 23493 38304 23949 38332
rect 21508 38236 21772 38264
rect 21508 38224 21514 38236
rect 22738 38224 22744 38276
rect 22796 38264 22802 38276
rect 22848 38264 22876 38295
rect 22796 38236 22876 38264
rect 22796 38224 22802 38236
rect 22002 38196 22008 38208
rect 20732 38168 22008 38196
rect 22002 38156 22008 38168
rect 22060 38196 22066 38208
rect 23198 38196 23204 38208
rect 22060 38168 23204 38196
rect 22060 38156 22066 38168
rect 23198 38156 23204 38168
rect 23256 38196 23262 38208
rect 23493 38196 23521 38304
rect 23937 38301 23949 38304
rect 23983 38301 23995 38335
rect 24760 38332 24768 38341
rect 24723 38304 24768 38332
rect 23937 38295 23995 38301
rect 24760 38295 24768 38304
rect 24762 38292 24768 38295
rect 24820 38292 24826 38344
rect 24964 38341 24992 38372
rect 24949 38335 25007 38341
rect 24949 38301 24961 38335
rect 24995 38301 25007 38335
rect 24949 38295 25007 38301
rect 25077 38335 25135 38341
rect 25077 38301 25089 38335
rect 25123 38301 25135 38335
rect 25077 38295 25135 38301
rect 25225 38335 25283 38341
rect 25225 38301 25237 38335
rect 25271 38332 25283 38335
rect 25866 38332 25872 38344
rect 25271 38304 25872 38332
rect 25271 38301 25283 38304
rect 25225 38295 25283 38301
rect 23750 38224 23756 38276
rect 23808 38264 23814 38276
rect 24857 38267 24915 38273
rect 24857 38264 24869 38267
rect 23808 38236 24869 38264
rect 23808 38224 23814 38236
rect 24857 38233 24869 38236
rect 24903 38233 24915 38267
rect 24857 38227 24915 38233
rect 23256 38168 23521 38196
rect 23256 38156 23262 38168
rect 23566 38156 23572 38208
rect 23624 38196 23630 38208
rect 25092 38196 25120 38295
rect 25866 38292 25872 38304
rect 25924 38292 25930 38344
rect 26234 38292 26240 38344
rect 26292 38332 26298 38344
rect 26375 38335 26433 38341
rect 26375 38332 26387 38335
rect 26292 38304 26387 38332
rect 26292 38292 26298 38304
rect 26375 38301 26387 38304
rect 26421 38301 26433 38335
rect 26528 38332 26556 38372
rect 29638 38360 29644 38412
rect 29696 38400 29702 38412
rect 31481 38403 31539 38409
rect 29696 38372 30972 38400
rect 29696 38360 29702 38372
rect 26528 38304 26648 38332
rect 26375 38295 26433 38301
rect 26620 38276 26648 38304
rect 26694 38292 26700 38344
rect 26752 38341 26758 38344
rect 26752 38335 26791 38341
rect 26779 38301 26791 38335
rect 26752 38295 26791 38301
rect 26881 38335 26939 38341
rect 26881 38301 26893 38335
rect 26927 38332 26939 38335
rect 26970 38332 26976 38344
rect 26927 38304 26976 38332
rect 26927 38301 26939 38304
rect 26881 38295 26939 38301
rect 26752 38292 26758 38295
rect 26970 38292 26976 38304
rect 27028 38332 27034 38344
rect 27982 38332 27988 38344
rect 27028 38304 27988 38332
rect 27028 38292 27034 38304
rect 27982 38292 27988 38304
rect 28040 38292 28046 38344
rect 28166 38341 28172 38344
rect 28133 38335 28172 38341
rect 28133 38301 28145 38335
rect 28133 38295 28172 38301
rect 28166 38292 28172 38295
rect 28224 38292 28230 38344
rect 28350 38292 28356 38344
rect 28408 38292 28414 38344
rect 28491 38335 28549 38341
rect 28491 38301 28503 38335
rect 28537 38332 28549 38335
rect 28626 38332 28632 38344
rect 28537 38304 28632 38332
rect 28537 38301 28549 38304
rect 28491 38295 28549 38301
rect 28626 38292 28632 38304
rect 28684 38332 28690 38344
rect 30834 38332 30840 38344
rect 28684 38304 30840 38332
rect 28684 38292 28690 38304
rect 30834 38292 30840 38304
rect 30892 38292 30898 38344
rect 26513 38267 26571 38273
rect 26513 38233 26525 38267
rect 26559 38233 26571 38267
rect 26513 38227 26571 38233
rect 23624 38168 25120 38196
rect 23624 38156 23630 38168
rect 25682 38156 25688 38208
rect 25740 38156 25746 38208
rect 26237 38199 26295 38205
rect 26237 38165 26249 38199
rect 26283 38196 26295 38199
rect 26326 38196 26332 38208
rect 26283 38168 26332 38196
rect 26283 38165 26295 38168
rect 26237 38159 26295 38165
rect 26326 38156 26332 38168
rect 26384 38156 26390 38208
rect 26528 38196 26556 38227
rect 26602 38224 26608 38276
rect 26660 38264 26666 38276
rect 28261 38267 28319 38273
rect 28261 38264 28273 38267
rect 26660 38236 28273 38264
rect 26660 38224 26666 38236
rect 28261 38233 28273 38236
rect 28307 38233 28319 38267
rect 28261 38227 28319 38233
rect 26878 38196 26884 38208
rect 26528 38168 26884 38196
rect 26878 38156 26884 38168
rect 26936 38156 26942 38208
rect 27890 38156 27896 38208
rect 27948 38196 27954 38208
rect 28166 38196 28172 38208
rect 27948 38168 28172 38196
rect 27948 38156 27954 38168
rect 28166 38156 28172 38168
rect 28224 38156 28230 38208
rect 28276 38196 28304 38227
rect 29914 38224 29920 38276
rect 29972 38224 29978 38276
rect 30101 38267 30159 38273
rect 30101 38233 30113 38267
rect 30147 38264 30159 38267
rect 30190 38264 30196 38276
rect 30147 38236 30196 38264
rect 30147 38233 30159 38236
rect 30101 38227 30159 38233
rect 30190 38224 30196 38236
rect 30248 38224 30254 38276
rect 30006 38196 30012 38208
rect 28276 38168 30012 38196
rect 30006 38156 30012 38168
rect 30064 38156 30070 38208
rect 30944 38196 30972 38372
rect 31481 38369 31493 38403
rect 31527 38400 31539 38403
rect 32306 38400 32312 38412
rect 31527 38372 32312 38400
rect 31527 38369 31539 38372
rect 31481 38363 31539 38369
rect 32306 38360 32312 38372
rect 32364 38360 32370 38412
rect 32766 38360 32772 38412
rect 32824 38360 32830 38412
rect 34146 38400 34152 38412
rect 33704 38372 34152 38400
rect 31018 38292 31024 38344
rect 31076 38332 31082 38344
rect 31665 38335 31723 38341
rect 31665 38332 31677 38335
rect 31076 38304 31677 38332
rect 31076 38292 31082 38304
rect 31665 38301 31677 38304
rect 31711 38301 31723 38335
rect 31665 38295 31723 38301
rect 31757 38335 31815 38341
rect 31757 38301 31769 38335
rect 31803 38301 31815 38335
rect 31757 38295 31815 38301
rect 31570 38224 31576 38276
rect 31628 38264 31634 38276
rect 31772 38264 31800 38295
rect 33318 38292 33324 38344
rect 33376 38292 33382 38344
rect 33410 38292 33416 38344
rect 33468 38292 33474 38344
rect 33704 38341 33732 38372
rect 34146 38360 34152 38372
rect 34204 38360 34210 38412
rect 39390 38400 39396 38412
rect 34440 38372 39396 38400
rect 34440 38344 34468 38372
rect 33689 38335 33747 38341
rect 33689 38301 33701 38335
rect 33735 38301 33747 38335
rect 33689 38295 33747 38301
rect 33781 38335 33839 38341
rect 33781 38301 33793 38335
rect 33827 38332 33839 38335
rect 34422 38332 34428 38344
rect 33827 38304 34428 38332
rect 33827 38301 33839 38304
rect 33781 38295 33839 38301
rect 31628 38236 31800 38264
rect 31628 38224 31634 38236
rect 32214 38224 32220 38276
rect 32272 38264 32278 38276
rect 33042 38264 33048 38276
rect 32272 38236 33048 38264
rect 32272 38224 32278 38236
rect 33042 38224 33048 38236
rect 33100 38224 33106 38276
rect 33226 38224 33232 38276
rect 33284 38264 33290 38276
rect 33796 38264 33824 38295
rect 34422 38292 34428 38304
rect 34480 38292 34486 38344
rect 34882 38292 34888 38344
rect 34940 38292 34946 38344
rect 35253 38335 35311 38341
rect 35253 38332 35265 38335
rect 34992 38304 35265 38332
rect 33284 38236 33824 38264
rect 33284 38224 33290 38236
rect 34514 38224 34520 38276
rect 34572 38264 34578 38276
rect 34992 38264 35020 38304
rect 35253 38301 35265 38304
rect 35299 38332 35311 38335
rect 36814 38332 36820 38344
rect 35299 38304 36820 38332
rect 35299 38301 35311 38304
rect 35253 38295 35311 38301
rect 36814 38292 36820 38304
rect 36872 38292 36878 38344
rect 37016 38341 37044 38372
rect 39390 38360 39396 38372
rect 39448 38360 39454 38412
rect 41046 38360 41052 38412
rect 41104 38360 41110 38412
rect 41509 38403 41567 38409
rect 41509 38369 41521 38403
rect 41555 38400 41567 38403
rect 41555 38372 42104 38400
rect 41555 38369 41567 38372
rect 41509 38363 41567 38369
rect 37001 38335 37059 38341
rect 37001 38301 37013 38335
rect 37047 38301 37059 38335
rect 37001 38295 37059 38301
rect 37090 38292 37096 38344
rect 37148 38292 37154 38344
rect 37366 38292 37372 38344
rect 37424 38292 37430 38344
rect 37642 38292 37648 38344
rect 37700 38292 37706 38344
rect 37826 38292 37832 38344
rect 37884 38292 37890 38344
rect 40034 38292 40040 38344
rect 40092 38292 40098 38344
rect 40126 38292 40132 38344
rect 40184 38292 40190 38344
rect 41138 38292 41144 38344
rect 41196 38292 41202 38344
rect 41874 38292 41880 38344
rect 41932 38332 41938 38344
rect 41969 38335 42027 38341
rect 41969 38332 41981 38335
rect 41932 38304 41981 38332
rect 41932 38292 41938 38304
rect 41969 38301 41981 38304
rect 42015 38301 42027 38335
rect 42076 38332 42104 38372
rect 42225 38335 42283 38341
rect 42225 38332 42237 38335
rect 42076 38304 42237 38332
rect 41969 38295 42027 38301
rect 42225 38301 42237 38304
rect 42271 38301 42283 38335
rect 42225 38295 42283 38301
rect 34572 38236 35020 38264
rect 34572 38224 34578 38236
rect 35066 38224 35072 38276
rect 35124 38224 35130 38276
rect 35158 38224 35164 38276
rect 35216 38224 35222 38276
rect 35820 38236 36860 38264
rect 35820 38196 35848 38236
rect 30944 38168 35848 38196
rect 35986 38156 35992 38208
rect 36044 38196 36050 38208
rect 36630 38196 36636 38208
rect 36044 38168 36636 38196
rect 36044 38156 36050 38168
rect 36630 38156 36636 38168
rect 36688 38156 36694 38208
rect 36832 38196 36860 38236
rect 36998 38196 37004 38208
rect 36832 38168 37004 38196
rect 36998 38156 37004 38168
rect 37056 38156 37062 38208
rect 37660 38196 37688 38292
rect 37918 38224 37924 38276
rect 37976 38264 37982 38276
rect 39025 38267 39083 38273
rect 39025 38264 39037 38267
rect 37976 38236 39037 38264
rect 37976 38224 37982 38236
rect 39025 38233 39037 38236
rect 39071 38233 39083 38267
rect 39025 38227 39083 38233
rect 40313 38267 40371 38273
rect 40313 38233 40325 38267
rect 40359 38264 40371 38267
rect 40678 38264 40684 38276
rect 40359 38236 40684 38264
rect 40359 38233 40371 38236
rect 40313 38227 40371 38233
rect 40678 38224 40684 38236
rect 40736 38224 40742 38276
rect 38470 38196 38476 38208
rect 37660 38168 38476 38196
rect 38470 38156 38476 38168
rect 38528 38156 38534 38208
rect 39850 38156 39856 38208
rect 39908 38196 39914 38208
rect 43349 38199 43407 38205
rect 43349 38196 43361 38199
rect 39908 38168 43361 38196
rect 39908 38156 39914 38168
rect 43349 38165 43361 38168
rect 43395 38165 43407 38199
rect 43349 38159 43407 38165
rect 1104 38106 43884 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 43884 38106
rect 1104 38032 43884 38054
rect 18230 37952 18236 38004
rect 18288 37952 18294 38004
rect 18877 37995 18935 38001
rect 18877 37961 18889 37995
rect 18923 37961 18935 37995
rect 18877 37955 18935 37961
rect 15194 37884 15200 37936
rect 15252 37884 15258 37936
rect 18417 37859 18475 37865
rect 18417 37825 18429 37859
rect 18463 37856 18475 37859
rect 18892 37856 18920 37955
rect 19242 37952 19248 38004
rect 19300 37992 19306 38004
rect 19300 37964 22324 37992
rect 19300 37952 19306 37964
rect 22296 37936 22324 37964
rect 23934 37952 23940 38004
rect 23992 37992 23998 38004
rect 24670 37992 24676 38004
rect 23992 37964 24676 37992
rect 23992 37952 23998 37964
rect 24670 37952 24676 37964
rect 24728 37952 24734 38004
rect 25130 37952 25136 38004
rect 25188 37952 25194 38004
rect 26602 37992 26608 38004
rect 25240 37964 25406 37992
rect 20162 37884 20168 37936
rect 20220 37924 20226 37936
rect 20257 37927 20315 37933
rect 20257 37924 20269 37927
rect 20220 37896 20269 37924
rect 20220 37884 20226 37896
rect 20257 37893 20269 37896
rect 20303 37893 20315 37927
rect 20257 37887 20315 37893
rect 20806 37884 20812 37936
rect 20864 37924 20870 37936
rect 21082 37924 21088 37936
rect 20864 37896 21088 37924
rect 20864 37884 20870 37896
rect 21082 37884 21088 37896
rect 21140 37884 21146 37936
rect 22278 37884 22284 37936
rect 22336 37884 22342 37936
rect 22373 37927 22431 37933
rect 22373 37893 22385 37927
rect 22419 37924 22431 37927
rect 23106 37924 23112 37936
rect 22419 37896 23112 37924
rect 22419 37893 22431 37896
rect 22373 37887 22431 37893
rect 23106 37884 23112 37896
rect 23164 37924 23170 37936
rect 23164 37896 23244 37924
rect 23164 37884 23170 37896
rect 18463 37828 18920 37856
rect 18463 37825 18475 37828
rect 18417 37819 18475 37825
rect 20898 37816 20904 37868
rect 20956 37816 20962 37868
rect 21266 37816 21272 37868
rect 21324 37816 21330 37868
rect 21450 37816 21456 37868
rect 21508 37816 21514 37868
rect 22094 37816 22100 37868
rect 22152 37865 22158 37868
rect 22152 37859 22201 37865
rect 22152 37825 22155 37859
rect 22189 37825 22201 37859
rect 22501 37859 22559 37865
rect 22501 37856 22513 37859
rect 22152 37819 22201 37825
rect 22480 37825 22513 37856
rect 22547 37825 22559 37859
rect 22480 37819 22559 37825
rect 22152 37816 22158 37819
rect 18506 37748 18512 37800
rect 18564 37788 18570 37800
rect 19242 37788 19248 37800
rect 18564 37760 19248 37788
rect 18564 37748 18570 37760
rect 19242 37748 19248 37760
rect 19300 37788 19306 37800
rect 19337 37791 19395 37797
rect 19337 37788 19349 37791
rect 19300 37760 19349 37788
rect 19300 37748 19306 37760
rect 19337 37757 19349 37760
rect 19383 37757 19395 37791
rect 19337 37751 19395 37757
rect 19426 37748 19432 37800
rect 19484 37748 19490 37800
rect 20990 37748 20996 37800
rect 21048 37748 21054 37800
rect 22480 37788 22508 37819
rect 22646 37816 22652 37868
rect 22704 37816 22710 37868
rect 23216 37856 23244 37896
rect 23290 37884 23296 37936
rect 23348 37924 23354 37936
rect 23569 37927 23627 37933
rect 23569 37924 23581 37927
rect 23348 37896 23581 37924
rect 23348 37884 23354 37896
rect 23569 37893 23581 37896
rect 23615 37893 23627 37927
rect 23569 37887 23627 37893
rect 23216 37828 23612 37856
rect 23584 37800 23612 37828
rect 24210 37816 24216 37868
rect 24268 37816 24274 37868
rect 24581 37859 24639 37865
rect 24581 37825 24593 37859
rect 24627 37856 24639 37859
rect 24670 37856 24676 37868
rect 24627 37828 24676 37856
rect 24627 37825 24639 37828
rect 24581 37819 24639 37825
rect 24670 37816 24676 37828
rect 24728 37816 24734 37868
rect 24762 37816 24768 37868
rect 24820 37816 24826 37868
rect 23290 37788 23296 37800
rect 21376 37760 23296 37788
rect 21376 37732 21404 37760
rect 23290 37748 23296 37760
rect 23348 37748 23354 37800
rect 23566 37748 23572 37800
rect 23624 37748 23630 37800
rect 24026 37748 24032 37800
rect 24084 37748 24090 37800
rect 15749 37723 15807 37729
rect 15749 37689 15761 37723
rect 15795 37720 15807 37723
rect 17218 37720 17224 37732
rect 15795 37692 17224 37720
rect 15795 37689 15807 37692
rect 15749 37683 15807 37689
rect 17218 37680 17224 37692
rect 17276 37680 17282 37732
rect 17773 37723 17831 37729
rect 17773 37689 17785 37723
rect 17819 37720 17831 37723
rect 21358 37720 21364 37732
rect 17819 37692 21364 37720
rect 17819 37689 17831 37692
rect 17773 37683 17831 37689
rect 21358 37680 21364 37692
rect 21416 37680 21422 37732
rect 25148 37720 25176 37952
rect 25240 37868 25268 37964
rect 25378 37924 25406 37964
rect 25608 37964 26608 37992
rect 25608 37933 25636 37964
rect 26602 37952 26608 37964
rect 26660 37952 26666 38004
rect 27264 37964 28064 37992
rect 25501 37927 25559 37933
rect 25501 37924 25513 37927
rect 25378 37896 25513 37924
rect 25501 37893 25513 37896
rect 25547 37893 25559 37927
rect 25501 37887 25559 37893
rect 25593 37927 25651 37933
rect 25593 37893 25605 37927
rect 25639 37893 25651 37927
rect 25593 37887 25651 37893
rect 26326 37884 26332 37936
rect 26384 37884 26390 37936
rect 27264 37924 27292 37964
rect 26436 37896 27292 37924
rect 25222 37816 25228 37868
rect 25280 37816 25286 37868
rect 25404 37859 25462 37865
rect 25404 37856 25416 37859
rect 25332 37828 25416 37856
rect 25332 37788 25360 37828
rect 25404 37825 25416 37828
rect 25450 37825 25462 37859
rect 25404 37819 25462 37825
rect 25682 37816 25688 37868
rect 25740 37865 25746 37868
rect 25740 37859 25779 37865
rect 25767 37825 25779 37859
rect 25740 37819 25779 37825
rect 25740 37816 25746 37819
rect 25866 37816 25872 37868
rect 25924 37816 25930 37868
rect 26142 37816 26148 37868
rect 26200 37856 26206 37868
rect 26436 37856 26464 37896
rect 26200 37828 26464 37856
rect 26513 37859 26571 37865
rect 26200 37816 26206 37828
rect 26513 37825 26525 37859
rect 26559 37825 26571 37859
rect 26513 37819 26571 37825
rect 26605 37859 26663 37865
rect 26605 37825 26617 37859
rect 26651 37856 26663 37859
rect 26786 37856 26792 37868
rect 26651 37828 26792 37856
rect 26651 37825 26663 37828
rect 26605 37819 26663 37825
rect 26234 37788 26240 37800
rect 25332 37760 26240 37788
rect 26234 37748 26240 37760
rect 26292 37748 26298 37800
rect 26528 37788 26556 37819
rect 26786 37816 26792 37828
rect 26844 37816 26850 37868
rect 27264 37865 27292 37896
rect 27617 37927 27675 37933
rect 27617 37893 27629 37927
rect 27663 37924 27675 37927
rect 27890 37924 27896 37936
rect 27663 37896 27896 37924
rect 27663 37893 27675 37896
rect 27617 37887 27675 37893
rect 27890 37884 27896 37896
rect 27948 37884 27954 37936
rect 27430 37865 27436 37868
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 27397 37859 27436 37865
rect 27397 37825 27409 37859
rect 27397 37819 27436 37825
rect 27430 37816 27436 37819
rect 27488 37816 27494 37868
rect 27522 37816 27528 37868
rect 27580 37816 27586 37868
rect 27755 37859 27813 37865
rect 27755 37825 27767 37859
rect 27801 37825 27813 37859
rect 28036 37862 28064 37964
rect 28644 37964 30512 37992
rect 28644 37936 28672 37964
rect 28626 37884 28632 37936
rect 28684 37884 28690 37936
rect 28721 37927 28779 37933
rect 28721 37893 28733 37927
rect 28767 37924 28779 37927
rect 30374 37924 30380 37936
rect 28767 37896 30380 37924
rect 28767 37893 28779 37896
rect 28721 37887 28779 37893
rect 30374 37884 30380 37896
rect 30432 37884 30438 37936
rect 30484 37924 30512 37964
rect 30558 37952 30564 38004
rect 30616 37992 30622 38004
rect 30653 37995 30711 38001
rect 30653 37992 30665 37995
rect 30616 37964 30665 37992
rect 30616 37952 30622 37964
rect 30653 37961 30665 37964
rect 30699 37961 30711 37995
rect 30653 37955 30711 37961
rect 30742 37952 30748 38004
rect 30800 37952 30806 38004
rect 31754 37952 31760 38004
rect 31812 37952 31818 38004
rect 32306 37952 32312 38004
rect 32364 37952 32370 38004
rect 34517 37995 34575 38001
rect 32600 37964 34284 37992
rect 30760 37924 30788 37952
rect 32398 37924 32404 37936
rect 30484 37896 30788 37924
rect 31588 37896 32404 37924
rect 28036 37846 28120 37862
rect 28353 37859 28411 37865
rect 28353 37856 28365 37859
rect 28276 37846 28365 37856
rect 28036 37834 28365 37846
rect 27755 37819 27813 37825
rect 28092 37828 28365 37834
rect 26528 37760 27292 37788
rect 27264 37732 27292 37760
rect 25225 37723 25283 37729
rect 25225 37720 25237 37723
rect 25148 37692 25237 37720
rect 25225 37689 25237 37692
rect 25271 37689 25283 37723
rect 25225 37683 25283 37689
rect 26329 37723 26387 37729
rect 26329 37689 26341 37723
rect 26375 37720 26387 37723
rect 26510 37720 26516 37732
rect 26375 37692 26516 37720
rect 26375 37689 26387 37692
rect 26329 37683 26387 37689
rect 26510 37680 26516 37692
rect 26568 37680 26574 37732
rect 27246 37680 27252 37732
rect 27304 37680 27310 37732
rect 27338 37680 27344 37732
rect 27396 37720 27402 37732
rect 27770 37720 27798 37819
rect 28092 37818 28304 37828
rect 28353 37825 28365 37828
rect 28399 37825 28411 37859
rect 28353 37819 28411 37825
rect 28442 37816 28448 37868
rect 28500 37865 28506 37868
rect 28500 37859 28531 37865
rect 28519 37825 28531 37859
rect 28500 37819 28531 37825
rect 28500 37816 28506 37819
rect 28810 37816 28816 37868
rect 28868 37865 28874 37868
rect 28868 37856 28876 37865
rect 29641 37859 29699 37865
rect 28868 37828 28913 37856
rect 28868 37819 28876 37828
rect 29641 37825 29653 37859
rect 29687 37825 29699 37859
rect 29641 37819 29699 37825
rect 28868 37816 28874 37819
rect 27982 37748 27988 37800
rect 28040 37788 28046 37800
rect 29178 37788 29184 37800
rect 28040 37760 29184 37788
rect 28040 37748 28046 37760
rect 29178 37748 29184 37760
rect 29236 37748 29242 37800
rect 27396 37692 28028 37720
rect 27396 37680 27402 37692
rect 16206 37612 16212 37664
rect 16264 37612 16270 37664
rect 17126 37612 17132 37664
rect 17184 37612 17190 37664
rect 21910 37612 21916 37664
rect 21968 37652 21974 37664
rect 22005 37655 22063 37661
rect 22005 37652 22017 37655
rect 21968 37624 22017 37652
rect 21968 37612 21974 37624
rect 22005 37621 22017 37624
rect 22051 37621 22063 37655
rect 22005 37615 22063 37621
rect 22554 37612 22560 37664
rect 22612 37652 22618 37664
rect 26878 37652 26884 37664
rect 22612 37624 26884 37652
rect 22612 37612 22618 37624
rect 26878 37612 26884 37624
rect 26936 37652 26942 37664
rect 27706 37652 27712 37664
rect 26936 37624 27712 37652
rect 26936 37612 26942 37624
rect 27706 37612 27712 37624
rect 27764 37612 27770 37664
rect 27890 37612 27896 37664
rect 27948 37612 27954 37664
rect 28000 37652 28028 37692
rect 28166 37680 28172 37732
rect 28224 37720 28230 37732
rect 29656 37720 29684 37819
rect 30466 37816 30472 37868
rect 30524 37816 30530 37868
rect 30650 37816 30656 37868
rect 30708 37856 30714 37868
rect 30745 37859 30803 37865
rect 30745 37856 30757 37859
rect 30708 37828 30757 37856
rect 30708 37816 30714 37828
rect 30745 37825 30757 37828
rect 30791 37825 30803 37859
rect 30745 37819 30803 37825
rect 31205 37859 31263 37865
rect 31205 37825 31217 37859
rect 31251 37825 31263 37859
rect 31205 37819 31263 37825
rect 31389 37859 31447 37865
rect 31389 37825 31401 37859
rect 31435 37825 31447 37859
rect 31389 37819 31447 37825
rect 29730 37748 29736 37800
rect 29788 37788 29794 37800
rect 30190 37788 30196 37800
rect 29788 37760 30196 37788
rect 29788 37748 29794 37760
rect 30190 37748 30196 37760
rect 30248 37748 30254 37800
rect 29914 37720 29920 37732
rect 28224 37692 29592 37720
rect 29656 37692 29920 37720
rect 28224 37680 28230 37692
rect 28810 37652 28816 37664
rect 28000 37624 28816 37652
rect 28810 37612 28816 37624
rect 28868 37612 28874 37664
rect 28994 37612 29000 37664
rect 29052 37612 29058 37664
rect 29564 37652 29592 37692
rect 29914 37680 29920 37692
rect 29972 37720 29978 37732
rect 30469 37723 30527 37729
rect 30469 37720 30481 37723
rect 29972 37692 30481 37720
rect 29972 37680 29978 37692
rect 30469 37689 30481 37692
rect 30515 37689 30527 37723
rect 31220 37720 31248 37819
rect 31404 37788 31432 37819
rect 31478 37816 31484 37868
rect 31536 37816 31542 37868
rect 31588 37865 31616 37896
rect 32398 37884 32404 37896
rect 32456 37884 32462 37936
rect 32600 37868 32628 37964
rect 34256 37933 34284 37964
rect 34517 37961 34529 37995
rect 34563 37992 34575 37995
rect 34563 37964 34928 37992
rect 34563 37961 34575 37964
rect 34517 37955 34575 37961
rect 34241 37927 34299 37933
rect 34241 37893 34253 37927
rect 34287 37924 34299 37927
rect 34698 37924 34704 37936
rect 34287 37896 34704 37924
rect 34287 37893 34299 37896
rect 34241 37887 34299 37893
rect 34698 37884 34704 37896
rect 34756 37884 34762 37936
rect 31573 37859 31631 37865
rect 31573 37825 31585 37859
rect 31619 37825 31631 37859
rect 31573 37819 31631 37825
rect 32493 37859 32551 37865
rect 32493 37825 32505 37859
rect 32539 37825 32551 37859
rect 32493 37819 32551 37825
rect 32508 37788 32536 37819
rect 32582 37816 32588 37868
rect 32640 37816 32646 37868
rect 32766 37816 32772 37868
rect 32824 37816 32830 37868
rect 32858 37816 32864 37868
rect 32916 37816 32922 37868
rect 33594 37816 33600 37868
rect 33652 37856 33658 37868
rect 33873 37859 33931 37865
rect 33873 37856 33885 37859
rect 33652 37828 33885 37856
rect 33652 37816 33658 37828
rect 33873 37825 33885 37828
rect 33919 37825 33931 37859
rect 33873 37819 33931 37825
rect 33962 37816 33968 37868
rect 34020 37856 34026 37868
rect 34020 37828 34065 37856
rect 34020 37816 34026 37828
rect 34146 37816 34152 37868
rect 34204 37816 34210 37868
rect 34422 37865 34428 37868
rect 34379 37859 34428 37865
rect 34379 37825 34391 37859
rect 34425 37825 34428 37859
rect 34379 37819 34428 37825
rect 34422 37816 34428 37819
rect 34480 37816 34486 37868
rect 34900 37856 34928 37964
rect 35250 37952 35256 38004
rect 35308 37952 35314 38004
rect 35805 37995 35863 38001
rect 35805 37961 35817 37995
rect 35851 37992 35863 37995
rect 36078 37992 36084 38004
rect 35851 37964 36084 37992
rect 35851 37961 35863 37964
rect 35805 37955 35863 37961
rect 36078 37952 36084 37964
rect 36136 37952 36142 38004
rect 36817 37995 36875 38001
rect 36817 37961 36829 37995
rect 36863 37992 36875 37995
rect 37366 37992 37372 38004
rect 36863 37964 37372 37992
rect 36863 37961 36875 37964
rect 36817 37955 36875 37961
rect 37366 37952 37372 37964
rect 37424 37952 37430 38004
rect 39022 37992 39028 38004
rect 38212 37964 39028 37992
rect 35268 37865 35296 37952
rect 35161 37859 35219 37865
rect 35161 37856 35173 37859
rect 34900 37828 35173 37856
rect 35161 37825 35173 37828
rect 35207 37825 35219 37859
rect 35268 37859 35339 37865
rect 35268 37828 35293 37859
rect 35161 37819 35219 37825
rect 35281 37825 35293 37828
rect 35327 37825 35339 37859
rect 35281 37819 35339 37825
rect 35437 37859 35495 37865
rect 35437 37825 35449 37859
rect 35483 37825 35495 37859
rect 35437 37819 35495 37825
rect 35452 37788 35480 37819
rect 35526 37816 35532 37868
rect 35584 37816 35590 37868
rect 35667 37859 35725 37865
rect 35667 37825 35679 37859
rect 35713 37856 35725 37859
rect 35894 37856 35900 37868
rect 35713 37828 35900 37856
rect 35713 37825 35725 37828
rect 35667 37819 35725 37825
rect 35894 37816 35900 37828
rect 35952 37816 35958 37868
rect 36265 37859 36323 37865
rect 36265 37825 36277 37859
rect 36311 37825 36323 37859
rect 36265 37819 36323 37825
rect 35802 37788 35808 37800
rect 31404 37760 35112 37788
rect 35452 37760 35808 37788
rect 35084 37732 35112 37760
rect 35802 37748 35808 37760
rect 35860 37748 35866 37800
rect 36280 37788 36308 37819
rect 36446 37816 36452 37868
rect 36504 37816 36510 37868
rect 36538 37816 36544 37868
rect 36596 37816 36602 37868
rect 36633 37859 36691 37865
rect 36633 37825 36645 37859
rect 36679 37856 36691 37859
rect 36814 37856 36820 37868
rect 36679 37828 36820 37856
rect 36679 37825 36691 37828
rect 36633 37819 36691 37825
rect 36814 37816 36820 37828
rect 36872 37816 36878 37868
rect 36998 37816 37004 37868
rect 37056 37856 37062 37868
rect 38212 37865 38240 37964
rect 39022 37952 39028 37964
rect 39080 37952 39086 38004
rect 39482 37952 39488 38004
rect 39540 37952 39546 38004
rect 40034 37952 40040 38004
rect 40092 37992 40098 38004
rect 40681 37995 40739 38001
rect 40681 37992 40693 37995
rect 40092 37964 40693 37992
rect 40092 37952 40098 37964
rect 40681 37961 40693 37964
rect 40727 37961 40739 37995
rect 40681 37955 40739 37961
rect 40405 37927 40463 37933
rect 40405 37893 40417 37927
rect 40451 37924 40463 37927
rect 40954 37924 40960 37936
rect 40451 37896 40960 37924
rect 40451 37893 40463 37896
rect 40405 37887 40463 37893
rect 40954 37884 40960 37896
rect 41012 37884 41018 37936
rect 41138 37884 41144 37936
rect 41196 37884 41202 37936
rect 41322 37884 41328 37936
rect 41380 37933 41386 37936
rect 41380 37927 41399 37933
rect 41387 37893 41399 37927
rect 41380 37887 41399 37893
rect 41380 37884 41386 37887
rect 38197 37859 38255 37865
rect 38197 37856 38209 37859
rect 37056 37828 38209 37856
rect 37056 37816 37062 37828
rect 38197 37825 38209 37828
rect 38243 37825 38255 37859
rect 38197 37819 38255 37825
rect 38470 37816 38476 37868
rect 38528 37816 38534 37868
rect 38749 37859 38807 37865
rect 38749 37825 38761 37859
rect 38795 37825 38807 37859
rect 38749 37819 38807 37825
rect 36722 37788 36728 37800
rect 36280 37760 36728 37788
rect 36722 37748 36728 37760
rect 36780 37748 36786 37800
rect 36906 37748 36912 37800
rect 36964 37788 36970 37800
rect 38764 37788 38792 37819
rect 39022 37816 39028 37868
rect 39080 37816 39086 37868
rect 39117 37859 39175 37865
rect 39117 37825 39129 37859
rect 39163 37856 39175 37859
rect 39390 37856 39396 37868
rect 39163 37828 39396 37856
rect 39163 37825 39175 37828
rect 39117 37819 39175 37825
rect 39390 37816 39396 37828
rect 39448 37816 39454 37868
rect 40034 37816 40040 37868
rect 40092 37816 40098 37868
rect 40185 37859 40243 37865
rect 40185 37825 40197 37859
rect 40231 37856 40243 37859
rect 40231 37825 40264 37856
rect 40185 37819 40264 37825
rect 36964 37760 38792 37788
rect 40236 37788 40264 37819
rect 40310 37816 40316 37868
rect 40368 37816 40374 37868
rect 40586 37865 40592 37868
rect 40543 37859 40592 37865
rect 40543 37825 40555 37859
rect 40589 37825 40592 37859
rect 40543 37819 40592 37825
rect 40586 37816 40592 37819
rect 40644 37816 40650 37868
rect 40402 37788 40408 37800
rect 40236 37760 40408 37788
rect 36964 37748 36970 37760
rect 40402 37748 40408 37760
rect 40460 37748 40466 37800
rect 40770 37748 40776 37800
rect 40828 37788 40834 37800
rect 41969 37791 42027 37797
rect 41969 37788 41981 37791
rect 40828 37760 41981 37788
rect 40828 37748 40834 37760
rect 41969 37757 41981 37760
rect 42015 37757 42027 37791
rect 41969 37751 42027 37757
rect 32214 37720 32220 37732
rect 31220 37692 32220 37720
rect 30469 37683 30527 37689
rect 32214 37680 32220 37692
rect 32272 37680 32278 37732
rect 33413 37723 33471 37729
rect 33413 37689 33425 37723
rect 33459 37720 33471 37723
rect 34790 37720 34796 37732
rect 33459 37692 34796 37720
rect 33459 37689 33471 37692
rect 33413 37683 33471 37689
rect 29822 37652 29828 37664
rect 29564 37624 29828 37652
rect 29822 37612 29828 37624
rect 29880 37612 29886 37664
rect 30006 37612 30012 37664
rect 30064 37612 30070 37664
rect 31202 37612 31208 37664
rect 31260 37652 31266 37664
rect 33428 37652 33456 37683
rect 34790 37680 34796 37692
rect 34848 37680 34854 37732
rect 35066 37680 35072 37732
rect 35124 37720 35130 37732
rect 36446 37720 36452 37732
rect 35124 37692 36452 37720
rect 35124 37680 35130 37692
rect 36446 37680 36452 37692
rect 36504 37680 36510 37732
rect 38194 37720 38200 37732
rect 36556 37692 38200 37720
rect 31260 37624 33456 37652
rect 31260 37612 31266 37624
rect 33502 37612 33508 37664
rect 33560 37652 33566 37664
rect 34514 37652 34520 37664
rect 33560 37624 34520 37652
rect 33560 37612 33566 37624
rect 34514 37612 34520 37624
rect 34572 37612 34578 37664
rect 34698 37612 34704 37664
rect 34756 37652 34762 37664
rect 36556 37652 36584 37692
rect 38194 37680 38200 37692
rect 38252 37720 38258 37732
rect 43165 37723 43223 37729
rect 43165 37720 43177 37723
rect 38252 37692 40448 37720
rect 38252 37680 38258 37692
rect 34756 37624 36584 37652
rect 34756 37612 34762 37624
rect 36630 37612 36636 37664
rect 36688 37652 36694 37664
rect 37553 37655 37611 37661
rect 37553 37652 37565 37655
rect 36688 37624 37565 37652
rect 36688 37612 36694 37624
rect 37553 37621 37565 37624
rect 37599 37652 37611 37655
rect 39206 37652 39212 37664
rect 37599 37624 39212 37652
rect 37599 37621 37611 37624
rect 37553 37615 37611 37621
rect 39206 37612 39212 37624
rect 39264 37612 39270 37664
rect 40420 37652 40448 37692
rect 40604 37692 43177 37720
rect 40604 37652 40632 37692
rect 43165 37689 43177 37692
rect 43211 37689 43223 37723
rect 43165 37683 43223 37689
rect 40420 37624 40632 37652
rect 41138 37612 41144 37664
rect 41196 37652 41202 37664
rect 41325 37655 41383 37661
rect 41325 37652 41337 37655
rect 41196 37624 41337 37652
rect 41196 37612 41202 37624
rect 41325 37621 41337 37624
rect 41371 37621 41383 37655
rect 41325 37615 41383 37621
rect 41506 37612 41512 37664
rect 41564 37612 41570 37664
rect 42058 37612 42064 37664
rect 42116 37652 42122 37664
rect 42613 37655 42671 37661
rect 42613 37652 42625 37655
rect 42116 37624 42625 37652
rect 42116 37612 42122 37624
rect 42613 37621 42625 37624
rect 42659 37621 42671 37655
rect 42613 37615 42671 37621
rect 1104 37562 43884 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 43884 37562
rect 1104 37488 43884 37510
rect 14458 37408 14464 37460
rect 14516 37408 14522 37460
rect 15562 37408 15568 37460
rect 15620 37408 15626 37460
rect 16114 37408 16120 37460
rect 16172 37408 16178 37460
rect 16666 37408 16672 37460
rect 16724 37408 16730 37460
rect 17218 37408 17224 37460
rect 17276 37408 17282 37460
rect 17770 37408 17776 37460
rect 17828 37448 17834 37460
rect 23934 37448 23940 37460
rect 17828 37420 23940 37448
rect 17828 37408 17834 37420
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 24029 37451 24087 37457
rect 24029 37417 24041 37451
rect 24075 37417 24087 37451
rect 24029 37411 24087 37417
rect 15013 37383 15071 37389
rect 15013 37349 15025 37383
rect 15059 37380 15071 37383
rect 16574 37380 16580 37392
rect 15059 37352 16580 37380
rect 15059 37349 15071 37352
rect 15013 37343 15071 37349
rect 16574 37340 16580 37352
rect 16632 37340 16638 37392
rect 18325 37383 18383 37389
rect 18325 37349 18337 37383
rect 18371 37380 18383 37383
rect 18877 37383 18935 37389
rect 18877 37380 18889 37383
rect 18371 37352 18889 37380
rect 18371 37349 18383 37352
rect 18325 37343 18383 37349
rect 18877 37349 18889 37352
rect 18923 37380 18935 37383
rect 19426 37380 19432 37392
rect 18923 37352 19432 37380
rect 18923 37349 18935 37352
rect 18877 37343 18935 37349
rect 19426 37340 19432 37352
rect 19484 37380 19490 37392
rect 20070 37380 20076 37392
rect 19484 37352 20076 37380
rect 19484 37340 19490 37352
rect 20070 37340 20076 37352
rect 20128 37340 20134 37392
rect 21266 37340 21272 37392
rect 21324 37380 21330 37392
rect 22646 37380 22652 37392
rect 21324 37352 22652 37380
rect 21324 37340 21330 37352
rect 16206 37272 16212 37324
rect 16264 37312 16270 37324
rect 20809 37315 20867 37321
rect 20809 37312 20821 37315
rect 16264 37284 20821 37312
rect 16264 37272 16270 37284
rect 20809 37281 20821 37284
rect 20855 37281 20867 37315
rect 20809 37275 20867 37281
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19392 37216 19625 37244
rect 19392 37204 19398 37216
rect 19613 37213 19625 37216
rect 19659 37213 19671 37247
rect 20824 37244 20852 37275
rect 21910 37272 21916 37324
rect 21968 37272 21974 37324
rect 22005 37247 22063 37253
rect 20824 37216 21956 37244
rect 19613 37207 19671 37213
rect 19242 37136 19248 37188
rect 19300 37176 19306 37188
rect 21361 37179 21419 37185
rect 21361 37176 21373 37179
rect 19300 37148 21373 37176
rect 19300 37136 19306 37148
rect 21361 37145 21373 37148
rect 21407 37145 21419 37179
rect 21928 37176 21956 37216
rect 22005 37213 22017 37247
rect 22051 37244 22063 37247
rect 22186 37244 22192 37256
rect 22051 37216 22192 37244
rect 22051 37213 22063 37216
rect 22005 37207 22063 37213
rect 22186 37204 22192 37216
rect 22244 37204 22250 37256
rect 22388 37253 22416 37352
rect 22646 37340 22652 37352
rect 22704 37340 22710 37392
rect 24044 37324 24072 37411
rect 24118 37408 24124 37460
rect 24176 37448 24182 37460
rect 25682 37448 25688 37460
rect 24176 37420 25688 37448
rect 24176 37408 24182 37420
rect 25682 37408 25688 37420
rect 25740 37408 25746 37460
rect 25866 37408 25872 37460
rect 25924 37448 25930 37460
rect 27522 37448 27528 37460
rect 25924 37420 27528 37448
rect 25924 37408 25930 37420
rect 27522 37408 27528 37420
rect 27580 37448 27586 37460
rect 28626 37448 28632 37460
rect 27580 37420 28632 37448
rect 27580 37408 27586 37420
rect 28626 37408 28632 37420
rect 28684 37408 28690 37460
rect 31018 37448 31024 37460
rect 29196 37420 31024 37448
rect 26326 37380 26332 37392
rect 24688 37352 26332 37380
rect 22480 37284 23521 37312
rect 22373 37247 22431 37253
rect 22373 37213 22385 37247
rect 22419 37213 22431 37247
rect 22373 37207 22431 37213
rect 22480 37176 22508 37284
rect 23493 37256 23521 37284
rect 24026 37272 24032 37324
rect 24084 37272 24090 37324
rect 24302 37272 24308 37324
rect 24360 37312 24366 37324
rect 24578 37312 24584 37324
rect 24360 37284 24584 37312
rect 24360 37272 24366 37284
rect 24578 37272 24584 37284
rect 24636 37272 24642 37324
rect 22557 37247 22615 37253
rect 22557 37213 22569 37247
rect 22603 37244 22615 37247
rect 23106 37244 23112 37256
rect 22603 37216 23112 37244
rect 22603 37213 22615 37216
rect 22557 37207 22615 37213
rect 21928 37148 22508 37176
rect 21361 37139 21419 37145
rect 19426 37068 19432 37120
rect 19484 37068 19490 37120
rect 20254 37068 20260 37120
rect 20312 37068 20318 37120
rect 22370 37068 22376 37120
rect 22428 37108 22434 37120
rect 22572 37108 22600 37207
rect 23106 37204 23112 37216
rect 23164 37204 23170 37256
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23256 37216 23397 37244
rect 23256 37204 23262 37216
rect 23385 37213 23397 37216
rect 23431 37213 23443 37247
rect 23385 37207 23443 37213
rect 23474 37204 23480 37256
rect 23532 37204 23538 37256
rect 23842 37204 23848 37256
rect 23900 37253 23906 37256
rect 23900 37244 23908 37253
rect 24688 37244 24716 37352
rect 26326 37340 26332 37352
rect 26384 37340 26390 37392
rect 27246 37340 27252 37392
rect 27304 37380 27310 37392
rect 28166 37380 28172 37392
rect 27304 37352 28172 37380
rect 27304 37340 27310 37352
rect 28166 37340 28172 37352
rect 28224 37340 28230 37392
rect 25222 37272 25228 37324
rect 25280 37272 25286 37324
rect 27890 37272 27896 37324
rect 27948 37312 27954 37324
rect 28077 37315 28135 37321
rect 28077 37312 28089 37315
rect 27948 37284 28089 37312
rect 27948 37272 27954 37284
rect 28077 37281 28089 37284
rect 28123 37281 28135 37315
rect 28077 37275 28135 37281
rect 28442 37272 28448 37324
rect 28500 37312 28506 37324
rect 28537 37315 28595 37321
rect 28537 37312 28549 37315
rect 28500 37284 28549 37312
rect 28500 37272 28506 37284
rect 28537 37281 28549 37284
rect 28583 37312 28595 37315
rect 29086 37312 29092 37324
rect 28583 37284 29092 37312
rect 28583 37281 28595 37284
rect 28537 37275 28595 37281
rect 29086 37272 29092 37284
rect 29144 37272 29150 37324
rect 23900 37216 24716 37244
rect 23900 37207 23908 37216
rect 23900 37204 23906 37207
rect 24854 37204 24860 37256
rect 24912 37204 24918 37256
rect 25409 37247 25467 37253
rect 25409 37213 25421 37247
rect 25455 37244 25467 37247
rect 26050 37244 26056 37256
rect 25455 37216 26056 37244
rect 25455 37213 25467 37216
rect 25409 37207 25467 37213
rect 26050 37204 26056 37216
rect 26108 37204 26114 37256
rect 26418 37204 26424 37256
rect 26476 37204 26482 37256
rect 26605 37247 26663 37253
rect 26605 37213 26617 37247
rect 26651 37244 26663 37247
rect 26786 37244 26792 37256
rect 26651 37216 26792 37244
rect 26651 37213 26663 37216
rect 26605 37207 26663 37213
rect 26786 37204 26792 37216
rect 26844 37204 26850 37256
rect 26973 37247 27031 37253
rect 26973 37213 26985 37247
rect 27019 37213 27031 37247
rect 26973 37207 27031 37213
rect 27157 37247 27215 37253
rect 27157 37213 27169 37247
rect 27203 37244 27215 37247
rect 27246 37244 27252 37256
rect 27203 37216 27252 37244
rect 27203 37213 27215 37216
rect 27157 37207 27215 37213
rect 23566 37136 23572 37188
rect 23624 37176 23630 37188
rect 23661 37179 23719 37185
rect 23661 37176 23673 37179
rect 23624 37148 23673 37176
rect 23624 37136 23630 37148
rect 23661 37145 23673 37148
rect 23707 37145 23719 37179
rect 23661 37139 23719 37145
rect 23753 37179 23811 37185
rect 23753 37145 23765 37179
rect 23799 37176 23811 37179
rect 24118 37176 24124 37188
rect 23799 37148 24124 37176
rect 23799 37145 23811 37148
rect 23753 37139 23811 37145
rect 24118 37136 24124 37148
rect 24176 37136 24182 37188
rect 24946 37136 24952 37188
rect 25004 37176 25010 37188
rect 25041 37179 25099 37185
rect 25041 37176 25053 37179
rect 25004 37148 25053 37176
rect 25004 37136 25010 37148
rect 25041 37145 25053 37148
rect 25087 37145 25099 37179
rect 25041 37139 25099 37145
rect 25774 37136 25780 37188
rect 25832 37176 25838 37188
rect 25961 37179 26019 37185
rect 25961 37176 25973 37179
rect 25832 37148 25973 37176
rect 25832 37136 25838 37148
rect 25961 37145 25973 37148
rect 26007 37145 26019 37179
rect 25961 37139 26019 37145
rect 26988 37176 27016 37207
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 27614 37204 27620 37256
rect 27672 37204 27678 37256
rect 28258 37204 28264 37256
rect 28316 37204 28322 37256
rect 28629 37247 28687 37253
rect 28629 37213 28641 37247
rect 28675 37244 28687 37247
rect 29196 37244 29224 37420
rect 31018 37408 31024 37420
rect 31076 37408 31082 37460
rect 31478 37408 31484 37460
rect 31536 37448 31542 37460
rect 32214 37448 32220 37460
rect 31536 37420 32220 37448
rect 31536 37408 31542 37420
rect 32214 37408 32220 37420
rect 32272 37408 32278 37460
rect 32953 37451 33011 37457
rect 32953 37448 32965 37451
rect 32876 37420 32965 37448
rect 31754 37340 31760 37392
rect 31812 37380 31818 37392
rect 32582 37380 32588 37392
rect 31812 37352 32588 37380
rect 31812 37340 31818 37352
rect 32582 37340 32588 37352
rect 32640 37340 32646 37392
rect 31018 37272 31024 37324
rect 31076 37312 31082 37324
rect 32876 37312 32904 37420
rect 32953 37417 32965 37420
rect 32999 37448 33011 37451
rect 36354 37448 36360 37460
rect 32999 37420 36360 37448
rect 32999 37417 33011 37420
rect 32953 37411 33011 37417
rect 36354 37408 36360 37420
rect 36412 37408 36418 37460
rect 36906 37408 36912 37460
rect 36964 37408 36970 37460
rect 37458 37408 37464 37460
rect 37516 37408 37522 37460
rect 39850 37448 39856 37460
rect 37752 37420 39856 37448
rect 34146 37340 34152 37392
rect 34204 37340 34210 37392
rect 34790 37340 34796 37392
rect 34848 37380 34854 37392
rect 34848 37352 35296 37380
rect 34848 37340 34854 37352
rect 31076 37284 32904 37312
rect 31076 37272 31082 37284
rect 33042 37272 33048 37324
rect 33100 37312 33106 37324
rect 33962 37312 33968 37324
rect 33100 37284 33824 37312
rect 33100 37272 33106 37284
rect 29270 37244 29276 37256
rect 28675 37216 29276 37244
rect 28675 37213 28687 37216
rect 28629 37207 28687 37213
rect 28644 37176 28672 37207
rect 29270 37204 29276 37216
rect 29328 37204 29334 37256
rect 29914 37204 29920 37256
rect 29972 37204 29978 37256
rect 30006 37204 30012 37256
rect 30064 37244 30070 37256
rect 30173 37247 30231 37253
rect 30173 37244 30185 37247
rect 30064 37216 30185 37244
rect 30064 37204 30070 37216
rect 30173 37213 30185 37216
rect 30219 37213 30231 37247
rect 30173 37207 30231 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31895 37247 31953 37253
rect 31895 37244 31907 37247
rect 30984 37216 31907 37244
rect 30984 37204 30990 37216
rect 31895 37213 31907 37216
rect 31941 37213 31953 37247
rect 31895 37207 31953 37213
rect 32030 37204 32036 37256
rect 32088 37204 32094 37256
rect 32253 37247 32311 37253
rect 32253 37244 32265 37247
rect 32232 37213 32265 37244
rect 32299 37213 32311 37247
rect 32232 37207 32311 37213
rect 32401 37247 32459 37253
rect 32401 37213 32413 37247
rect 32447 37244 32459 37247
rect 32582 37244 32588 37256
rect 32447 37216 32588 37244
rect 32447 37213 32459 37216
rect 32401 37207 32459 37213
rect 26988 37148 28672 37176
rect 22428 37080 22600 37108
rect 22428 37068 22434 37080
rect 22646 37068 22652 37120
rect 22704 37108 22710 37120
rect 24670 37108 24676 37120
rect 22704 37080 24676 37108
rect 22704 37068 22710 37080
rect 24670 37068 24676 37080
rect 24728 37108 24734 37120
rect 26988 37108 27016 37148
rect 29362 37136 29368 37188
rect 29420 37176 29426 37188
rect 30282 37176 30288 37188
rect 29420 37148 30288 37176
rect 29420 37136 29426 37148
rect 30282 37136 30288 37148
rect 30340 37136 30346 37188
rect 30374 37136 30380 37188
rect 30432 37176 30438 37188
rect 30432 37148 31984 37176
rect 30432 37136 30438 37148
rect 24728 37080 27016 37108
rect 24728 37068 24734 37080
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 30558 37108 30564 37120
rect 27764 37080 30564 37108
rect 27764 37068 27770 37080
rect 30558 37068 30564 37080
rect 30616 37108 30622 37120
rect 31297 37111 31355 37117
rect 31297 37108 31309 37111
rect 30616 37080 31309 37108
rect 30616 37068 30622 37080
rect 31297 37077 31309 37080
rect 31343 37077 31355 37111
rect 31297 37071 31355 37077
rect 31757 37111 31815 37117
rect 31757 37077 31769 37111
rect 31803 37108 31815 37111
rect 31846 37108 31852 37120
rect 31803 37080 31852 37108
rect 31803 37077 31815 37080
rect 31757 37071 31815 37077
rect 31846 37068 31852 37080
rect 31904 37068 31910 37120
rect 31956 37108 31984 37148
rect 32122 37136 32128 37188
rect 32180 37136 32186 37188
rect 32232 37108 32260 37207
rect 32582 37204 32588 37216
rect 32640 37244 32646 37256
rect 33594 37244 33600 37256
rect 32640 37216 33600 37244
rect 32640 37204 32646 37216
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 33690 37247 33748 37253
rect 33690 37213 33702 37247
rect 33736 37213 33748 37247
rect 33690 37207 33748 37213
rect 33226 37136 33232 37188
rect 33284 37176 33290 37188
rect 33704 37176 33732 37207
rect 33284 37148 33732 37176
rect 33796 37176 33824 37284
rect 33888 37284 33968 37312
rect 33888 37253 33916 37284
rect 33962 37272 33968 37284
rect 34020 37312 34026 37324
rect 34164 37312 34192 37340
rect 34020 37284 35204 37312
rect 34020 37272 34026 37284
rect 35176 37256 35204 37284
rect 34146 37253 34152 37256
rect 33873 37247 33931 37253
rect 33873 37213 33885 37247
rect 33919 37213 33931 37247
rect 33873 37207 33931 37213
rect 34103 37247 34152 37253
rect 34103 37213 34115 37247
rect 34149 37213 34152 37247
rect 34103 37207 34152 37213
rect 34146 37204 34152 37207
rect 34204 37244 34210 37256
rect 34514 37244 34520 37256
rect 34204 37216 34520 37244
rect 34204 37204 34210 37216
rect 34514 37204 34520 37216
rect 34572 37244 34578 37256
rect 34790 37244 34796 37256
rect 34572 37216 34796 37244
rect 34572 37204 34578 37216
rect 34790 37204 34796 37216
rect 34848 37204 34854 37256
rect 35066 37253 35072 37256
rect 34885 37247 34943 37253
rect 34885 37213 34897 37247
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 35033 37247 35072 37253
rect 35033 37213 35045 37247
rect 35033 37207 35072 37213
rect 33965 37179 34023 37185
rect 33965 37176 33977 37179
rect 33796 37148 33977 37176
rect 33284 37136 33290 37148
rect 33965 37145 33977 37148
rect 34011 37145 34023 37179
rect 34422 37176 34428 37188
rect 33965 37139 34023 37145
rect 34169 37148 34428 37176
rect 31956 37080 32260 37108
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 33502 37108 33508 37120
rect 32456 37080 33508 37108
rect 32456 37068 32462 37080
rect 33502 37068 33508 37080
rect 33560 37068 33566 37120
rect 33594 37068 33600 37120
rect 33652 37108 33658 37120
rect 34169 37108 34197 37148
rect 34422 37136 34428 37148
rect 34480 37176 34486 37188
rect 34900 37176 34928 37207
rect 35066 37204 35072 37207
rect 35124 37204 35130 37256
rect 35158 37204 35164 37256
rect 35216 37204 35222 37256
rect 35268 37253 35296 37352
rect 37090 37340 37096 37392
rect 37148 37380 37154 37392
rect 37752 37380 37780 37420
rect 39850 37408 39856 37420
rect 39908 37408 39914 37460
rect 40678 37408 40684 37460
rect 40736 37408 40742 37460
rect 39390 37380 39396 37392
rect 37148 37352 37780 37380
rect 37844 37352 39396 37380
rect 37148 37340 37154 37352
rect 36630 37312 36636 37324
rect 35728 37284 36636 37312
rect 35253 37247 35311 37253
rect 35253 37213 35265 37247
rect 35299 37213 35311 37247
rect 35253 37207 35311 37213
rect 35391 37247 35449 37253
rect 35391 37213 35403 37247
rect 35437 37244 35449 37247
rect 35618 37244 35624 37256
rect 35437 37216 35624 37244
rect 35437 37213 35449 37216
rect 35391 37207 35449 37213
rect 35618 37204 35624 37216
rect 35676 37204 35682 37256
rect 35728 37176 35756 37284
rect 36630 37272 36636 37284
rect 36688 37272 36694 37324
rect 36357 37247 36415 37253
rect 36357 37213 36369 37247
rect 36403 37244 36415 37247
rect 36446 37244 36452 37256
rect 36403 37216 36452 37244
rect 36403 37213 36415 37216
rect 36357 37207 36415 37213
rect 36446 37204 36452 37216
rect 36504 37204 36510 37256
rect 36725 37247 36783 37253
rect 36725 37213 36737 37247
rect 36771 37244 36783 37247
rect 36814 37244 36820 37256
rect 36771 37216 36820 37244
rect 36771 37213 36783 37216
rect 36725 37207 36783 37213
rect 36814 37204 36820 37216
rect 36872 37204 36878 37256
rect 37844 37253 37872 37352
rect 39390 37340 39396 37352
rect 39448 37340 39454 37392
rect 39574 37340 39580 37392
rect 39632 37380 39638 37392
rect 40770 37380 40776 37392
rect 39632 37352 40776 37380
rect 39632 37340 39638 37352
rect 40770 37340 40776 37352
rect 40828 37340 40834 37392
rect 41414 37340 41420 37392
rect 41472 37340 41478 37392
rect 39298 37272 39304 37324
rect 39356 37312 39362 37324
rect 39356 37284 40448 37312
rect 39356 37272 39362 37284
rect 37829 37247 37887 37253
rect 37829 37213 37841 37247
rect 37875 37213 37887 37247
rect 37829 37207 37887 37213
rect 38102 37204 38108 37256
rect 38160 37204 38166 37256
rect 38194 37204 38200 37256
rect 38252 37204 38258 37256
rect 38286 37204 38292 37256
rect 38344 37244 38350 37256
rect 38470 37244 38476 37256
rect 38344 37216 38476 37244
rect 38344 37204 38350 37216
rect 38470 37204 38476 37216
rect 38528 37204 38534 37256
rect 38654 37204 38660 37256
rect 38712 37204 38718 37256
rect 40218 37253 40224 37256
rect 40037 37247 40095 37253
rect 40037 37244 40049 37247
rect 38764 37216 40049 37244
rect 34480 37148 34928 37176
rect 34992 37148 35756 37176
rect 34480 37136 34486 37148
rect 33652 37080 34197 37108
rect 33652 37068 33658 37080
rect 34238 37068 34244 37120
rect 34296 37068 34302 37120
rect 34606 37068 34612 37120
rect 34664 37108 34670 37120
rect 34992 37108 35020 37148
rect 36170 37136 36176 37188
rect 36228 37176 36234 37188
rect 36538 37176 36544 37188
rect 36228 37148 36544 37176
rect 36228 37136 36234 37148
rect 36538 37136 36544 37148
rect 36596 37136 36602 37188
rect 36633 37179 36691 37185
rect 36633 37145 36645 37179
rect 36679 37176 36691 37179
rect 37182 37176 37188 37188
rect 36679 37148 37188 37176
rect 36679 37145 36691 37148
rect 36633 37139 36691 37145
rect 37182 37136 37188 37148
rect 37240 37136 37246 37188
rect 37384 37148 37688 37176
rect 34664 37080 35020 37108
rect 34664 37068 34670 37080
rect 35066 37068 35072 37120
rect 35124 37108 35130 37120
rect 35434 37108 35440 37120
rect 35124 37080 35440 37108
rect 35124 37068 35130 37080
rect 35434 37068 35440 37080
rect 35492 37068 35498 37120
rect 35529 37111 35587 37117
rect 35529 37077 35541 37111
rect 35575 37108 35587 37111
rect 37384 37108 37412 37148
rect 35575 37080 37412 37108
rect 37660 37108 37688 37148
rect 38764 37108 38792 37216
rect 40037 37213 40049 37216
rect 40083 37213 40095 37247
rect 40037 37207 40095 37213
rect 40185 37247 40224 37253
rect 40185 37213 40197 37247
rect 40185 37207 40224 37213
rect 40218 37204 40224 37207
rect 40276 37204 40282 37256
rect 40420 37253 40448 37284
rect 40586 37253 40592 37256
rect 40405 37247 40463 37253
rect 40405 37213 40417 37247
rect 40451 37213 40463 37247
rect 40405 37207 40463 37213
rect 40543 37247 40592 37253
rect 40543 37213 40555 37247
rect 40589 37213 40592 37247
rect 40543 37207 40592 37213
rect 40586 37204 40592 37207
rect 40644 37204 40650 37256
rect 41138 37204 41144 37256
rect 41196 37204 41202 37256
rect 41230 37204 41236 37256
rect 41288 37204 41294 37256
rect 41874 37204 41880 37256
rect 41932 37204 41938 37256
rect 40310 37136 40316 37188
rect 40368 37136 40374 37188
rect 40770 37136 40776 37188
rect 40828 37176 40834 37188
rect 41322 37176 41328 37188
rect 40828 37148 41328 37176
rect 40828 37136 40834 37148
rect 41322 37136 41328 37148
rect 41380 37176 41386 37188
rect 41417 37179 41475 37185
rect 41417 37176 41429 37179
rect 41380 37148 41429 37176
rect 41380 37136 41386 37148
rect 41417 37145 41429 37148
rect 41463 37145 41475 37179
rect 41417 37139 41475 37145
rect 41966 37136 41972 37188
rect 42024 37176 42030 37188
rect 42122 37179 42180 37185
rect 42122 37176 42134 37179
rect 42024 37148 42134 37176
rect 42024 37136 42030 37148
rect 42122 37145 42134 37148
rect 42168 37145 42180 37179
rect 42122 37139 42180 37145
rect 37660 37080 38792 37108
rect 35575 37077 35587 37080
rect 35529 37071 35587 37077
rect 40218 37068 40224 37120
rect 40276 37108 40282 37120
rect 43257 37111 43315 37117
rect 43257 37108 43269 37111
rect 40276 37080 43269 37108
rect 40276 37068 40282 37080
rect 43257 37077 43269 37080
rect 43303 37077 43315 37111
rect 43257 37071 43315 37077
rect 1104 37018 43884 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 43884 37018
rect 1104 36944 43884 36966
rect 14645 36907 14703 36913
rect 14645 36873 14657 36907
rect 14691 36904 14703 36907
rect 16206 36904 16212 36916
rect 14691 36876 16212 36904
rect 14691 36873 14703 36876
rect 14645 36867 14703 36873
rect 16206 36864 16212 36876
rect 16264 36864 16270 36916
rect 16301 36907 16359 36913
rect 16301 36873 16313 36907
rect 16347 36904 16359 36907
rect 18233 36907 18291 36913
rect 18233 36904 18245 36907
rect 16347 36876 18245 36904
rect 16347 36873 16359 36876
rect 16301 36867 16359 36873
rect 18233 36873 18245 36876
rect 18279 36904 18291 36907
rect 22370 36904 22376 36916
rect 18279 36876 22376 36904
rect 18279 36873 18291 36876
rect 18233 36867 18291 36873
rect 22370 36864 22376 36876
rect 22428 36864 22434 36916
rect 22462 36864 22468 36916
rect 22520 36904 22526 36916
rect 22741 36907 22799 36913
rect 22741 36904 22753 36907
rect 22520 36876 22753 36904
rect 22520 36864 22526 36876
rect 22741 36873 22753 36876
rect 22787 36873 22799 36907
rect 22741 36867 22799 36873
rect 23658 36864 23664 36916
rect 23716 36904 23722 36916
rect 23937 36907 23995 36913
rect 23937 36904 23949 36907
rect 23716 36876 23949 36904
rect 23716 36864 23722 36876
rect 23937 36873 23949 36876
rect 23983 36873 23995 36907
rect 23937 36867 23995 36873
rect 25866 36864 25872 36916
rect 25924 36864 25930 36916
rect 26160 36876 26372 36904
rect 15749 36839 15807 36845
rect 15749 36805 15761 36839
rect 15795 36836 15807 36839
rect 16114 36836 16120 36848
rect 15795 36808 16120 36836
rect 15795 36805 15807 36808
rect 15749 36799 15807 36805
rect 16114 36796 16120 36808
rect 16172 36796 16178 36848
rect 17494 36836 17500 36848
rect 16868 36808 17500 36836
rect 16868 36780 16896 36808
rect 17494 36796 17500 36808
rect 17552 36836 17558 36848
rect 20714 36836 20720 36848
rect 17552 36808 20720 36836
rect 17552 36796 17558 36808
rect 16850 36728 16856 36780
rect 16908 36728 16914 36780
rect 18800 36777 18828 36808
rect 20714 36796 20720 36808
rect 20772 36796 20778 36848
rect 23106 36796 23112 36848
rect 23164 36836 23170 36848
rect 24213 36839 24271 36845
rect 24213 36836 24225 36839
rect 23164 36808 24225 36836
rect 23164 36796 23170 36808
rect 24213 36805 24225 36808
rect 24259 36836 24271 36839
rect 24394 36836 24400 36848
rect 24259 36808 24400 36836
rect 24259 36805 24271 36808
rect 24213 36799 24271 36805
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 24762 36836 24768 36848
rect 24504 36808 24768 36836
rect 17109 36771 17167 36777
rect 17109 36768 17121 36771
rect 16960 36740 17121 36768
rect 16206 36660 16212 36712
rect 16264 36700 16270 36712
rect 16960 36700 16988 36740
rect 17109 36737 17121 36740
rect 17155 36737 17167 36771
rect 17109 36731 17167 36737
rect 18785 36771 18843 36777
rect 18785 36737 18797 36771
rect 18831 36737 18843 36771
rect 18785 36731 18843 36737
rect 19052 36771 19110 36777
rect 19052 36737 19064 36771
rect 19098 36768 19110 36771
rect 19426 36768 19432 36780
rect 19098 36740 19432 36768
rect 19098 36737 19110 36740
rect 19052 36731 19110 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 20254 36728 20260 36780
rect 20312 36768 20318 36780
rect 22465 36771 22523 36777
rect 20312 36740 22232 36768
rect 20312 36728 20318 36740
rect 22204 36709 22232 36740
rect 22465 36737 22477 36771
rect 22511 36768 22523 36771
rect 22646 36768 22652 36780
rect 22511 36740 22652 36768
rect 22511 36737 22523 36740
rect 22465 36731 22523 36737
rect 22646 36728 22652 36740
rect 22704 36728 22710 36780
rect 24118 36777 24124 36780
rect 24116 36731 24124 36777
rect 24118 36728 24124 36731
rect 24176 36728 24182 36780
rect 24302 36728 24308 36780
rect 24360 36728 24366 36780
rect 24504 36777 24532 36808
rect 24762 36796 24768 36808
rect 24820 36796 24826 36848
rect 25884 36836 25912 36864
rect 26160 36845 26188 36876
rect 26053 36839 26111 36845
rect 26053 36836 26065 36839
rect 25884 36808 26065 36836
rect 26053 36805 26065 36808
rect 26099 36805 26111 36839
rect 26053 36799 26111 36805
rect 26145 36839 26203 36845
rect 26145 36805 26157 36839
rect 26191 36805 26203 36839
rect 26344 36836 26372 36876
rect 26418 36864 26424 36916
rect 26476 36864 26482 36916
rect 27338 36864 27344 36916
rect 27396 36864 27402 36916
rect 28534 36864 28540 36916
rect 28592 36864 28598 36916
rect 30466 36864 30472 36916
rect 30524 36864 30530 36916
rect 30558 36864 30564 36916
rect 30616 36904 30622 36916
rect 32122 36904 32128 36916
rect 30616 36876 32128 36904
rect 30616 36864 30622 36876
rect 32122 36864 32128 36876
rect 32180 36864 32186 36916
rect 32858 36864 32864 36916
rect 32916 36904 32922 36916
rect 33045 36907 33103 36913
rect 33045 36904 33057 36907
rect 32916 36876 33057 36904
rect 32916 36864 32922 36876
rect 33045 36873 33057 36876
rect 33091 36873 33103 36907
rect 33045 36867 33103 36873
rect 33226 36864 33232 36916
rect 33284 36904 33290 36916
rect 33778 36904 33784 36916
rect 33284 36876 33784 36904
rect 33284 36864 33290 36876
rect 33778 36864 33784 36876
rect 33836 36864 33842 36916
rect 33888 36876 34376 36904
rect 26694 36836 26700 36848
rect 26344 36808 26700 36836
rect 26145 36799 26203 36805
rect 26694 36796 26700 36808
rect 26752 36796 26758 36848
rect 27356 36836 27384 36864
rect 26804 36808 27384 36836
rect 27433 36839 27491 36845
rect 24488 36771 24546 36777
rect 24488 36737 24500 36771
rect 24534 36737 24546 36771
rect 24488 36731 24546 36737
rect 24581 36771 24639 36777
rect 24581 36737 24593 36771
rect 24627 36768 24639 36771
rect 24670 36768 24676 36780
rect 24627 36740 24676 36768
rect 24627 36737 24639 36740
rect 24581 36731 24639 36737
rect 24670 36728 24676 36740
rect 24728 36728 24734 36780
rect 25038 36728 25044 36780
rect 25096 36728 25102 36780
rect 25225 36771 25283 36777
rect 25225 36737 25237 36771
rect 25271 36768 25283 36771
rect 25406 36768 25412 36780
rect 25271 36740 25412 36768
rect 25271 36737 25283 36740
rect 25225 36731 25283 36737
rect 25406 36728 25412 36740
rect 25464 36728 25470 36780
rect 25774 36728 25780 36780
rect 25832 36728 25838 36780
rect 25866 36728 25872 36780
rect 25924 36768 25930 36780
rect 26326 36777 26332 36780
rect 26283 36771 26332 36777
rect 25924 36740 25969 36768
rect 25924 36728 25930 36740
rect 26283 36737 26295 36771
rect 26329 36737 26332 36771
rect 26283 36731 26332 36737
rect 26326 36728 26332 36731
rect 26384 36768 26390 36780
rect 26804 36768 26832 36808
rect 27433 36805 27445 36839
rect 27479 36836 27491 36839
rect 33888 36836 33916 36876
rect 34348 36848 34376 36876
rect 35342 36864 35348 36916
rect 35400 36904 35406 36916
rect 35621 36907 35679 36913
rect 35621 36904 35633 36907
rect 35400 36876 35633 36904
rect 35400 36864 35406 36876
rect 35621 36873 35633 36876
rect 35667 36873 35679 36907
rect 35621 36867 35679 36873
rect 36909 36907 36967 36913
rect 36909 36873 36921 36907
rect 36955 36904 36967 36907
rect 38194 36904 38200 36916
rect 36955 36876 38200 36904
rect 36955 36873 36967 36876
rect 36909 36867 36967 36873
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 39114 36864 39120 36916
rect 39172 36904 39178 36916
rect 39172 36876 40724 36904
rect 39172 36864 39178 36876
rect 27479 36808 33916 36836
rect 27479 36805 27491 36808
rect 27433 36799 27491 36805
rect 33962 36796 33968 36848
rect 34020 36796 34026 36848
rect 34330 36796 34336 36848
rect 34388 36836 34394 36848
rect 35253 36839 35311 36845
rect 34388 36808 35112 36836
rect 34388 36796 34394 36808
rect 26384 36740 26832 36768
rect 27341 36771 27399 36777
rect 26384 36728 26390 36740
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 16264 36672 16988 36700
rect 21453 36703 21511 36709
rect 16264 36660 16270 36672
rect 21453 36669 21465 36703
rect 21499 36700 21511 36703
rect 22097 36703 22155 36709
rect 21499 36672 21588 36700
rect 21499 36669 21511 36672
rect 21453 36663 21511 36669
rect 21560 36644 21588 36672
rect 22097 36669 22109 36703
rect 22143 36669 22155 36703
rect 22097 36663 22155 36669
rect 22189 36703 22247 36709
rect 22189 36669 22201 36703
rect 22235 36700 22247 36703
rect 22278 36700 22284 36712
rect 22235 36672 22284 36700
rect 22235 36669 22247 36672
rect 22189 36663 22247 36669
rect 14090 36592 14096 36644
rect 14148 36592 14154 36644
rect 15197 36635 15255 36641
rect 15197 36601 15209 36635
rect 15243 36632 15255 36635
rect 20901 36635 20959 36641
rect 15243 36604 16896 36632
rect 15243 36601 15255 36604
rect 15197 36595 15255 36601
rect 16868 36564 16896 36604
rect 20901 36601 20913 36635
rect 20947 36632 20959 36635
rect 20947 36604 21496 36632
rect 20947 36601 20959 36604
rect 20901 36595 20959 36601
rect 19978 36564 19984 36576
rect 16868 36536 19984 36564
rect 19978 36524 19984 36536
rect 20036 36524 20042 36576
rect 20162 36524 20168 36576
rect 20220 36524 20226 36576
rect 21468 36564 21496 36604
rect 21542 36592 21548 36644
rect 21600 36632 21606 36644
rect 22112 36632 22140 36663
rect 22278 36660 22284 36672
rect 22336 36660 22342 36712
rect 22554 36660 22560 36712
rect 22612 36660 22618 36712
rect 23382 36700 23388 36712
rect 22664 36672 23388 36700
rect 22664 36632 22692 36672
rect 23382 36660 23388 36672
rect 23440 36660 23446 36712
rect 25792 36700 25820 36728
rect 26142 36700 26148 36712
rect 25792 36672 26148 36700
rect 26142 36660 26148 36672
rect 26200 36660 26206 36712
rect 26510 36660 26516 36712
rect 26568 36700 26574 36712
rect 27062 36700 27068 36712
rect 26568 36672 27068 36700
rect 26568 36660 26574 36672
rect 27062 36660 27068 36672
rect 27120 36660 27126 36712
rect 27356 36700 27384 36731
rect 27522 36728 27528 36780
rect 27580 36728 27586 36780
rect 27709 36771 27767 36777
rect 27709 36737 27721 36771
rect 27755 36768 27767 36771
rect 28074 36768 28080 36780
rect 27755 36740 28080 36768
rect 27755 36737 27767 36740
rect 27709 36731 27767 36737
rect 28074 36728 28080 36740
rect 28132 36728 28138 36780
rect 28905 36771 28963 36777
rect 28905 36737 28917 36771
rect 28951 36768 28963 36771
rect 29086 36768 29092 36780
rect 28951 36740 29092 36768
rect 28951 36737 28963 36740
rect 28905 36731 28963 36737
rect 29086 36728 29092 36740
rect 29144 36728 29150 36780
rect 29270 36728 29276 36780
rect 29328 36728 29334 36780
rect 29454 36728 29460 36780
rect 29512 36728 29518 36780
rect 29917 36771 29975 36777
rect 29917 36737 29929 36771
rect 29963 36737 29975 36771
rect 29917 36731 29975 36737
rect 27430 36700 27436 36712
rect 27356 36672 27436 36700
rect 27430 36660 27436 36672
rect 27488 36660 27494 36712
rect 28813 36703 28871 36709
rect 28813 36669 28825 36703
rect 28859 36700 28871 36703
rect 28994 36700 29000 36712
rect 28859 36672 29000 36700
rect 28859 36669 28871 36672
rect 28813 36663 28871 36669
rect 28994 36660 29000 36672
rect 29052 36660 29058 36712
rect 29932 36700 29960 36731
rect 30098 36728 30104 36780
rect 30156 36728 30162 36780
rect 30190 36728 30196 36780
rect 30248 36728 30254 36780
rect 30282 36728 30288 36780
rect 30340 36728 30346 36780
rect 30926 36728 30932 36780
rect 30984 36768 30990 36780
rect 31202 36768 31208 36780
rect 30984 36740 31208 36768
rect 30984 36728 30990 36740
rect 31202 36728 31208 36740
rect 31260 36728 31266 36780
rect 31570 36728 31576 36780
rect 31628 36768 31634 36780
rect 32490 36768 32496 36780
rect 31628 36740 32496 36768
rect 31628 36728 31634 36740
rect 32490 36728 32496 36740
rect 32548 36728 32554 36780
rect 32674 36728 32680 36780
rect 32732 36728 32738 36780
rect 32766 36728 32772 36780
rect 32824 36728 32830 36780
rect 32861 36771 32919 36777
rect 32861 36737 32873 36771
rect 32907 36768 32919 36771
rect 33502 36768 33508 36780
rect 32907 36740 33508 36768
rect 32907 36737 32919 36740
rect 32861 36731 32919 36737
rect 33502 36728 33508 36740
rect 33560 36728 33566 36780
rect 33594 36728 33600 36780
rect 33652 36768 33658 36780
rect 33689 36771 33747 36777
rect 33689 36768 33701 36771
rect 33652 36740 33701 36768
rect 33652 36728 33658 36740
rect 33689 36737 33701 36740
rect 33735 36737 33747 36771
rect 33689 36731 33747 36737
rect 33782 36771 33840 36777
rect 33782 36737 33794 36771
rect 33828 36737 33840 36771
rect 33782 36731 33840 36737
rect 29380 36672 29960 36700
rect 30116 36700 30144 36728
rect 30558 36700 30564 36712
rect 30116 36672 30564 36700
rect 21600 36604 22692 36632
rect 21600 36592 21606 36604
rect 22830 36592 22836 36644
rect 22888 36632 22894 36644
rect 29380 36632 29408 36672
rect 30558 36660 30564 36672
rect 30616 36660 30622 36712
rect 32306 36660 32312 36712
rect 32364 36700 32370 36712
rect 33134 36700 33140 36712
rect 32364 36672 33140 36700
rect 32364 36660 32370 36672
rect 33134 36660 33140 36672
rect 33192 36700 33198 36712
rect 33796 36700 33824 36731
rect 33870 36728 33876 36780
rect 33928 36768 33934 36780
rect 34057 36771 34115 36777
rect 34057 36768 34069 36771
rect 33928 36740 34069 36768
rect 33928 36728 33934 36740
rect 34057 36737 34069 36740
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 34146 36728 34152 36780
rect 34204 36777 34210 36780
rect 35084 36777 35112 36808
rect 35253 36805 35265 36839
rect 35299 36836 35311 36839
rect 35802 36836 35808 36848
rect 35299 36808 35808 36836
rect 35299 36805 35311 36808
rect 35253 36799 35311 36805
rect 35802 36796 35808 36808
rect 35860 36796 35866 36848
rect 36170 36796 36176 36848
rect 36228 36836 36234 36848
rect 36541 36839 36599 36845
rect 36541 36836 36553 36839
rect 36228 36808 36553 36836
rect 36228 36796 36234 36808
rect 36541 36805 36553 36808
rect 36587 36805 36599 36839
rect 36541 36799 36599 36805
rect 38286 36796 38292 36848
rect 38344 36836 38350 36848
rect 38344 36808 38608 36836
rect 38344 36796 38350 36808
rect 34204 36768 34212 36777
rect 34977 36771 35035 36777
rect 34977 36768 34989 36771
rect 34204 36740 34249 36768
rect 34348 36740 34989 36768
rect 34204 36731 34212 36740
rect 34204 36728 34210 36731
rect 33192 36672 33824 36700
rect 33192 36660 33198 36672
rect 22888 36604 29408 36632
rect 22888 36592 22894 36604
rect 33594 36592 33600 36644
rect 33652 36632 33658 36644
rect 34146 36632 34152 36644
rect 33652 36604 34152 36632
rect 33652 36592 33658 36604
rect 34146 36592 34152 36604
rect 34204 36592 34210 36644
rect 34348 36641 34376 36740
rect 34977 36737 34989 36740
rect 35023 36737 35035 36771
rect 34977 36731 35035 36737
rect 35070 36771 35128 36777
rect 35070 36737 35082 36771
rect 35116 36737 35128 36771
rect 35070 36731 35128 36737
rect 35158 36728 35164 36780
rect 35216 36768 35222 36780
rect 35345 36771 35403 36777
rect 35345 36768 35357 36771
rect 35216 36740 35357 36768
rect 35216 36728 35222 36740
rect 35345 36737 35357 36740
rect 35391 36737 35403 36771
rect 35345 36731 35403 36737
rect 35483 36771 35541 36777
rect 35483 36737 35495 36771
rect 35529 36768 35541 36771
rect 35894 36768 35900 36780
rect 35529 36740 35900 36768
rect 35529 36737 35541 36740
rect 35483 36731 35541 36737
rect 35894 36728 35900 36740
rect 35952 36728 35958 36780
rect 36354 36728 36360 36780
rect 36412 36728 36418 36780
rect 36630 36728 36636 36780
rect 36688 36728 36694 36780
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 36814 36768 36820 36780
rect 36771 36740 36820 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 36814 36728 36820 36740
rect 36872 36728 36878 36780
rect 37642 36728 37648 36780
rect 37700 36768 37706 36780
rect 38378 36768 38384 36780
rect 37700 36740 38384 36768
rect 37700 36728 37706 36740
rect 38378 36728 38384 36740
rect 38436 36728 38442 36780
rect 38580 36777 38608 36808
rect 39666 36796 39672 36848
rect 39724 36796 39730 36848
rect 39942 36796 39948 36848
rect 40000 36836 40006 36848
rect 40497 36839 40555 36845
rect 40497 36836 40509 36839
rect 40000 36808 40509 36836
rect 40000 36796 40006 36808
rect 40497 36805 40509 36808
rect 40543 36805 40555 36839
rect 40696 36836 40724 36876
rect 40770 36864 40776 36916
rect 40828 36864 40834 36916
rect 41414 36864 41420 36916
rect 41472 36864 41478 36916
rect 41966 36864 41972 36916
rect 42024 36864 42030 36916
rect 41432 36836 41460 36864
rect 40696 36808 40816 36836
rect 41432 36808 42104 36836
rect 40497 36799 40555 36805
rect 38565 36771 38623 36777
rect 38565 36737 38577 36771
rect 38611 36737 38623 36771
rect 38565 36731 38623 36737
rect 38841 36771 38899 36777
rect 38841 36737 38853 36771
rect 38887 36737 38899 36771
rect 38841 36731 38899 36737
rect 39117 36771 39175 36777
rect 39117 36737 39129 36771
rect 39163 36737 39175 36771
rect 39117 36731 39175 36737
rect 39209 36771 39267 36777
rect 39209 36737 39221 36771
rect 39255 36768 39267 36771
rect 39390 36768 39396 36780
rect 39255 36740 39396 36768
rect 39255 36737 39267 36740
rect 39209 36731 39267 36737
rect 34333 36635 34391 36641
rect 34333 36601 34345 36635
rect 34379 36601 34391 36635
rect 34333 36595 34391 36601
rect 35894 36592 35900 36644
rect 35952 36632 35958 36644
rect 36998 36632 37004 36644
rect 35952 36604 37004 36632
rect 35952 36592 35958 36604
rect 36998 36592 37004 36604
rect 37056 36592 37062 36644
rect 37553 36635 37611 36641
rect 37553 36601 37565 36635
rect 37599 36632 37611 36635
rect 37918 36632 37924 36644
rect 37599 36604 37924 36632
rect 37599 36601 37611 36604
rect 37553 36595 37611 36601
rect 37918 36592 37924 36604
rect 37976 36592 37982 36644
rect 38010 36592 38016 36644
rect 38068 36632 38074 36644
rect 38654 36632 38660 36644
rect 38068 36604 38660 36632
rect 38068 36592 38074 36604
rect 38654 36592 38660 36604
rect 38712 36592 38718 36644
rect 38856 36632 38884 36731
rect 39132 36700 39160 36731
rect 39390 36728 39396 36740
rect 39448 36728 39454 36780
rect 40126 36728 40132 36780
rect 40184 36728 40190 36780
rect 40218 36728 40224 36780
rect 40276 36728 40282 36780
rect 40310 36728 40316 36780
rect 40368 36768 40374 36780
rect 40405 36771 40463 36777
rect 40405 36768 40417 36771
rect 40368 36740 40417 36768
rect 40368 36728 40374 36740
rect 40405 36737 40417 36740
rect 40451 36737 40463 36771
rect 40405 36731 40463 36737
rect 40586 36728 40592 36780
rect 40644 36777 40650 36780
rect 40644 36768 40652 36777
rect 40644 36740 40689 36768
rect 40644 36731 40652 36740
rect 40644 36728 40650 36731
rect 39482 36700 39488 36712
rect 39132 36672 39488 36700
rect 39482 36660 39488 36672
rect 39540 36660 39546 36712
rect 40236 36700 40264 36728
rect 40144 36672 40264 36700
rect 38930 36632 38936 36644
rect 38856 36604 38936 36632
rect 38930 36592 38936 36604
rect 38988 36592 38994 36644
rect 22370 36564 22376 36576
rect 21468 36536 22376 36564
rect 22370 36524 22376 36536
rect 22428 36564 22434 36576
rect 23198 36564 23204 36576
rect 22428 36536 23204 36564
rect 22428 36524 22434 36536
rect 23198 36524 23204 36536
rect 23256 36524 23262 36576
rect 23382 36524 23388 36576
rect 23440 36564 23446 36576
rect 23477 36567 23535 36573
rect 23477 36564 23489 36567
rect 23440 36536 23489 36564
rect 23440 36524 23446 36536
rect 23477 36533 23489 36536
rect 23523 36564 23535 36567
rect 23658 36564 23664 36576
rect 23523 36536 23664 36564
rect 23523 36533 23535 36536
rect 23477 36527 23535 36533
rect 23658 36524 23664 36536
rect 23716 36524 23722 36576
rect 25130 36524 25136 36576
rect 25188 36524 25194 36576
rect 26326 36524 26332 36576
rect 26384 36564 26390 36576
rect 27157 36567 27215 36573
rect 27157 36564 27169 36567
rect 26384 36536 27169 36564
rect 26384 36524 26390 36536
rect 27157 36533 27169 36536
rect 27203 36533 27215 36567
rect 27157 36527 27215 36533
rect 27614 36524 27620 36576
rect 27672 36564 27678 36576
rect 30374 36564 30380 36576
rect 27672 36536 30380 36564
rect 27672 36524 27678 36536
rect 30374 36524 30380 36536
rect 30432 36524 30438 36576
rect 31021 36567 31079 36573
rect 31021 36533 31033 36567
rect 31067 36564 31079 36567
rect 31202 36564 31208 36576
rect 31067 36536 31208 36564
rect 31067 36533 31079 36536
rect 31021 36527 31079 36533
rect 31202 36524 31208 36536
rect 31260 36524 31266 36576
rect 31573 36567 31631 36573
rect 31573 36533 31585 36567
rect 31619 36564 31631 36567
rect 33686 36564 33692 36576
rect 31619 36536 33692 36564
rect 31619 36533 31631 36536
rect 31573 36527 31631 36533
rect 33686 36524 33692 36536
rect 33744 36564 33750 36576
rect 33870 36564 33876 36576
rect 33744 36536 33876 36564
rect 33744 36524 33750 36536
rect 33870 36524 33876 36536
rect 33928 36524 33934 36576
rect 36354 36524 36360 36576
rect 36412 36564 36418 36576
rect 37734 36564 37740 36576
rect 36412 36536 37740 36564
rect 36412 36524 36418 36536
rect 37734 36524 37740 36536
rect 37792 36524 37798 36576
rect 38102 36524 38108 36576
rect 38160 36564 38166 36576
rect 40144 36564 40172 36672
rect 40788 36632 40816 36808
rect 41230 36728 41236 36780
rect 41288 36728 41294 36780
rect 41417 36771 41475 36777
rect 41417 36737 41429 36771
rect 41463 36768 41475 36771
rect 41506 36768 41512 36780
rect 41463 36740 41512 36768
rect 41463 36737 41475 36740
rect 41417 36731 41475 36737
rect 41506 36728 41512 36740
rect 41564 36768 41570 36780
rect 42076 36777 42104 36808
rect 41877 36771 41935 36777
rect 41877 36768 41889 36771
rect 41564 36740 41889 36768
rect 41564 36728 41570 36740
rect 41877 36737 41889 36740
rect 41923 36737 41935 36771
rect 41877 36731 41935 36737
rect 42061 36771 42119 36777
rect 42061 36737 42073 36771
rect 42107 36737 42119 36771
rect 42061 36731 42119 36737
rect 43346 36728 43352 36780
rect 43404 36768 43410 36780
rect 43990 36768 43996 36780
rect 43404 36740 43996 36768
rect 43404 36728 43410 36740
rect 43990 36728 43996 36740
rect 44048 36728 44054 36780
rect 41046 36660 41052 36712
rect 41104 36700 41110 36712
rect 42518 36700 42524 36712
rect 41104 36672 42524 36700
rect 41104 36660 41110 36672
rect 42518 36660 42524 36672
rect 42576 36660 42582 36712
rect 41782 36632 41788 36644
rect 40788 36604 41788 36632
rect 41782 36592 41788 36604
rect 41840 36592 41846 36644
rect 38160 36536 40172 36564
rect 38160 36524 38166 36536
rect 41322 36524 41328 36576
rect 41380 36524 41386 36576
rect 42242 36524 42248 36576
rect 42300 36564 42306 36576
rect 42613 36567 42671 36573
rect 42613 36564 42625 36567
rect 42300 36536 42625 36564
rect 42300 36524 42306 36536
rect 42613 36533 42625 36536
rect 42659 36533 42671 36567
rect 42613 36527 42671 36533
rect 42978 36524 42984 36576
rect 43036 36564 43042 36576
rect 43165 36567 43223 36573
rect 43165 36564 43177 36567
rect 43036 36536 43177 36564
rect 43036 36524 43042 36536
rect 43165 36533 43177 36536
rect 43211 36533 43223 36567
rect 43165 36527 43223 36533
rect 1104 36474 43884 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 43884 36474
rect 1104 36400 43884 36422
rect 9674 36320 9680 36372
rect 9732 36320 9738 36372
rect 17770 36320 17776 36372
rect 17828 36320 17834 36372
rect 19334 36320 19340 36372
rect 19392 36360 19398 36372
rect 19429 36363 19487 36369
rect 19429 36360 19441 36363
rect 19392 36332 19441 36360
rect 19392 36320 19398 36332
rect 19429 36329 19441 36332
rect 19475 36329 19487 36363
rect 19429 36323 19487 36329
rect 21361 36363 21419 36369
rect 21361 36329 21373 36363
rect 21407 36360 21419 36363
rect 21542 36360 21548 36372
rect 21407 36332 21548 36360
rect 21407 36329 21419 36332
rect 21361 36323 21419 36329
rect 21542 36320 21548 36332
rect 21600 36320 21606 36372
rect 22922 36320 22928 36372
rect 22980 36360 22986 36372
rect 24946 36360 24952 36372
rect 22980 36332 24952 36360
rect 22980 36320 22986 36332
rect 24946 36320 24952 36332
rect 25004 36360 25010 36372
rect 26602 36360 26608 36372
rect 25004 36332 26608 36360
rect 25004 36320 25010 36332
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 26786 36320 26792 36372
rect 26844 36360 26850 36372
rect 28902 36360 28908 36372
rect 26844 36332 28908 36360
rect 26844 36320 26850 36332
rect 28902 36320 28908 36332
rect 28960 36320 28966 36372
rect 30466 36320 30472 36372
rect 30524 36360 30530 36372
rect 30834 36360 30840 36372
rect 30524 36332 30840 36360
rect 30524 36320 30530 36332
rect 30834 36320 30840 36332
rect 30892 36320 30898 36372
rect 31297 36363 31355 36369
rect 31297 36329 31309 36363
rect 31343 36360 31355 36363
rect 31386 36360 31392 36372
rect 31343 36332 31392 36360
rect 31343 36329 31355 36332
rect 31297 36323 31355 36329
rect 31386 36320 31392 36332
rect 31444 36320 31450 36372
rect 32674 36320 32680 36372
rect 32732 36320 32738 36372
rect 33686 36320 33692 36372
rect 33744 36320 33750 36372
rect 33870 36360 33876 36372
rect 33796 36332 33876 36360
rect 21913 36295 21971 36301
rect 21913 36292 21925 36295
rect 19904 36264 21925 36292
rect 16209 36227 16267 36233
rect 16209 36193 16221 36227
rect 16255 36224 16267 36227
rect 16850 36224 16856 36236
rect 16255 36196 16856 36224
rect 16255 36193 16267 36196
rect 16209 36187 16267 36193
rect 9861 36159 9919 36165
rect 9861 36125 9873 36159
rect 9907 36156 9919 36159
rect 14277 36159 14335 36165
rect 9907 36128 10456 36156
rect 9907 36125 9919 36128
rect 9861 36119 9919 36125
rect 10428 36032 10456 36128
rect 14277 36125 14289 36159
rect 14323 36156 14335 36159
rect 16224 36156 16252 36187
rect 16850 36184 16856 36196
rect 16908 36184 16914 36236
rect 19150 36184 19156 36236
rect 19208 36224 19214 36236
rect 19904 36233 19932 36264
rect 21913 36261 21925 36264
rect 21959 36261 21971 36295
rect 21913 36255 21971 36261
rect 23477 36295 23535 36301
rect 23477 36261 23489 36295
rect 23523 36261 23535 36295
rect 23477 36255 23535 36261
rect 19889 36227 19947 36233
rect 19889 36224 19901 36227
rect 19208 36196 19901 36224
rect 19208 36184 19214 36196
rect 19889 36193 19901 36196
rect 19935 36193 19947 36227
rect 19889 36187 19947 36193
rect 20070 36184 20076 36236
rect 20128 36184 20134 36236
rect 22557 36227 22615 36233
rect 22557 36193 22569 36227
rect 22603 36224 22615 36227
rect 23492 36224 23520 36255
rect 23566 36252 23572 36304
rect 23624 36292 23630 36304
rect 23624 36264 23980 36292
rect 23624 36252 23630 36264
rect 23842 36224 23848 36236
rect 22603 36196 23520 36224
rect 23584 36196 23848 36224
rect 22603 36193 22615 36196
rect 22557 36187 22615 36193
rect 14323 36128 16252 36156
rect 14323 36125 14335 36128
rect 14277 36119 14335 36125
rect 16482 36116 16488 36168
rect 16540 36116 16546 36168
rect 19797 36159 19855 36165
rect 19797 36125 19809 36159
rect 19843 36156 19855 36159
rect 20162 36156 20168 36168
rect 19843 36128 20168 36156
rect 19843 36125 19855 36128
rect 19797 36119 19855 36125
rect 20162 36116 20168 36128
rect 20220 36156 20226 36168
rect 20220 36128 22094 36156
rect 20220 36116 20226 36128
rect 12618 36048 12624 36100
rect 12676 36088 12682 36100
rect 14522 36091 14580 36097
rect 14522 36088 14534 36091
rect 12676 36060 14534 36088
rect 12676 36048 12682 36060
rect 14522 36057 14534 36060
rect 14568 36057 14580 36091
rect 20070 36088 20076 36100
rect 14522 36051 14580 36057
rect 18708 36060 20076 36088
rect 10410 35980 10416 36032
rect 10468 35980 10474 36032
rect 15657 36023 15715 36029
rect 15657 35989 15669 36023
rect 15703 36020 15715 36023
rect 17126 36020 17132 36032
rect 15703 35992 17132 36020
rect 15703 35989 15715 35992
rect 15657 35983 15715 35989
rect 17126 35980 17132 35992
rect 17184 36020 17190 36032
rect 18708 36020 18736 36060
rect 20070 36048 20076 36060
rect 20128 36048 20134 36100
rect 22066 36088 22094 36128
rect 22462 36116 22468 36168
rect 22520 36116 22526 36168
rect 22830 36116 22836 36168
rect 22888 36116 22894 36168
rect 22922 36116 22928 36168
rect 22980 36156 22986 36168
rect 23017 36159 23075 36165
rect 23017 36156 23029 36159
rect 22980 36128 23029 36156
rect 22980 36116 22986 36128
rect 23017 36125 23029 36128
rect 23063 36156 23075 36159
rect 23584 36156 23612 36196
rect 23842 36184 23848 36196
rect 23900 36184 23906 36236
rect 23063 36128 23612 36156
rect 23063 36125 23075 36128
rect 23017 36119 23075 36125
rect 23658 36116 23664 36168
rect 23716 36116 23722 36168
rect 22848 36088 22876 36116
rect 23753 36091 23811 36097
rect 23753 36088 23765 36091
rect 22066 36060 22876 36088
rect 23216 36060 23765 36088
rect 17184 35992 18736 36020
rect 17184 35980 17190 35992
rect 18782 35980 18788 36032
rect 18840 35980 18846 36032
rect 20809 36023 20867 36029
rect 20809 35989 20821 36023
rect 20855 36020 20867 36023
rect 23216 36020 23244 36060
rect 23753 36057 23765 36060
rect 23799 36057 23811 36091
rect 23753 36051 23811 36057
rect 23845 36091 23903 36097
rect 23845 36057 23857 36091
rect 23891 36088 23903 36091
rect 23952 36088 23980 36264
rect 24026 36252 24032 36304
rect 24084 36292 24090 36304
rect 24486 36292 24492 36304
rect 24084 36264 24492 36292
rect 24084 36252 24090 36264
rect 24486 36252 24492 36264
rect 24544 36252 24550 36304
rect 26050 36252 26056 36304
rect 26108 36252 26114 36304
rect 28445 36295 28503 36301
rect 28445 36261 28457 36295
rect 28491 36292 28503 36295
rect 29270 36292 29276 36304
rect 28491 36264 29276 36292
rect 28491 36261 28503 36264
rect 28445 36255 28503 36261
rect 29270 36252 29276 36264
rect 29328 36252 29334 36304
rect 31389 36227 31447 36233
rect 31389 36224 31401 36227
rect 26436 36196 30052 36224
rect 26436 36168 26464 36196
rect 24029 36159 24087 36165
rect 24029 36125 24041 36159
rect 24075 36156 24087 36159
rect 24578 36156 24584 36168
rect 24075 36128 24584 36156
rect 24075 36125 24087 36128
rect 24029 36119 24087 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25225 36159 25283 36165
rect 25225 36153 25237 36159
rect 25216 36125 25237 36153
rect 25271 36125 25283 36159
rect 25216 36119 25283 36125
rect 23891 36060 23980 36088
rect 23891 36057 23903 36060
rect 23845 36051 23903 36057
rect 20855 35992 23244 36020
rect 23768 36020 23796 36051
rect 23934 36020 23940 36032
rect 23768 35992 23940 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 23934 35980 23940 35992
rect 23992 35980 23998 36032
rect 24762 35980 24768 36032
rect 24820 36020 24826 36032
rect 25041 36023 25099 36029
rect 25041 36020 25053 36023
rect 24820 35992 25053 36020
rect 24820 35980 24826 35992
rect 25041 35989 25053 35992
rect 25087 35989 25099 36023
rect 25216 36020 25244 36119
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 25593 36159 25651 36165
rect 25593 36156 25605 36159
rect 25556 36128 25605 36156
rect 25556 36116 25562 36128
rect 25593 36125 25605 36128
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 26234 36116 26240 36168
rect 26292 36116 26298 36168
rect 26418 36116 26424 36168
rect 26476 36116 26482 36168
rect 26602 36116 26608 36168
rect 26660 36116 26666 36168
rect 26694 36116 26700 36168
rect 26752 36156 26758 36168
rect 27062 36156 27068 36168
rect 26752 36128 27068 36156
rect 26752 36116 26758 36128
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27249 36159 27307 36165
rect 27249 36125 27261 36159
rect 27295 36125 27307 36159
rect 27249 36119 27307 36125
rect 27617 36159 27675 36165
rect 27617 36125 27629 36159
rect 27663 36156 27675 36159
rect 27798 36156 27804 36168
rect 27663 36128 27804 36156
rect 27663 36125 27675 36128
rect 27617 36119 27675 36125
rect 25314 36048 25320 36100
rect 25372 36048 25378 36100
rect 25409 36091 25467 36097
rect 25409 36057 25421 36091
rect 25455 36088 25467 36091
rect 26050 36088 26056 36100
rect 25455 36060 26056 36088
rect 25455 36057 25467 36060
rect 25409 36051 25467 36057
rect 26050 36048 26056 36060
rect 26108 36048 26114 36100
rect 26329 36091 26387 36097
rect 26329 36057 26341 36091
rect 26375 36088 26387 36091
rect 26510 36088 26516 36100
rect 26375 36060 26516 36088
rect 26375 36057 26387 36060
rect 26329 36051 26387 36057
rect 26510 36048 26516 36060
rect 26568 36048 26574 36100
rect 27264 36088 27292 36119
rect 27798 36116 27804 36128
rect 27856 36116 27862 36168
rect 29178 36116 29184 36168
rect 29236 36156 29242 36168
rect 29917 36159 29975 36165
rect 29917 36156 29929 36159
rect 29236 36128 29929 36156
rect 29236 36116 29242 36128
rect 29917 36125 29929 36128
rect 29963 36125 29975 36159
rect 29917 36119 29975 36125
rect 26620 36060 27292 36088
rect 26142 36020 26148 36032
rect 25216 35992 26148 36020
rect 25041 35983 25099 35989
rect 26142 35980 26148 35992
rect 26200 36020 26206 36032
rect 26620 36020 26648 36060
rect 27338 36048 27344 36100
rect 27396 36048 27402 36100
rect 27433 36091 27491 36097
rect 27433 36057 27445 36091
rect 27479 36088 27491 36091
rect 27522 36088 27528 36100
rect 27479 36060 27528 36088
rect 27479 36057 27491 36060
rect 27433 36051 27491 36057
rect 27522 36048 27528 36060
rect 27580 36048 27586 36100
rect 28166 36048 28172 36100
rect 28224 36048 28230 36100
rect 28810 36048 28816 36100
rect 28868 36088 28874 36100
rect 30024 36088 30052 36196
rect 30300 36196 31401 36224
rect 30300 36165 30328 36196
rect 31389 36193 31401 36196
rect 31435 36224 31447 36227
rect 33594 36224 33600 36236
rect 31435 36196 33600 36224
rect 31435 36193 31447 36196
rect 31389 36187 31447 36193
rect 33594 36184 33600 36196
rect 33652 36184 33658 36236
rect 33796 36233 33824 36332
rect 33870 36320 33876 36332
rect 33928 36320 33934 36372
rect 34422 36320 34428 36372
rect 34480 36360 34486 36372
rect 35069 36363 35127 36369
rect 35069 36360 35081 36363
rect 34480 36332 35081 36360
rect 34480 36320 34486 36332
rect 35069 36329 35081 36332
rect 35115 36360 35127 36363
rect 36722 36360 36728 36372
rect 35115 36332 36728 36360
rect 35115 36329 35127 36332
rect 35069 36323 35127 36329
rect 36722 36320 36728 36332
rect 36780 36320 36786 36372
rect 36814 36320 36820 36372
rect 36872 36360 36878 36372
rect 38746 36360 38752 36372
rect 36872 36332 38752 36360
rect 36872 36320 36878 36332
rect 38746 36320 38752 36332
rect 38804 36320 38810 36372
rect 38930 36320 38936 36372
rect 38988 36320 38994 36372
rect 40681 36363 40739 36369
rect 40681 36329 40693 36363
rect 40727 36360 40739 36363
rect 41138 36360 41144 36372
rect 40727 36332 41144 36360
rect 40727 36329 40739 36332
rect 40681 36323 40739 36329
rect 41138 36320 41144 36332
rect 41196 36320 41202 36372
rect 42334 36360 42340 36372
rect 41708 36332 42340 36360
rect 34882 36252 34888 36304
rect 34940 36292 34946 36304
rect 35618 36292 35624 36304
rect 34940 36264 35624 36292
rect 34940 36252 34946 36264
rect 35618 36252 35624 36264
rect 35676 36292 35682 36304
rect 37274 36292 37280 36304
rect 35676 36264 37280 36292
rect 35676 36252 35682 36264
rect 37274 36252 37280 36264
rect 37332 36252 37338 36304
rect 37369 36295 37427 36301
rect 37369 36261 37381 36295
rect 37415 36292 37427 36295
rect 37415 36264 37688 36292
rect 37415 36261 37427 36264
rect 37369 36255 37427 36261
rect 33781 36227 33839 36233
rect 33781 36193 33793 36227
rect 33827 36193 33839 36227
rect 33781 36187 33839 36193
rect 35342 36184 35348 36236
rect 35400 36224 35406 36236
rect 36262 36224 36268 36236
rect 35400 36196 36268 36224
rect 35400 36184 35406 36196
rect 36262 36184 36268 36196
rect 36320 36224 36326 36236
rect 37660 36224 37688 36264
rect 37734 36252 37740 36304
rect 37792 36292 37798 36304
rect 38194 36292 38200 36304
rect 37792 36264 38200 36292
rect 37792 36252 37798 36264
rect 38194 36252 38200 36264
rect 38252 36252 38258 36304
rect 38473 36295 38531 36301
rect 38473 36261 38485 36295
rect 38519 36292 38531 36295
rect 40126 36292 40132 36304
rect 38519 36264 40132 36292
rect 38519 36261 38531 36264
rect 38473 36255 38531 36261
rect 40126 36252 40132 36264
rect 40184 36252 40190 36304
rect 41708 36236 41736 36332
rect 42334 36320 42340 36332
rect 42392 36320 42398 36372
rect 42610 36320 42616 36372
rect 42668 36360 42674 36372
rect 43349 36363 43407 36369
rect 43349 36360 43361 36363
rect 42668 36332 43361 36360
rect 42668 36320 42674 36332
rect 43349 36329 43361 36332
rect 43395 36329 43407 36363
rect 43349 36323 43407 36329
rect 41690 36224 41696 36236
rect 36320 36196 37412 36224
rect 37660 36196 40080 36224
rect 36320 36184 36326 36196
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36125 30343 36159
rect 30285 36119 30343 36125
rect 30466 36116 30472 36168
rect 30524 36116 30530 36168
rect 30745 36159 30803 36165
rect 30745 36125 30757 36159
rect 30791 36156 30803 36159
rect 31205 36159 31263 36165
rect 31205 36156 31217 36159
rect 30791 36128 31217 36156
rect 30791 36125 30803 36128
rect 30745 36119 30803 36125
rect 31205 36125 31217 36128
rect 31251 36156 31263 36159
rect 31478 36156 31484 36168
rect 31251 36128 31484 36156
rect 31251 36125 31263 36128
rect 31205 36119 31263 36125
rect 31478 36116 31484 36128
rect 31536 36116 31542 36168
rect 31573 36159 31631 36165
rect 31573 36125 31585 36159
rect 31619 36156 31631 36159
rect 33873 36159 33931 36165
rect 31619 36128 33732 36156
rect 31619 36125 31631 36128
rect 31573 36119 31631 36125
rect 30650 36088 30656 36100
rect 28868 36060 29776 36088
rect 30024 36060 30656 36088
rect 28868 36048 28874 36060
rect 26200 35992 26648 36020
rect 26200 35980 26206 35992
rect 26694 35980 26700 36032
rect 26752 36020 26758 36032
rect 27065 36023 27123 36029
rect 27065 36020 27077 36023
rect 26752 35992 27077 36020
rect 26752 35980 26758 35992
rect 27065 35989 27077 35992
rect 27111 35989 27123 36023
rect 27065 35983 27123 35989
rect 29089 36023 29147 36029
rect 29089 35989 29101 36023
rect 29135 36020 29147 36023
rect 29638 36020 29644 36032
rect 29135 35992 29644 36020
rect 29135 35989 29147 35992
rect 29089 35983 29147 35989
rect 29638 35980 29644 35992
rect 29696 35980 29702 36032
rect 29748 36020 29776 36060
rect 30650 36048 30656 36060
rect 30708 36048 30714 36100
rect 30834 36048 30840 36100
rect 30892 36088 30898 36100
rect 31588 36088 31616 36119
rect 30892 36060 31616 36088
rect 32769 36091 32827 36097
rect 30892 36048 30898 36060
rect 32769 36057 32781 36091
rect 32815 36057 32827 36091
rect 33704 36088 33732 36128
rect 33873 36125 33885 36159
rect 33919 36156 33931 36159
rect 34238 36156 34244 36168
rect 33919 36128 34244 36156
rect 33919 36125 33931 36128
rect 33873 36119 33931 36125
rect 34238 36116 34244 36128
rect 34296 36116 34302 36168
rect 34885 36159 34943 36165
rect 34885 36125 34897 36159
rect 34931 36156 34943 36159
rect 34931 36128 35204 36156
rect 34931 36125 34943 36128
rect 34885 36119 34943 36125
rect 35176 36100 35204 36128
rect 35894 36116 35900 36168
rect 35952 36116 35958 36168
rect 36722 36116 36728 36168
rect 36780 36116 36786 36168
rect 36814 36116 36820 36168
rect 36872 36156 36878 36168
rect 37016 36165 37044 36196
rect 37274 36165 37280 36168
rect 37001 36159 37059 36165
rect 36872 36128 36917 36156
rect 36872 36116 36878 36128
rect 37001 36125 37013 36159
rect 37047 36125 37059 36159
rect 37001 36119 37059 36125
rect 37231 36159 37280 36165
rect 37231 36125 37243 36159
rect 37277 36125 37280 36159
rect 37231 36119 37280 36125
rect 37274 36116 37280 36119
rect 37332 36116 37338 36168
rect 34974 36088 34980 36100
rect 33704 36060 34980 36088
rect 32769 36051 32827 36057
rect 30282 36020 30288 36032
rect 29748 35992 30288 36020
rect 30282 35980 30288 35992
rect 30340 35980 30346 36032
rect 30374 35980 30380 36032
rect 30432 36020 30438 36032
rect 31110 36020 31116 36032
rect 30432 35992 31116 36020
rect 30432 35980 30438 35992
rect 31110 35980 31116 35992
rect 31168 35980 31174 36032
rect 32784 36020 32812 36051
rect 34974 36048 34980 36060
rect 35032 36048 35038 36100
rect 35158 36048 35164 36100
rect 35216 36088 35222 36100
rect 36078 36088 36084 36100
rect 35216 36060 36084 36088
rect 35216 36048 35222 36060
rect 36078 36048 36084 36060
rect 36136 36048 36142 36100
rect 37093 36091 37151 36097
rect 37093 36057 37105 36091
rect 37139 36057 37151 36091
rect 37384 36088 37412 36196
rect 37734 36116 37740 36168
rect 37792 36156 37798 36168
rect 38010 36165 38016 36168
rect 37829 36159 37887 36165
rect 37829 36156 37841 36159
rect 37792 36128 37841 36156
rect 37792 36116 37798 36128
rect 37829 36125 37841 36128
rect 37875 36125 37887 36159
rect 37829 36119 37887 36125
rect 37977 36159 38016 36165
rect 37977 36125 37989 36159
rect 37977 36119 38016 36125
rect 38010 36116 38016 36119
rect 38068 36116 38074 36168
rect 38194 36116 38200 36168
rect 38252 36116 38258 36168
rect 38286 36116 38292 36168
rect 38344 36165 38350 36168
rect 38344 36156 38352 36165
rect 38344 36128 38389 36156
rect 38344 36119 38352 36128
rect 38344 36116 38350 36119
rect 38746 36116 38752 36168
rect 38804 36156 38810 36168
rect 39117 36159 39175 36165
rect 39117 36156 39129 36159
rect 38804 36128 39129 36156
rect 38804 36116 38810 36128
rect 39117 36125 39129 36128
rect 39163 36156 39175 36159
rect 39390 36156 39396 36168
rect 39163 36128 39396 36156
rect 39163 36125 39175 36128
rect 39117 36119 39175 36125
rect 39390 36116 39396 36128
rect 39448 36116 39454 36168
rect 40052 36165 40080 36196
rect 40420 36196 41696 36224
rect 39485 36159 39543 36165
rect 39485 36125 39497 36159
rect 39531 36156 39543 36159
rect 40037 36159 40095 36165
rect 39531 36128 39620 36156
rect 39531 36125 39543 36128
rect 39485 36119 39543 36125
rect 38105 36091 38163 36097
rect 38105 36088 38117 36091
rect 37384 36060 38117 36088
rect 37093 36051 37151 36057
rect 38105 36057 38117 36060
rect 38151 36057 38163 36091
rect 38105 36051 38163 36057
rect 33505 36023 33563 36029
rect 33505 36020 33517 36023
rect 32784 35992 33517 36020
rect 33505 35989 33517 35992
rect 33551 35989 33563 36023
rect 33505 35983 33563 35989
rect 35250 35980 35256 36032
rect 35308 36020 35314 36032
rect 35526 36020 35532 36032
rect 35308 35992 35532 36020
rect 35308 35980 35314 35992
rect 35526 35980 35532 35992
rect 35584 36020 35590 36032
rect 35713 36023 35771 36029
rect 35713 36020 35725 36023
rect 35584 35992 35725 36020
rect 35584 35980 35590 35992
rect 35713 35989 35725 35992
rect 35759 35989 35771 36023
rect 37108 36020 37136 36051
rect 39206 36048 39212 36100
rect 39264 36048 39270 36100
rect 39298 36048 39304 36100
rect 39356 36048 39362 36100
rect 37458 36020 37464 36032
rect 37108 35992 37464 36020
rect 35713 35983 35771 35989
rect 37458 35980 37464 35992
rect 37516 35980 37522 36032
rect 38470 35980 38476 36032
rect 38528 36020 38534 36032
rect 39592 36020 39620 36128
rect 40037 36125 40049 36159
rect 40083 36125 40095 36159
rect 40037 36119 40095 36125
rect 40130 36159 40188 36165
rect 40130 36125 40142 36159
rect 40176 36125 40188 36159
rect 40130 36119 40188 36125
rect 39850 36048 39856 36100
rect 39908 36088 39914 36100
rect 40144 36088 40172 36119
rect 40218 36116 40224 36168
rect 40276 36156 40282 36168
rect 40420 36165 40448 36196
rect 41690 36184 41696 36196
rect 41748 36184 41754 36236
rect 40405 36159 40463 36165
rect 40405 36156 40417 36159
rect 40276 36128 40417 36156
rect 40276 36116 40282 36128
rect 40405 36125 40417 36128
rect 40451 36125 40463 36159
rect 40405 36119 40463 36125
rect 40494 36116 40500 36168
rect 40552 36165 40558 36168
rect 40552 36156 40560 36165
rect 41141 36159 41199 36165
rect 40552 36128 40597 36156
rect 40552 36119 40560 36128
rect 41141 36125 41153 36159
rect 41187 36156 41199 36159
rect 41230 36156 41236 36168
rect 41187 36128 41236 36156
rect 41187 36125 41199 36128
rect 41141 36119 41199 36125
rect 40552 36116 40558 36119
rect 41230 36116 41236 36128
rect 41288 36116 41294 36168
rect 41325 36159 41383 36165
rect 41325 36125 41337 36159
rect 41371 36156 41383 36159
rect 41414 36156 41420 36168
rect 41371 36128 41420 36156
rect 41371 36125 41383 36128
rect 41325 36119 41383 36125
rect 41414 36116 41420 36128
rect 41472 36116 41478 36168
rect 41506 36116 41512 36168
rect 41564 36156 41570 36168
rect 41874 36156 41880 36168
rect 41564 36128 41880 36156
rect 41564 36116 41570 36128
rect 41874 36116 41880 36128
rect 41932 36156 41938 36168
rect 41969 36159 42027 36165
rect 41969 36156 41981 36159
rect 41932 36128 41981 36156
rect 41932 36116 41938 36128
rect 41969 36125 41981 36128
rect 42015 36125 42027 36159
rect 41969 36119 42027 36125
rect 39908 36060 40172 36088
rect 39908 36048 39914 36060
rect 40310 36048 40316 36100
rect 40368 36048 40374 36100
rect 42236 36091 42294 36097
rect 42236 36057 42248 36091
rect 42282 36088 42294 36091
rect 42610 36088 42616 36100
rect 42282 36060 42616 36088
rect 42282 36057 42294 36060
rect 42236 36051 42294 36057
rect 42610 36048 42616 36060
rect 42668 36048 42674 36100
rect 41046 36020 41052 36032
rect 38528 35992 41052 36020
rect 38528 35980 38534 35992
rect 41046 35980 41052 35992
rect 41104 35980 41110 36032
rect 41509 36023 41567 36029
rect 41509 35989 41521 36023
rect 41555 36020 41567 36023
rect 41782 36020 41788 36032
rect 41555 35992 41788 36020
rect 41555 35989 41567 35992
rect 41509 35983 41567 35989
rect 41782 35980 41788 35992
rect 41840 35980 41846 36032
rect 1104 35930 43884 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 43884 35930
rect 1104 35856 43884 35878
rect 1302 35776 1308 35828
rect 1360 35816 1366 35828
rect 14553 35819 14611 35825
rect 1360 35788 12434 35816
rect 1360 35776 1366 35788
rect 12406 35748 12434 35788
rect 14553 35785 14565 35819
rect 14599 35816 14611 35819
rect 15562 35816 15568 35828
rect 14599 35788 15568 35816
rect 14599 35785 14611 35788
rect 14553 35779 14611 35785
rect 15562 35776 15568 35788
rect 15620 35776 15626 35828
rect 16114 35776 16120 35828
rect 16172 35816 16178 35828
rect 16482 35816 16488 35828
rect 16172 35788 16488 35816
rect 16172 35776 16178 35788
rect 16482 35776 16488 35788
rect 16540 35776 16546 35828
rect 16592 35788 19932 35816
rect 16592 35748 16620 35788
rect 17954 35748 17960 35760
rect 12406 35720 16620 35748
rect 17052 35720 17960 35748
rect 13998 35640 14004 35692
rect 14056 35680 14062 35692
rect 15013 35683 15071 35689
rect 15013 35680 15025 35683
rect 14056 35652 15025 35680
rect 14056 35640 14062 35652
rect 15013 35649 15025 35652
rect 15059 35649 15071 35683
rect 15013 35643 15071 35649
rect 15470 35640 15476 35692
rect 15528 35680 15534 35692
rect 17052 35689 17080 35720
rect 17954 35708 17960 35720
rect 18012 35708 18018 35760
rect 15933 35683 15991 35689
rect 15933 35680 15945 35683
rect 15528 35652 15945 35680
rect 15528 35640 15534 35652
rect 15933 35649 15945 35652
rect 15979 35649 15991 35683
rect 15933 35643 15991 35649
rect 17037 35683 17095 35689
rect 17037 35649 17049 35683
rect 17083 35649 17095 35683
rect 17037 35643 17095 35649
rect 17126 35640 17132 35692
rect 17184 35640 17190 35692
rect 17313 35683 17371 35689
rect 17313 35649 17325 35683
rect 17359 35680 17371 35683
rect 17773 35683 17831 35689
rect 17773 35680 17785 35683
rect 17359 35652 17785 35680
rect 17359 35649 17371 35652
rect 17313 35643 17371 35649
rect 17773 35649 17785 35652
rect 17819 35649 17831 35683
rect 18693 35683 18751 35689
rect 18693 35680 18705 35683
rect 17773 35643 17831 35649
rect 17972 35652 18705 35680
rect 13449 35615 13507 35621
rect 13449 35581 13461 35615
rect 13495 35612 13507 35615
rect 16666 35612 16672 35624
rect 13495 35584 16672 35612
rect 13495 35581 13507 35584
rect 13449 35575 13507 35581
rect 16666 35572 16672 35584
rect 16724 35572 16730 35624
rect 15197 35547 15255 35553
rect 15197 35513 15209 35547
rect 15243 35544 15255 35547
rect 16206 35544 16212 35556
rect 15243 35516 16212 35544
rect 15243 35513 15255 35516
rect 15197 35507 15255 35513
rect 16206 35504 16212 35516
rect 16264 35504 16270 35556
rect 17972 35553 18000 35652
rect 18693 35649 18705 35652
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 18414 35572 18420 35624
rect 18472 35572 18478 35624
rect 17957 35547 18015 35553
rect 17957 35513 17969 35547
rect 18003 35513 18015 35547
rect 17957 35507 18015 35513
rect 14001 35479 14059 35485
rect 14001 35445 14013 35479
rect 14047 35476 14059 35479
rect 16942 35476 16948 35488
rect 14047 35448 16948 35476
rect 14047 35445 14059 35448
rect 14001 35439 14059 35445
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 17218 35436 17224 35488
rect 17276 35476 17282 35488
rect 18782 35476 18788 35488
rect 17276 35448 18788 35476
rect 17276 35436 17282 35448
rect 18782 35436 18788 35448
rect 18840 35436 18846 35488
rect 19904 35476 19932 35788
rect 19978 35776 19984 35828
rect 20036 35776 20042 35828
rect 20901 35819 20959 35825
rect 20901 35785 20913 35819
rect 20947 35816 20959 35819
rect 21453 35819 21511 35825
rect 21453 35816 21465 35819
rect 20947 35788 21465 35816
rect 20947 35785 20959 35788
rect 20901 35779 20959 35785
rect 21453 35785 21465 35788
rect 21499 35816 21511 35819
rect 21542 35816 21548 35828
rect 21499 35788 21548 35816
rect 21499 35785 21511 35788
rect 21453 35779 21511 35785
rect 21542 35776 21548 35788
rect 21600 35776 21606 35828
rect 22462 35776 22468 35828
rect 22520 35816 22526 35828
rect 23937 35819 23995 35825
rect 23937 35816 23949 35819
rect 22520 35788 23949 35816
rect 22520 35776 22526 35788
rect 23937 35785 23949 35788
rect 23983 35785 23995 35819
rect 28994 35816 29000 35828
rect 23937 35779 23995 35785
rect 24136 35788 29000 35816
rect 22002 35708 22008 35760
rect 22060 35708 22066 35760
rect 22094 35708 22100 35760
rect 22152 35748 22158 35760
rect 22922 35748 22928 35760
rect 22152 35720 22928 35748
rect 22152 35708 22158 35720
rect 22664 35689 22692 35720
rect 22922 35708 22928 35720
rect 22980 35708 22986 35760
rect 23658 35748 23664 35760
rect 23032 35720 23664 35748
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35649 22339 35683
rect 22281 35643 22339 35649
rect 22649 35683 22707 35689
rect 22649 35649 22661 35683
rect 22695 35649 22707 35683
rect 22649 35643 22707 35649
rect 22296 35612 22324 35643
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 23032 35689 23060 35720
rect 23658 35708 23664 35720
rect 23716 35708 23722 35760
rect 23017 35683 23075 35689
rect 23017 35680 23029 35683
rect 22888 35652 23029 35680
rect 22888 35640 22894 35652
rect 23017 35649 23029 35652
rect 23063 35649 23075 35683
rect 23017 35643 23075 35649
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35680 23535 35683
rect 23934 35680 23940 35692
rect 23523 35652 23940 35680
rect 23523 35649 23535 35652
rect 23477 35643 23535 35649
rect 23934 35640 23940 35652
rect 23992 35680 23998 35692
rect 24136 35680 24164 35788
rect 28994 35776 29000 35788
rect 29052 35776 29058 35828
rect 29086 35776 29092 35828
rect 29144 35816 29150 35828
rect 29181 35819 29239 35825
rect 29181 35816 29193 35819
rect 29144 35788 29193 35816
rect 29144 35776 29150 35788
rect 29181 35785 29193 35788
rect 29227 35785 29239 35819
rect 29181 35779 29239 35785
rect 29270 35776 29276 35828
rect 29328 35816 29334 35828
rect 29730 35816 29736 35828
rect 29328 35788 29736 35816
rect 29328 35776 29334 35788
rect 29730 35776 29736 35788
rect 29788 35776 29794 35828
rect 30834 35776 30840 35828
rect 30892 35776 30898 35828
rect 31662 35776 31668 35828
rect 31720 35776 31726 35828
rect 32122 35776 32128 35828
rect 32180 35816 32186 35828
rect 35618 35816 35624 35828
rect 32180 35788 35624 35816
rect 32180 35776 32186 35788
rect 35618 35776 35624 35788
rect 35676 35776 35682 35828
rect 35802 35776 35808 35828
rect 35860 35816 35866 35828
rect 40310 35816 40316 35828
rect 35860 35788 40316 35816
rect 35860 35776 35866 35788
rect 24578 35708 24584 35760
rect 24636 35708 24642 35760
rect 25317 35751 25375 35757
rect 25317 35717 25329 35751
rect 25363 35748 25375 35751
rect 27154 35748 27160 35760
rect 25363 35720 27160 35748
rect 25363 35717 25375 35720
rect 25317 35711 25375 35717
rect 27154 35708 27160 35720
rect 27212 35708 27218 35760
rect 27522 35708 27528 35760
rect 27580 35748 27586 35760
rect 27706 35748 27712 35760
rect 27580 35720 27712 35748
rect 27580 35708 27586 35720
rect 27706 35708 27712 35720
rect 27764 35748 27770 35760
rect 30009 35751 30067 35757
rect 30009 35748 30021 35751
rect 27764 35720 30021 35748
rect 27764 35708 27770 35720
rect 30009 35717 30021 35720
rect 30055 35748 30067 35751
rect 30098 35748 30104 35760
rect 30055 35720 30104 35748
rect 30055 35717 30067 35720
rect 30009 35711 30067 35717
rect 30098 35708 30104 35720
rect 30156 35708 30162 35760
rect 31680 35748 31708 35776
rect 30300 35720 31708 35748
rect 32861 35751 32919 35757
rect 23992 35652 24164 35680
rect 24213 35683 24271 35689
rect 23992 35640 23998 35652
rect 24213 35649 24225 35683
rect 24259 35680 24271 35683
rect 24394 35680 24400 35692
rect 24259 35652 24400 35680
rect 24259 35649 24271 35652
rect 24213 35643 24271 35649
rect 24394 35640 24400 35652
rect 24452 35680 24458 35692
rect 26053 35683 26111 35689
rect 24452 35652 26004 35680
rect 24452 35640 24458 35652
rect 23290 35612 23296 35624
rect 22296 35584 23296 35612
rect 23290 35572 23296 35584
rect 23348 35612 23354 35624
rect 23566 35612 23572 35624
rect 23348 35584 23572 35612
rect 23348 35572 23354 35584
rect 23566 35572 23572 35584
rect 23624 35572 23630 35624
rect 24121 35615 24179 35621
rect 24121 35581 24133 35615
rect 24167 35612 24179 35615
rect 24302 35612 24308 35624
rect 24167 35584 24308 35612
rect 24167 35581 24179 35584
rect 24121 35575 24179 35581
rect 24302 35572 24308 35584
rect 24360 35572 24366 35624
rect 24489 35615 24547 35621
rect 24489 35581 24501 35615
rect 24535 35612 24547 35615
rect 25314 35612 25320 35624
rect 24535 35584 25320 35612
rect 24535 35581 24547 35584
rect 24489 35575 24547 35581
rect 25314 35572 25320 35584
rect 25372 35612 25378 35624
rect 25774 35612 25780 35624
rect 25372 35584 25780 35612
rect 25372 35572 25378 35584
rect 25774 35572 25780 35584
rect 25832 35572 25838 35624
rect 25976 35612 26004 35652
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 26234 35680 26240 35692
rect 26099 35652 26240 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 26234 35640 26240 35652
rect 26292 35680 26298 35692
rect 26602 35680 26608 35692
rect 26292 35652 26608 35680
rect 26292 35640 26298 35652
rect 26602 35640 26608 35652
rect 26660 35640 26666 35692
rect 27433 35683 27491 35689
rect 27433 35680 27445 35683
rect 26712 35652 27445 35680
rect 26712 35612 26740 35652
rect 27433 35649 27445 35652
rect 27479 35680 27491 35683
rect 28902 35680 28908 35692
rect 27479 35652 28908 35680
rect 27479 35649 27491 35652
rect 27433 35643 27491 35649
rect 28902 35640 28908 35652
rect 28960 35640 28966 35692
rect 29270 35640 29276 35692
rect 29328 35680 29334 35692
rect 29779 35683 29837 35689
rect 29779 35680 29791 35683
rect 29328 35652 29791 35680
rect 29328 35640 29334 35652
rect 29779 35649 29791 35652
rect 29825 35649 29837 35683
rect 29779 35643 29837 35649
rect 29914 35640 29920 35692
rect 29972 35640 29978 35692
rect 30190 35640 30196 35692
rect 30248 35640 30254 35692
rect 30300 35689 30328 35720
rect 32861 35717 32873 35751
rect 32907 35748 32919 35751
rect 33134 35748 33140 35760
rect 32907 35720 33140 35748
rect 32907 35717 32919 35720
rect 32861 35711 32919 35717
rect 33134 35708 33140 35720
rect 33192 35708 33198 35760
rect 35066 35748 35072 35760
rect 34256 35720 35072 35748
rect 30285 35683 30343 35689
rect 30285 35649 30297 35683
rect 30331 35649 30343 35683
rect 30285 35643 30343 35649
rect 30374 35640 30380 35692
rect 30432 35680 30438 35692
rect 31297 35683 31355 35689
rect 31297 35680 31309 35683
rect 30432 35652 31309 35680
rect 30432 35640 30438 35652
rect 31297 35649 31309 35652
rect 31343 35649 31355 35683
rect 31297 35643 31355 35649
rect 31665 35683 31723 35689
rect 31665 35649 31677 35683
rect 31711 35680 31723 35683
rect 31754 35680 31760 35692
rect 31711 35652 31760 35680
rect 31711 35649 31723 35652
rect 31665 35643 31723 35649
rect 31754 35640 31760 35652
rect 31812 35640 31818 35692
rect 32122 35640 32128 35692
rect 32180 35680 32186 35692
rect 32677 35683 32735 35689
rect 32677 35680 32689 35683
rect 32180 35652 32689 35680
rect 32180 35640 32186 35652
rect 32677 35649 32689 35652
rect 32723 35649 32735 35683
rect 32677 35643 32735 35649
rect 32769 35683 32827 35689
rect 32769 35649 32781 35683
rect 32815 35680 32827 35683
rect 32950 35680 32956 35692
rect 32815 35652 32956 35680
rect 32815 35649 32827 35652
rect 32769 35643 32827 35649
rect 32950 35640 32956 35652
rect 33008 35640 33014 35692
rect 33045 35683 33103 35689
rect 33045 35649 33057 35683
rect 33091 35649 33103 35683
rect 33045 35643 33103 35649
rect 25976 35584 26740 35612
rect 27341 35615 27399 35621
rect 27341 35581 27353 35615
rect 27387 35612 27399 35615
rect 27522 35612 27528 35624
rect 27387 35584 27528 35612
rect 27387 35581 27399 35584
rect 27341 35575 27399 35581
rect 27522 35572 27528 35584
rect 27580 35572 27586 35624
rect 27614 35572 27620 35624
rect 27672 35612 27678 35624
rect 27709 35615 27767 35621
rect 27709 35612 27721 35615
rect 27672 35584 27721 35612
rect 27672 35572 27678 35584
rect 27709 35581 27721 35584
rect 27755 35581 27767 35615
rect 27709 35575 27767 35581
rect 27801 35615 27859 35621
rect 27801 35581 27813 35615
rect 27847 35612 27859 35615
rect 28534 35612 28540 35624
rect 27847 35584 28540 35612
rect 27847 35581 27859 35584
rect 27801 35575 27859 35581
rect 28534 35572 28540 35584
rect 28592 35572 28598 35624
rect 28626 35572 28632 35624
rect 28684 35572 28690 35624
rect 28994 35572 29000 35624
rect 29052 35572 29058 35624
rect 29086 35572 29092 35624
rect 29144 35612 29150 35624
rect 29144 35584 31432 35612
rect 29144 35572 29150 35584
rect 26602 35504 26608 35556
rect 26660 35544 26666 35556
rect 31202 35544 31208 35556
rect 26660 35516 31208 35544
rect 26660 35504 26666 35516
rect 31202 35504 31208 35516
rect 31260 35504 31266 35556
rect 24578 35476 24584 35488
rect 19904 35448 24584 35476
rect 24578 35436 24584 35448
rect 24636 35436 24642 35488
rect 26878 35436 26884 35488
rect 26936 35476 26942 35488
rect 27157 35479 27215 35485
rect 27157 35476 27169 35479
rect 26936 35448 27169 35476
rect 26936 35436 26942 35448
rect 27157 35445 27169 35448
rect 27203 35445 27215 35479
rect 27157 35439 27215 35445
rect 29362 35436 29368 35488
rect 29420 35476 29426 35488
rect 29641 35479 29699 35485
rect 29641 35476 29653 35479
rect 29420 35448 29653 35476
rect 29420 35436 29426 35448
rect 29641 35445 29653 35448
rect 29687 35445 29699 35479
rect 29641 35439 29699 35445
rect 30006 35436 30012 35488
rect 30064 35476 30070 35488
rect 31018 35476 31024 35488
rect 30064 35448 31024 35476
rect 30064 35436 30070 35448
rect 31018 35436 31024 35448
rect 31076 35436 31082 35488
rect 31404 35476 31432 35584
rect 31938 35572 31944 35624
rect 31996 35612 32002 35624
rect 32398 35612 32404 35624
rect 31996 35584 32404 35612
rect 31996 35572 32002 35584
rect 32398 35572 32404 35584
rect 32456 35612 32462 35624
rect 33060 35612 33088 35643
rect 34146 35640 34152 35692
rect 34204 35680 34210 35692
rect 34256 35689 34284 35720
rect 35066 35708 35072 35720
rect 35124 35708 35130 35760
rect 35250 35708 35256 35760
rect 35308 35748 35314 35760
rect 35308 35720 36032 35748
rect 35308 35708 35314 35720
rect 36004 35692 36032 35720
rect 37182 35708 37188 35760
rect 37240 35748 37246 35760
rect 37737 35751 37795 35757
rect 37737 35748 37749 35751
rect 37240 35720 37749 35748
rect 37240 35708 37246 35720
rect 37737 35717 37749 35720
rect 37783 35717 37795 35751
rect 38470 35748 38476 35760
rect 37737 35711 37795 35717
rect 37844 35720 38476 35748
rect 34241 35683 34299 35689
rect 34241 35680 34253 35683
rect 34204 35652 34253 35680
rect 34204 35640 34210 35652
rect 34241 35649 34253 35652
rect 34287 35649 34299 35683
rect 34241 35643 34299 35649
rect 34882 35640 34888 35692
rect 34940 35640 34946 35692
rect 35158 35640 35164 35692
rect 35216 35640 35222 35692
rect 35805 35683 35863 35689
rect 35805 35680 35817 35683
rect 35360 35652 35817 35680
rect 32456 35584 33088 35612
rect 32456 35572 32462 35584
rect 33318 35572 33324 35624
rect 33376 35612 33382 35624
rect 33965 35615 34023 35621
rect 33965 35612 33977 35615
rect 33376 35584 33977 35612
rect 33376 35572 33382 35584
rect 33965 35581 33977 35584
rect 34011 35581 34023 35615
rect 33965 35575 34023 35581
rect 34974 35572 34980 35624
rect 35032 35572 35038 35624
rect 31478 35504 31484 35556
rect 31536 35544 31542 35556
rect 35250 35544 35256 35556
rect 31536 35516 35256 35544
rect 31536 35504 31542 35516
rect 35250 35504 35256 35516
rect 35308 35504 35314 35556
rect 35360 35553 35388 35652
rect 35805 35649 35817 35652
rect 35851 35649 35863 35683
rect 35805 35643 35863 35649
rect 35986 35640 35992 35692
rect 36044 35640 36050 35692
rect 36722 35640 36728 35692
rect 36780 35680 36786 35692
rect 37642 35689 37648 35692
rect 37461 35683 37519 35689
rect 37461 35680 37473 35683
rect 36780 35652 37473 35680
rect 36780 35640 36786 35652
rect 37461 35649 37473 35652
rect 37507 35649 37519 35683
rect 37461 35643 37519 35649
rect 37609 35683 37648 35689
rect 37609 35649 37621 35683
rect 37609 35643 37648 35649
rect 37642 35640 37648 35643
rect 37700 35640 37706 35692
rect 37844 35689 37872 35720
rect 38470 35708 38476 35720
rect 38528 35708 38534 35760
rect 38657 35751 38715 35757
rect 38657 35717 38669 35751
rect 38703 35748 38715 35751
rect 39022 35748 39028 35760
rect 38703 35720 39028 35748
rect 38703 35717 38715 35720
rect 38657 35711 38715 35717
rect 39022 35708 39028 35720
rect 39080 35708 39086 35760
rect 39684 35757 39712 35788
rect 40310 35776 40316 35788
rect 40368 35776 40374 35828
rect 41141 35819 41199 35825
rect 41141 35785 41153 35819
rect 41187 35816 41199 35819
rect 41230 35816 41236 35828
rect 41187 35788 41236 35816
rect 41187 35785 41199 35788
rect 41141 35779 41199 35785
rect 41230 35776 41236 35788
rect 41288 35776 41294 35828
rect 42610 35776 42616 35828
rect 42668 35776 42674 35828
rect 42702 35776 42708 35828
rect 42760 35816 42766 35828
rect 43257 35819 43315 35825
rect 43257 35816 43269 35819
rect 42760 35788 43269 35816
rect 42760 35776 42766 35788
rect 43257 35785 43269 35788
rect 43303 35785 43315 35819
rect 43257 35779 43315 35785
rect 39669 35751 39727 35757
rect 39669 35717 39681 35751
rect 39715 35717 39727 35751
rect 39669 35711 39727 35717
rect 37829 35683 37887 35689
rect 37829 35649 37841 35683
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 37967 35683 38025 35689
rect 37967 35649 37979 35683
rect 38013 35649 38025 35683
rect 39393 35683 39451 35689
rect 39393 35680 39405 35683
rect 37967 35643 38025 35649
rect 38120 35652 39405 35680
rect 36814 35572 36820 35624
rect 36872 35612 36878 35624
rect 37844 35612 37872 35643
rect 36872 35584 37872 35612
rect 36872 35572 36878 35584
rect 35345 35547 35403 35553
rect 35345 35513 35357 35547
rect 35391 35513 35403 35547
rect 35345 35507 35403 35513
rect 35802 35504 35808 35556
rect 35860 35544 35866 35556
rect 35897 35547 35955 35553
rect 35897 35544 35909 35547
rect 35860 35516 35909 35544
rect 35860 35504 35866 35516
rect 35897 35513 35909 35516
rect 35943 35513 35955 35547
rect 35897 35507 35955 35513
rect 36170 35504 36176 35556
rect 36228 35544 36234 35556
rect 37826 35544 37832 35556
rect 36228 35516 37832 35544
rect 36228 35504 36234 35516
rect 37826 35504 37832 35516
rect 37884 35504 37890 35556
rect 32398 35476 32404 35488
rect 31404 35448 32404 35476
rect 32398 35436 32404 35448
rect 32456 35436 32462 35488
rect 32490 35436 32496 35488
rect 32548 35436 32554 35488
rect 33870 35436 33876 35488
rect 33928 35476 33934 35488
rect 34057 35479 34115 35485
rect 34057 35476 34069 35479
rect 33928 35448 34069 35476
rect 33928 35436 33934 35448
rect 34057 35445 34069 35448
rect 34103 35445 34115 35479
rect 34057 35439 34115 35445
rect 34422 35436 34428 35488
rect 34480 35436 34486 35488
rect 34606 35436 34612 35488
rect 34664 35476 34670 35488
rect 34885 35479 34943 35485
rect 34885 35476 34897 35479
rect 34664 35448 34897 35476
rect 34664 35436 34670 35448
rect 34885 35445 34897 35448
rect 34931 35445 34943 35479
rect 34885 35439 34943 35445
rect 35066 35436 35072 35488
rect 35124 35476 35130 35488
rect 36630 35476 36636 35488
rect 35124 35448 36636 35476
rect 35124 35436 35130 35448
rect 36630 35436 36636 35448
rect 36688 35436 36694 35488
rect 37274 35436 37280 35488
rect 37332 35476 37338 35488
rect 37992 35476 38020 35643
rect 38120 35553 38148 35652
rect 39393 35649 39405 35652
rect 39439 35649 39451 35683
rect 39393 35643 39451 35649
rect 39482 35640 39488 35692
rect 39540 35680 39546 35692
rect 39540 35652 39585 35680
rect 39540 35640 39546 35652
rect 39758 35640 39764 35692
rect 39816 35640 39822 35692
rect 39899 35683 39957 35689
rect 39899 35649 39911 35683
rect 39945 35680 39957 35683
rect 40402 35680 40408 35692
rect 39945 35652 40408 35680
rect 39945 35649 39957 35652
rect 39899 35643 39957 35649
rect 40402 35640 40408 35652
rect 40460 35640 40466 35692
rect 40494 35640 40500 35692
rect 40552 35640 40558 35692
rect 40586 35640 40592 35692
rect 40644 35689 40650 35692
rect 40644 35683 40693 35689
rect 40644 35649 40647 35683
rect 40681 35649 40693 35683
rect 40644 35643 40693 35649
rect 40773 35683 40831 35689
rect 40773 35649 40785 35683
rect 40819 35649 40831 35683
rect 40773 35643 40831 35649
rect 40644 35640 40650 35643
rect 40310 35572 40316 35624
rect 40368 35612 40374 35624
rect 40788 35612 40816 35643
rect 40862 35640 40868 35692
rect 40920 35640 40926 35692
rect 40962 35683 41020 35689
rect 40962 35649 40974 35683
rect 41008 35649 41020 35683
rect 40962 35643 41020 35649
rect 40368 35584 40816 35612
rect 40368 35572 40374 35584
rect 38105 35547 38163 35553
rect 38105 35513 38117 35547
rect 38151 35513 38163 35547
rect 38105 35507 38163 35513
rect 40402 35504 40408 35556
rect 40460 35544 40466 35556
rect 40972 35544 41000 35643
rect 41782 35640 41788 35692
rect 41840 35640 41846 35692
rect 41969 35683 42027 35689
rect 41969 35649 41981 35683
rect 42015 35680 42027 35683
rect 42797 35683 42855 35689
rect 42797 35680 42809 35683
rect 42015 35652 42809 35680
rect 42015 35649 42027 35652
rect 41969 35643 42027 35649
rect 42797 35649 42809 35652
rect 42843 35649 42855 35683
rect 42797 35643 42855 35649
rect 41322 35572 41328 35624
rect 41380 35612 41386 35624
rect 41601 35615 41659 35621
rect 41601 35612 41613 35615
rect 41380 35584 41613 35612
rect 41380 35572 41386 35584
rect 41601 35581 41613 35584
rect 41647 35581 41659 35615
rect 41601 35575 41659 35581
rect 40460 35516 41000 35544
rect 40460 35504 40466 35516
rect 38194 35476 38200 35488
rect 37332 35448 38200 35476
rect 37332 35436 37338 35448
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 40037 35479 40095 35485
rect 40037 35445 40049 35479
rect 40083 35476 40095 35479
rect 40586 35476 40592 35488
rect 40083 35448 40592 35476
rect 40083 35445 40095 35448
rect 40037 35439 40095 35445
rect 40586 35436 40592 35448
rect 40644 35436 40650 35488
rect 1104 35386 43884 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 43884 35386
rect 1104 35312 43884 35334
rect 5994 35232 6000 35284
rect 6052 35272 6058 35284
rect 15378 35272 15384 35284
rect 6052 35244 15384 35272
rect 6052 35232 6058 35244
rect 15378 35232 15384 35244
rect 15436 35232 15442 35284
rect 15470 35232 15476 35284
rect 15528 35232 15534 35284
rect 16206 35232 16212 35284
rect 16264 35232 16270 35284
rect 20165 35275 20223 35281
rect 20165 35241 20177 35275
rect 20211 35272 20223 35275
rect 20806 35272 20812 35284
rect 20211 35244 20812 35272
rect 20211 35241 20223 35244
rect 20165 35235 20223 35241
rect 20806 35232 20812 35244
rect 20864 35232 20870 35284
rect 20898 35232 20904 35284
rect 20956 35272 20962 35284
rect 21913 35275 21971 35281
rect 21913 35272 21925 35275
rect 20956 35244 21925 35272
rect 20956 35232 20962 35244
rect 21913 35241 21925 35244
rect 21959 35241 21971 35275
rect 21913 35235 21971 35241
rect 23658 35232 23664 35284
rect 23716 35232 23722 35284
rect 23845 35275 23903 35281
rect 23845 35241 23857 35275
rect 23891 35272 23903 35275
rect 23891 35244 25360 35272
rect 23891 35241 23903 35244
rect 23845 35235 23903 35241
rect 4614 35164 4620 35216
rect 4672 35204 4678 35216
rect 24762 35204 24768 35216
rect 4672 35176 15240 35204
rect 4672 35164 4678 35176
rect 2866 35096 2872 35148
rect 2924 35136 2930 35148
rect 15010 35136 15016 35148
rect 2924 35108 15016 35136
rect 2924 35096 2930 35108
rect 15010 35096 15016 35108
rect 15068 35096 15074 35148
rect 15212 35136 15240 35176
rect 15488 35176 24768 35204
rect 15488 35136 15516 35176
rect 24762 35164 24768 35176
rect 24820 35164 24826 35216
rect 24854 35164 24860 35216
rect 24912 35164 24918 35216
rect 25332 35204 25360 35244
rect 26602 35232 26608 35284
rect 26660 35272 26666 35284
rect 27706 35272 27712 35284
rect 26660 35244 27712 35272
rect 26660 35232 26666 35244
rect 27706 35232 27712 35244
rect 27764 35232 27770 35284
rect 28534 35232 28540 35284
rect 28592 35272 28598 35284
rect 29546 35272 29552 35284
rect 28592 35244 29552 35272
rect 28592 35232 28598 35244
rect 29546 35232 29552 35244
rect 29604 35232 29610 35284
rect 30742 35232 30748 35284
rect 30800 35272 30806 35284
rect 30837 35275 30895 35281
rect 30837 35272 30849 35275
rect 30800 35244 30849 35272
rect 30800 35232 30806 35244
rect 30837 35241 30849 35244
rect 30883 35241 30895 35275
rect 30837 35235 30895 35241
rect 33321 35275 33379 35281
rect 33321 35241 33333 35275
rect 33367 35272 33379 35275
rect 33410 35272 33416 35284
rect 33367 35244 33416 35272
rect 33367 35241 33379 35244
rect 33321 35235 33379 35241
rect 33410 35232 33416 35244
rect 33468 35232 33474 35284
rect 33594 35232 33600 35284
rect 33652 35272 33658 35284
rect 33778 35272 33784 35284
rect 33652 35244 33784 35272
rect 33652 35232 33658 35244
rect 33778 35232 33784 35244
rect 33836 35232 33842 35284
rect 33870 35232 33876 35284
rect 33928 35272 33934 35284
rect 35802 35272 35808 35284
rect 33928 35244 35808 35272
rect 33928 35232 33934 35244
rect 35802 35232 35808 35244
rect 35860 35232 35866 35284
rect 36262 35232 36268 35284
rect 36320 35232 36326 35284
rect 36998 35232 37004 35284
rect 37056 35272 37062 35284
rect 37737 35275 37795 35281
rect 37056 35244 37504 35272
rect 37056 35232 37062 35244
rect 28166 35204 28172 35216
rect 25332 35176 28172 35204
rect 28166 35164 28172 35176
rect 28224 35164 28230 35216
rect 30098 35164 30104 35216
rect 30156 35204 30162 35216
rect 31846 35204 31852 35216
rect 30156 35176 31852 35204
rect 30156 35164 30162 35176
rect 31846 35164 31852 35176
rect 31904 35204 31910 35216
rect 32122 35204 32128 35216
rect 31904 35176 32128 35204
rect 31904 35164 31910 35176
rect 32122 35164 32128 35176
rect 32180 35164 32186 35216
rect 32398 35164 32404 35216
rect 32456 35204 32462 35216
rect 33962 35204 33968 35216
rect 32456 35176 33968 35204
rect 32456 35164 32462 35176
rect 33962 35164 33968 35176
rect 34020 35164 34026 35216
rect 34882 35164 34888 35216
rect 34940 35164 34946 35216
rect 36170 35204 36176 35216
rect 34992 35176 36176 35204
rect 15212 35108 15516 35136
rect 16114 35096 16120 35148
rect 16172 35096 16178 35148
rect 16408 35108 18000 35136
rect 14369 35071 14427 35077
rect 14369 35037 14381 35071
rect 14415 35068 14427 35071
rect 14550 35068 14556 35080
rect 14415 35040 14556 35068
rect 14415 35037 14427 35040
rect 14369 35031 14427 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 15102 35028 15108 35080
rect 15160 35028 15166 35080
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35037 15347 35071
rect 15289 35031 15347 35037
rect 14458 34960 14464 35012
rect 14516 34960 14522 35012
rect 14645 35003 14703 35009
rect 14645 34969 14657 35003
rect 14691 35000 14703 35003
rect 15194 35000 15200 35012
rect 14691 34972 15200 35000
rect 14691 34969 14703 34972
rect 14645 34963 14703 34969
rect 15194 34960 15200 34972
rect 15252 34960 15258 35012
rect 13722 34892 13728 34944
rect 13780 34892 13786 34944
rect 14553 34935 14611 34941
rect 14553 34901 14565 34935
rect 14599 34932 14611 34935
rect 15304 34932 15332 35031
rect 16298 35028 16304 35080
rect 16356 35068 16362 35080
rect 16408 35077 16436 35108
rect 17972 35080 18000 35108
rect 18782 35096 18788 35148
rect 18840 35136 18846 35148
rect 22554 35136 22560 35148
rect 18840 35108 22560 35136
rect 18840 35096 18846 35108
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 16356 35040 16405 35068
rect 16356 35028 16362 35040
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 16393 35031 16451 35037
rect 16577 35071 16635 35077
rect 16577 35037 16589 35071
rect 16623 35068 16635 35071
rect 16850 35068 16856 35080
rect 16623 35040 16856 35068
rect 16623 35037 16635 35040
rect 16577 35031 16635 35037
rect 16850 35028 16856 35040
rect 16908 35068 16914 35080
rect 17126 35068 17132 35080
rect 16908 35040 17132 35068
rect 16908 35028 16914 35040
rect 17126 35028 17132 35040
rect 17184 35028 17190 35080
rect 17954 35028 17960 35080
rect 18012 35028 18018 35080
rect 18046 35028 18052 35080
rect 18104 35028 18110 35080
rect 18138 35028 18144 35080
rect 18196 35068 18202 35080
rect 18233 35071 18291 35077
rect 18233 35068 18245 35071
rect 18196 35040 18245 35068
rect 18196 35028 18202 35040
rect 18233 35037 18245 35040
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 18322 35028 18328 35080
rect 18380 35028 18386 35080
rect 20732 35077 20760 35108
rect 22554 35096 22560 35108
rect 22612 35136 22618 35148
rect 23106 35136 23112 35148
rect 22612 35108 23112 35136
rect 22612 35096 22618 35108
rect 23106 35096 23112 35108
rect 23164 35096 23170 35148
rect 23569 35139 23627 35145
rect 23569 35105 23581 35139
rect 23615 35136 23627 35139
rect 23842 35136 23848 35148
rect 23615 35108 23848 35136
rect 23615 35105 23627 35108
rect 23569 35099 23627 35105
rect 23842 35096 23848 35108
rect 23900 35096 23906 35148
rect 24578 35096 24584 35148
rect 24636 35096 24642 35148
rect 24872 35136 24900 35164
rect 25777 35139 25835 35145
rect 24872 35108 25360 35136
rect 20717 35071 20775 35077
rect 20717 35037 20729 35071
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 21453 35071 21511 35077
rect 21453 35037 21465 35071
rect 21499 35068 21511 35071
rect 22002 35068 22008 35080
rect 21499 35040 22008 35068
rect 21499 35037 21511 35040
rect 21453 35031 21511 35037
rect 22002 35028 22008 35040
rect 22060 35028 22066 35080
rect 22094 35028 22100 35080
rect 22152 35028 22158 35080
rect 22189 35071 22247 35077
rect 22189 35037 22201 35071
rect 22235 35068 22247 35071
rect 22646 35068 22652 35080
rect 22235 35040 22652 35068
rect 22235 35037 22247 35040
rect 22189 35031 22247 35037
rect 22646 35028 22652 35040
rect 22704 35068 22710 35080
rect 22704 35040 23152 35068
rect 22704 35028 22710 35040
rect 16022 34960 16028 35012
rect 16080 35000 16086 35012
rect 16485 35003 16543 35009
rect 16485 35000 16497 35003
rect 16080 34972 16497 35000
rect 16080 34960 16086 34972
rect 16485 34969 16497 34972
rect 16531 34969 16543 35003
rect 20993 35003 21051 35009
rect 20993 35000 21005 35003
rect 16485 34963 16543 34969
rect 16592 34972 21005 35000
rect 14599 34904 15332 34932
rect 14599 34901 14611 34904
rect 14553 34895 14611 34901
rect 15378 34892 15384 34944
rect 15436 34932 15442 34944
rect 16592 34932 16620 34972
rect 20993 34969 21005 34972
rect 21039 34969 21051 35003
rect 20993 34963 21051 34969
rect 22462 34960 22468 35012
rect 22520 34960 22526 35012
rect 22557 35003 22615 35009
rect 22557 34969 22569 35003
rect 22603 35000 22615 35003
rect 22830 35000 22836 35012
rect 22603 34972 22836 35000
rect 22603 34969 22615 34972
rect 22557 34963 22615 34969
rect 22830 34960 22836 34972
rect 22888 34960 22894 35012
rect 15436 34904 16620 34932
rect 16853 34935 16911 34941
rect 15436 34892 15442 34904
rect 16853 34901 16865 34935
rect 16899 34932 16911 34935
rect 17126 34932 17132 34944
rect 16899 34904 17132 34932
rect 16899 34901 16911 34904
rect 16853 34895 16911 34901
rect 17126 34892 17132 34904
rect 17184 34892 17190 34944
rect 17218 34892 17224 34944
rect 17276 34932 17282 34944
rect 17313 34935 17371 34941
rect 17313 34932 17325 34935
rect 17276 34904 17325 34932
rect 17276 34892 17282 34904
rect 17313 34901 17325 34904
rect 17359 34901 17371 34935
rect 17313 34895 17371 34901
rect 17402 34892 17408 34944
rect 17460 34932 17466 34944
rect 17865 34935 17923 34941
rect 17865 34932 17877 34935
rect 17460 34904 17877 34932
rect 17460 34892 17466 34904
rect 17865 34901 17877 34904
rect 17911 34901 17923 34935
rect 17865 34895 17923 34901
rect 18506 34892 18512 34944
rect 18564 34932 18570 34944
rect 18785 34935 18843 34941
rect 18785 34932 18797 34935
rect 18564 34904 18797 34932
rect 18564 34892 18570 34904
rect 18785 34901 18797 34904
rect 18831 34901 18843 34935
rect 18785 34895 18843 34901
rect 19705 34935 19763 34941
rect 19705 34901 19717 34935
rect 19751 34932 19763 34935
rect 22094 34932 22100 34944
rect 19751 34904 22100 34932
rect 19751 34901 19763 34904
rect 19705 34895 19763 34901
rect 22094 34892 22100 34904
rect 22152 34892 22158 34944
rect 22480 34932 22508 34960
rect 22738 34932 22744 34944
rect 22480 34904 22744 34932
rect 22738 34892 22744 34904
rect 22796 34892 22802 34944
rect 23124 34932 23152 35040
rect 23198 35028 23204 35080
rect 23256 35068 23262 35080
rect 23661 35071 23719 35077
rect 23661 35068 23673 35071
rect 23256 35040 23673 35068
rect 23256 35028 23262 35040
rect 23661 35037 23673 35040
rect 23707 35068 23719 35071
rect 23934 35068 23940 35080
rect 23707 35040 23940 35068
rect 23707 35037 23719 35040
rect 23661 35031 23719 35037
rect 23934 35028 23940 35040
rect 23992 35028 23998 35080
rect 24854 35028 24860 35080
rect 24912 35068 24918 35080
rect 25332 35077 25360 35108
rect 25777 35105 25789 35139
rect 25823 35136 25835 35139
rect 26326 35136 26332 35148
rect 25823 35108 26332 35136
rect 25823 35105 25835 35108
rect 25777 35099 25835 35105
rect 26326 35096 26332 35108
rect 26384 35096 26390 35148
rect 27890 35136 27896 35148
rect 26436 35108 27896 35136
rect 25133 35071 25191 35077
rect 25133 35068 25145 35071
rect 24912 35040 25145 35068
rect 24912 35028 24918 35040
rect 25133 35037 25145 35040
rect 25179 35037 25191 35071
rect 25133 35031 25191 35037
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 25406 35028 25412 35080
rect 25464 35068 25470 35080
rect 25593 35071 25651 35077
rect 25593 35068 25605 35071
rect 25464 35040 25605 35068
rect 25464 35028 25470 35040
rect 25593 35037 25605 35040
rect 25639 35068 25651 35071
rect 25866 35068 25872 35080
rect 25639 35040 25872 35068
rect 25639 35037 25651 35040
rect 25593 35031 25651 35037
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 26050 35028 26056 35080
rect 26108 35068 26114 35080
rect 26436 35068 26464 35108
rect 26108 35040 26464 35068
rect 26108 35028 26114 35040
rect 26602 35028 26608 35080
rect 26660 35077 26666 35080
rect 26660 35071 26709 35077
rect 26660 35037 26663 35071
rect 26697 35037 26709 35071
rect 26660 35031 26709 35037
rect 26660 35028 26666 35031
rect 23290 34960 23296 35012
rect 23348 35000 23354 35012
rect 23385 35003 23443 35009
rect 23385 35000 23397 35003
rect 23348 34972 23397 35000
rect 23348 34960 23354 34972
rect 23385 34969 23397 34972
rect 23431 34969 23443 35003
rect 24394 35000 24400 35012
rect 23385 34963 23443 34969
rect 23492 34972 24400 35000
rect 23492 34932 23520 34972
rect 24394 34960 24400 34972
rect 24452 34960 24458 35012
rect 25884 35000 25912 35028
rect 25884 34972 26740 35000
rect 23124 34904 23520 34932
rect 23566 34892 23572 34944
rect 23624 34932 23630 34944
rect 26513 34935 26571 34941
rect 26513 34932 26525 34935
rect 23624 34904 26525 34932
rect 23624 34892 23630 34904
rect 26513 34901 26525 34904
rect 26559 34901 26571 34935
rect 26712 34932 26740 34972
rect 26786 34960 26792 35012
rect 26844 34960 26850 35012
rect 26896 35009 26924 35108
rect 27890 35096 27896 35108
rect 27948 35136 27954 35148
rect 28721 35139 28779 35145
rect 28721 35136 28733 35139
rect 27948 35108 28733 35136
rect 27948 35096 27954 35108
rect 28721 35105 28733 35108
rect 28767 35136 28779 35139
rect 33134 35136 33140 35148
rect 28767 35108 33140 35136
rect 28767 35105 28779 35108
rect 28721 35099 28779 35105
rect 33134 35096 33140 35108
rect 33192 35096 33198 35148
rect 34992 35136 35020 35176
rect 36170 35164 36176 35176
rect 36228 35164 36234 35216
rect 36280 35204 36308 35232
rect 37182 35204 37188 35216
rect 36280 35176 37188 35204
rect 37182 35164 37188 35176
rect 37240 35204 37246 35216
rect 37476 35204 37504 35244
rect 37737 35241 37749 35275
rect 37783 35272 37795 35275
rect 40494 35272 40500 35284
rect 37783 35244 40500 35272
rect 37783 35241 37795 35244
rect 37737 35235 37795 35241
rect 40494 35232 40500 35244
rect 40552 35232 40558 35284
rect 42889 35275 42947 35281
rect 42889 35272 42901 35275
rect 41386 35244 42901 35272
rect 37240 35176 37320 35204
rect 37476 35176 38424 35204
rect 37240 35164 37246 35176
rect 33520 35108 35020 35136
rect 35069 35139 35127 35145
rect 33520 35080 33548 35108
rect 35069 35105 35081 35139
rect 35115 35136 35127 35139
rect 36814 35136 36820 35148
rect 35115 35108 36820 35136
rect 35115 35105 35127 35108
rect 35069 35099 35127 35105
rect 36814 35096 36820 35108
rect 36872 35096 36878 35148
rect 36906 35096 36912 35148
rect 36964 35136 36970 35148
rect 36964 35108 37228 35136
rect 36964 35096 36970 35108
rect 27062 35068 27068 35080
rect 27023 35040 27068 35068
rect 27062 35028 27068 35040
rect 27120 35028 27126 35080
rect 27157 35071 27215 35077
rect 27157 35037 27169 35071
rect 27203 35037 27215 35071
rect 27157 35031 27215 35037
rect 26881 35003 26939 35009
rect 26881 34969 26893 35003
rect 26927 34969 26939 35003
rect 26881 34963 26939 34969
rect 27172 34932 27200 35031
rect 27798 35028 27804 35080
rect 27856 35068 27862 35080
rect 28261 35071 28319 35077
rect 28261 35068 28273 35071
rect 27856 35040 28273 35068
rect 27856 35028 27862 35040
rect 28261 35037 28273 35040
rect 28307 35037 28319 35071
rect 28261 35031 28319 35037
rect 28350 35028 28356 35080
rect 28408 35028 28414 35080
rect 29270 35028 29276 35080
rect 29328 35068 29334 35080
rect 29914 35068 29920 35080
rect 29328 35040 29920 35068
rect 29328 35028 29334 35040
rect 29914 35028 29920 35040
rect 29972 35028 29978 35080
rect 30098 35028 30104 35080
rect 30156 35028 30162 35080
rect 30282 35028 30288 35080
rect 30340 35028 30346 35080
rect 31113 35071 31171 35077
rect 31113 35037 31125 35071
rect 31159 35068 31171 35071
rect 31386 35068 31392 35080
rect 31159 35040 31392 35068
rect 31159 35037 31171 35040
rect 31113 35031 31171 35037
rect 31386 35028 31392 35040
rect 31444 35028 31450 35080
rect 31662 35028 31668 35080
rect 31720 35068 31726 35080
rect 32217 35071 32275 35077
rect 32217 35068 32229 35071
rect 31720 35040 32229 35068
rect 31720 35028 31726 35040
rect 32217 35037 32229 35040
rect 32263 35037 32275 35071
rect 32217 35031 32275 35037
rect 32401 35071 32459 35077
rect 32401 35037 32413 35071
rect 32447 35068 32459 35071
rect 32582 35068 32588 35080
rect 32447 35040 32588 35068
rect 32447 35037 32459 35040
rect 32401 35031 32459 35037
rect 32582 35028 32588 35040
rect 32640 35028 32646 35080
rect 32674 35028 32680 35080
rect 32732 35068 32738 35080
rect 33318 35068 33324 35080
rect 32732 35040 33324 35068
rect 32732 35028 32738 35040
rect 33318 35028 33324 35040
rect 33376 35028 33382 35080
rect 33502 35028 33508 35080
rect 33560 35028 33566 35080
rect 33594 35028 33600 35080
rect 33652 35028 33658 35080
rect 33778 35028 33784 35080
rect 33836 35028 33842 35080
rect 33873 35071 33931 35077
rect 33873 35037 33885 35071
rect 33919 35068 33931 35071
rect 33962 35068 33968 35080
rect 33919 35040 33968 35068
rect 33919 35037 33931 35040
rect 33873 35031 33931 35037
rect 33962 35028 33968 35040
rect 34020 35028 34026 35080
rect 35161 35071 35219 35077
rect 35161 35037 35173 35071
rect 35207 35037 35219 35071
rect 35161 35031 35219 35037
rect 28626 34960 28632 35012
rect 28684 34960 28690 35012
rect 29454 34960 29460 35012
rect 29512 35000 29518 35012
rect 29822 35000 29828 35012
rect 29512 34972 29828 35000
rect 29512 34960 29518 34972
rect 29822 34960 29828 34972
rect 29880 35000 29886 35012
rect 30009 35003 30067 35009
rect 30009 35000 30021 35003
rect 29880 34972 30021 35000
rect 29880 34960 29886 34972
rect 30009 34969 30021 34972
rect 30055 34969 30067 35003
rect 30009 34963 30067 34969
rect 31202 34960 31208 35012
rect 31260 35000 31266 35012
rect 32766 35000 32772 35012
rect 31260 34972 32772 35000
rect 31260 34960 31266 34972
rect 32766 34960 32772 34972
rect 32824 34960 32830 35012
rect 33410 34960 33416 35012
rect 33468 35000 33474 35012
rect 34514 35000 34520 35012
rect 33468 34972 34520 35000
rect 33468 34960 33474 34972
rect 34514 34960 34520 34972
rect 34572 34960 34578 35012
rect 34606 34960 34612 35012
rect 34664 35000 34670 35012
rect 35176 35000 35204 35031
rect 35342 35028 35348 35080
rect 35400 35068 35406 35080
rect 35437 35071 35495 35077
rect 35437 35068 35449 35071
rect 35400 35040 35449 35068
rect 35400 35028 35406 35040
rect 35437 35037 35449 35040
rect 35483 35037 35495 35071
rect 35437 35031 35495 35037
rect 35526 35028 35532 35080
rect 35584 35028 35590 35080
rect 36722 35028 36728 35080
rect 36780 35068 36786 35080
rect 37200 35077 37228 35108
rect 37093 35071 37151 35077
rect 37093 35068 37105 35071
rect 36780 35040 37105 35068
rect 36780 35028 36786 35040
rect 37093 35037 37105 35040
rect 37139 35037 37151 35071
rect 37093 35031 37151 35037
rect 37186 35071 37244 35077
rect 37186 35037 37198 35071
rect 37232 35037 37244 35071
rect 37292 35068 37320 35176
rect 38286 35096 38292 35148
rect 38344 35096 38350 35148
rect 38396 35136 38424 35176
rect 39482 35164 39488 35216
rect 39540 35204 39546 35216
rect 41386 35204 41414 35244
rect 42889 35241 42901 35244
rect 42935 35241 42947 35275
rect 42889 35235 42947 35241
rect 39540 35176 41414 35204
rect 39540 35164 39546 35176
rect 40402 35136 40408 35148
rect 38396 35108 40408 35136
rect 40402 35096 40408 35108
rect 40460 35096 40466 35148
rect 40586 35096 40592 35148
rect 40644 35096 40650 35148
rect 41506 35096 41512 35148
rect 41564 35096 41570 35148
rect 37369 35071 37427 35077
rect 37369 35068 37381 35071
rect 37292 35040 37381 35068
rect 37186 35031 37244 35037
rect 37369 35037 37381 35040
rect 37415 35037 37427 35071
rect 37369 35031 37427 35037
rect 37599 35071 37657 35077
rect 37599 35037 37611 35071
rect 37645 35068 37657 35071
rect 38194 35068 38200 35080
rect 37645 35040 38200 35068
rect 37645 35037 37657 35040
rect 37599 35031 37657 35037
rect 38194 35028 38200 35040
rect 38252 35028 38258 35080
rect 38381 35071 38439 35077
rect 38381 35037 38393 35071
rect 38427 35068 38439 35071
rect 38470 35068 38476 35080
rect 38427 35040 38476 35068
rect 38427 35037 38439 35040
rect 38381 35031 38439 35037
rect 38470 35028 38476 35040
rect 38528 35028 38534 35080
rect 38933 35071 38991 35077
rect 38933 35037 38945 35071
rect 38979 35068 38991 35071
rect 40126 35068 40132 35080
rect 38979 35040 40132 35068
rect 38979 35037 38991 35040
rect 38933 35031 38991 35037
rect 40126 35028 40132 35040
rect 40184 35028 40190 35080
rect 40681 35071 40739 35077
rect 40681 35037 40693 35071
rect 40727 35068 40739 35071
rect 41322 35068 41328 35080
rect 40727 35040 41328 35068
rect 40727 35037 40739 35040
rect 40681 35031 40739 35037
rect 41322 35028 41328 35040
rect 41380 35028 41386 35080
rect 34664 34972 35204 35000
rect 34664 34960 34670 34972
rect 35618 34960 35624 35012
rect 35676 35000 35682 35012
rect 35989 35003 36047 35009
rect 35989 35000 36001 35003
rect 35676 34972 36001 35000
rect 35676 34960 35682 34972
rect 35989 34969 36001 34972
rect 36035 34969 36047 35003
rect 35989 34963 36047 34969
rect 36170 34960 36176 35012
rect 36228 34960 36234 35012
rect 36354 34960 36360 35012
rect 36412 35000 36418 35012
rect 37461 35003 37519 35009
rect 37461 35000 37473 35003
rect 36412 34972 37473 35000
rect 36412 34960 36418 34972
rect 37461 34969 37473 34972
rect 37507 34969 37519 35003
rect 37461 34963 37519 34969
rect 37826 34960 37832 35012
rect 37884 35000 37890 35012
rect 39298 35000 39304 35012
rect 37884 34972 39304 35000
rect 37884 34960 37890 34972
rect 39298 34960 39304 34972
rect 39356 34960 39362 35012
rect 39485 35003 39543 35009
rect 39485 34969 39497 35003
rect 39531 35000 39543 35003
rect 39666 35000 39672 35012
rect 39531 34972 39672 35000
rect 39531 34969 39543 34972
rect 39485 34963 39543 34969
rect 39666 34960 39672 34972
rect 39724 35000 39730 35012
rect 40954 35000 40960 35012
rect 39724 34972 40960 35000
rect 39724 34960 39730 34972
rect 40954 34960 40960 34972
rect 41012 34960 41018 35012
rect 41754 35003 41812 35009
rect 41754 35000 41766 35003
rect 41386 34972 41766 35000
rect 26712 34904 27200 34932
rect 26513 34895 26571 34901
rect 27982 34892 27988 34944
rect 28040 34932 28046 34944
rect 28077 34935 28135 34941
rect 28077 34932 28089 34935
rect 28040 34904 28089 34932
rect 28040 34892 28046 34904
rect 28077 34901 28089 34904
rect 28123 34901 28135 34935
rect 28077 34895 28135 34901
rect 28166 34892 28172 34944
rect 28224 34932 28230 34944
rect 29733 34935 29791 34941
rect 29733 34932 29745 34935
rect 28224 34904 29745 34932
rect 28224 34892 28230 34904
rect 29733 34901 29745 34904
rect 29779 34901 29791 34935
rect 29733 34895 29791 34901
rect 32585 34935 32643 34941
rect 32585 34901 32597 34935
rect 32631 34932 32643 34935
rect 34698 34932 34704 34944
rect 32631 34904 34704 34932
rect 32631 34901 32643 34904
rect 32585 34895 32643 34901
rect 34698 34892 34704 34904
rect 34756 34892 34762 34944
rect 35802 34892 35808 34944
rect 35860 34932 35866 34944
rect 40494 34932 40500 34944
rect 35860 34904 40500 34932
rect 35860 34892 35866 34904
rect 40494 34892 40500 34904
rect 40552 34892 40558 34944
rect 41049 34935 41107 34941
rect 41049 34901 41061 34935
rect 41095 34932 41107 34935
rect 41386 34932 41414 34972
rect 41754 34969 41766 34972
rect 41800 34969 41812 35003
rect 41754 34963 41812 34969
rect 41095 34904 41414 34932
rect 41095 34901 41107 34904
rect 41049 34895 41107 34901
rect 1104 34842 43884 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 43884 34842
rect 1104 34768 43884 34790
rect 13998 34688 14004 34740
rect 14056 34688 14062 34740
rect 16298 34688 16304 34740
rect 16356 34688 16362 34740
rect 22097 34731 22155 34737
rect 22097 34728 22109 34731
rect 16408 34700 22109 34728
rect 15010 34620 15016 34672
rect 15068 34660 15074 34672
rect 16408 34660 16436 34700
rect 22097 34697 22109 34700
rect 22143 34697 22155 34731
rect 22097 34691 22155 34697
rect 23290 34688 23296 34740
rect 23348 34728 23354 34740
rect 27798 34728 27804 34740
rect 23348 34700 27804 34728
rect 23348 34688 23354 34700
rect 27798 34688 27804 34700
rect 27856 34688 27862 34740
rect 28994 34688 29000 34740
rect 29052 34688 29058 34740
rect 31662 34728 31668 34740
rect 29196 34700 31668 34728
rect 22922 34660 22928 34672
rect 15068 34632 16436 34660
rect 19444 34632 22928 34660
rect 15068 34620 15074 34632
rect 13814 34552 13820 34604
rect 13872 34552 13878 34604
rect 14458 34552 14464 34604
rect 14516 34552 14522 34604
rect 14553 34595 14611 34601
rect 14553 34561 14565 34595
rect 14599 34592 14611 34595
rect 14642 34592 14648 34604
rect 14599 34564 14648 34592
rect 14599 34561 14611 34564
rect 14553 34555 14611 34561
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 14737 34595 14795 34601
rect 14737 34561 14749 34595
rect 14783 34592 14795 34595
rect 15194 34592 15200 34604
rect 14783 34564 15200 34592
rect 14783 34561 14795 34564
rect 14737 34555 14795 34561
rect 15194 34552 15200 34564
rect 15252 34592 15258 34604
rect 15562 34592 15568 34604
rect 15252 34564 15568 34592
rect 15252 34552 15258 34564
rect 15562 34552 15568 34564
rect 15620 34552 15626 34604
rect 15841 34595 15899 34601
rect 15841 34561 15853 34595
rect 15887 34561 15899 34595
rect 15841 34555 15899 34561
rect 13633 34527 13691 34533
rect 13633 34493 13645 34527
rect 13679 34524 13691 34527
rect 14476 34524 14504 34552
rect 13679 34496 14504 34524
rect 14921 34527 14979 34533
rect 13679 34493 13691 34496
rect 13633 34487 13691 34493
rect 14921 34493 14933 34527
rect 14967 34524 14979 34527
rect 15102 34524 15108 34536
rect 14967 34496 15108 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 15102 34484 15108 34496
rect 15160 34524 15166 34536
rect 15856 34524 15884 34555
rect 15930 34552 15936 34604
rect 15988 34552 15994 34604
rect 16117 34595 16175 34601
rect 16117 34561 16129 34595
rect 16163 34592 16175 34595
rect 16574 34592 16580 34604
rect 16163 34564 16580 34592
rect 16163 34561 16175 34564
rect 16117 34555 16175 34561
rect 16574 34552 16580 34564
rect 16632 34552 16638 34604
rect 17126 34552 17132 34604
rect 17184 34552 17190 34604
rect 17310 34552 17316 34604
rect 17368 34552 17374 34604
rect 17402 34552 17408 34604
rect 17460 34552 17466 34604
rect 17586 34552 17592 34604
rect 17644 34592 17650 34604
rect 17865 34595 17923 34601
rect 17865 34592 17877 34595
rect 17644 34564 17877 34592
rect 17644 34552 17650 34564
rect 17865 34561 17877 34564
rect 17911 34592 17923 34595
rect 18414 34592 18420 34604
rect 17911 34564 18420 34592
rect 17911 34561 17923 34564
rect 17865 34555 17923 34561
rect 18414 34552 18420 34564
rect 18472 34552 18478 34604
rect 18506 34552 18512 34604
rect 18564 34592 18570 34604
rect 19444 34592 19472 34632
rect 18564 34564 19472 34592
rect 19521 34595 19579 34601
rect 18564 34552 18570 34564
rect 19521 34561 19533 34595
rect 19567 34592 19579 34595
rect 20070 34592 20076 34604
rect 19567 34564 20076 34592
rect 19567 34561 19579 34564
rect 19521 34555 19579 34561
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 20916 34601 20944 34632
rect 22922 34620 22928 34632
rect 22980 34620 22986 34672
rect 24213 34663 24271 34669
rect 24213 34629 24225 34663
rect 24259 34660 24271 34663
rect 26234 34660 26240 34672
rect 24259 34632 26240 34660
rect 24259 34629 24271 34632
rect 24213 34623 24271 34629
rect 26234 34620 26240 34632
rect 26292 34620 26298 34672
rect 27338 34620 27344 34672
rect 27396 34620 27402 34672
rect 27816 34660 27844 34688
rect 29086 34660 29092 34672
rect 27816 34632 29092 34660
rect 29086 34620 29092 34632
rect 29144 34620 29150 34672
rect 20533 34595 20591 34601
rect 20533 34561 20545 34595
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20901 34595 20959 34601
rect 20901 34561 20913 34595
rect 20947 34561 20959 34595
rect 20901 34555 20959 34561
rect 16758 34524 16764 34536
rect 15160 34496 16764 34524
rect 15160 34484 15166 34496
rect 16758 34484 16764 34496
rect 16816 34484 16822 34536
rect 16945 34527 17003 34533
rect 16945 34493 16957 34527
rect 16991 34524 17003 34527
rect 18141 34527 18199 34533
rect 18141 34524 18153 34527
rect 16991 34496 18153 34524
rect 16991 34493 17003 34496
rect 16945 34487 17003 34493
rect 18141 34493 18153 34496
rect 18187 34493 18199 34527
rect 20548 34524 20576 34555
rect 22278 34552 22284 34604
rect 22336 34552 22342 34604
rect 22373 34595 22431 34601
rect 22373 34561 22385 34595
rect 22419 34592 22431 34595
rect 23566 34592 23572 34604
rect 22419 34564 23572 34592
rect 22419 34561 22431 34564
rect 22373 34555 22431 34561
rect 23566 34552 23572 34564
rect 23624 34552 23630 34604
rect 24762 34552 24768 34604
rect 24820 34592 24826 34604
rect 24857 34595 24915 34601
rect 24857 34592 24869 34595
rect 24820 34564 24869 34592
rect 24820 34552 24826 34564
rect 24857 34561 24869 34564
rect 24903 34561 24915 34595
rect 24857 34555 24915 34561
rect 25130 34552 25136 34604
rect 25188 34592 25194 34604
rect 25409 34595 25467 34601
rect 25409 34592 25421 34595
rect 25188 34564 25421 34592
rect 25188 34552 25194 34564
rect 25409 34561 25421 34564
rect 25455 34561 25467 34595
rect 25409 34555 25467 34561
rect 25590 34552 25596 34604
rect 25648 34552 25654 34604
rect 25682 34552 25688 34604
rect 25740 34552 25746 34604
rect 25866 34552 25872 34604
rect 25924 34552 25930 34604
rect 27982 34552 27988 34604
rect 28040 34552 28046 34604
rect 28077 34595 28135 34601
rect 28077 34561 28089 34595
rect 28123 34592 28135 34595
rect 28166 34592 28172 34604
rect 28123 34564 28172 34592
rect 28123 34561 28135 34564
rect 28077 34555 28135 34561
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 28350 34552 28356 34604
rect 28408 34552 28414 34604
rect 29196 34592 29224 34700
rect 31662 34688 31668 34700
rect 31720 34688 31726 34740
rect 31754 34688 31760 34740
rect 31812 34688 31818 34740
rect 33502 34728 33508 34740
rect 32048 34700 33508 34728
rect 30834 34620 30840 34672
rect 30892 34620 30898 34672
rect 28966 34564 29224 34592
rect 20622 34524 20628 34536
rect 20548 34496 20628 34524
rect 18141 34487 18199 34493
rect 20622 34484 20628 34496
rect 20680 34484 20686 34536
rect 20806 34484 20812 34536
rect 20864 34524 20870 34536
rect 21361 34527 21419 34533
rect 21361 34524 21373 34527
rect 20864 34496 21373 34524
rect 20864 34484 20870 34496
rect 21361 34493 21373 34496
rect 21407 34524 21419 34527
rect 22649 34527 22707 34533
rect 22649 34524 22661 34527
rect 21407 34496 22661 34524
rect 21407 34493 21419 34496
rect 21361 34487 21419 34493
rect 22649 34493 22661 34496
rect 22695 34524 22707 34527
rect 23290 34524 23296 34536
rect 22695 34496 23296 34524
rect 22695 34493 22707 34496
rect 22649 34487 22707 34493
rect 23290 34484 23296 34496
rect 23348 34484 23354 34536
rect 23385 34527 23443 34533
rect 23385 34493 23397 34527
rect 23431 34493 23443 34527
rect 23385 34487 23443 34493
rect 20530 34416 20536 34468
rect 20588 34416 20594 34468
rect 20714 34416 20720 34468
rect 20772 34456 20778 34468
rect 23400 34456 23428 34487
rect 23658 34484 23664 34536
rect 23716 34484 23722 34536
rect 24118 34484 24124 34536
rect 24176 34524 24182 34536
rect 25222 34524 25228 34536
rect 24176 34496 25228 34524
rect 24176 34484 24182 34496
rect 25222 34484 25228 34496
rect 25280 34484 25286 34536
rect 25498 34484 25504 34536
rect 25556 34524 25562 34536
rect 26050 34524 26056 34536
rect 25556 34496 26056 34524
rect 25556 34484 25562 34496
rect 26050 34484 26056 34496
rect 26108 34484 26114 34536
rect 27430 34484 27436 34536
rect 27488 34524 27494 34536
rect 28445 34527 28503 34533
rect 28445 34524 28457 34527
rect 27488 34496 28457 34524
rect 27488 34484 27494 34496
rect 28445 34493 28457 34496
rect 28491 34524 28503 34527
rect 28966 34524 28994 34564
rect 29362 34552 29368 34604
rect 29420 34552 29426 34604
rect 30006 34552 30012 34604
rect 30064 34592 30070 34604
rect 30561 34595 30619 34601
rect 30561 34592 30573 34595
rect 30064 34564 30573 34592
rect 30064 34552 30070 34564
rect 30561 34561 30573 34564
rect 30607 34561 30619 34595
rect 30561 34555 30619 34561
rect 30745 34595 30803 34601
rect 30745 34561 30757 34595
rect 30791 34592 30803 34595
rect 30852 34592 30880 34620
rect 31389 34595 31447 34601
rect 30791 34564 30972 34592
rect 30791 34561 30803 34564
rect 30745 34555 30803 34561
rect 28491 34496 28994 34524
rect 28491 34493 28503 34496
rect 28445 34487 28503 34493
rect 29270 34484 29276 34536
rect 29328 34484 29334 34536
rect 29730 34484 29736 34536
rect 29788 34524 29794 34536
rect 29825 34527 29883 34533
rect 29825 34524 29837 34527
rect 29788 34496 29837 34524
rect 29788 34484 29794 34496
rect 29825 34493 29837 34496
rect 29871 34493 29883 34527
rect 29825 34487 29883 34493
rect 30837 34527 30895 34533
rect 30837 34493 30849 34527
rect 30883 34493 30895 34527
rect 30944 34524 30972 34564
rect 31389 34561 31401 34595
rect 31435 34592 31447 34595
rect 32048 34592 32076 34700
rect 33502 34688 33508 34700
rect 33560 34688 33566 34740
rect 33962 34728 33968 34740
rect 33612 34700 33968 34728
rect 33612 34660 33640 34700
rect 33962 34688 33968 34700
rect 34020 34688 34026 34740
rect 35342 34728 35348 34740
rect 35084 34700 35348 34728
rect 31435 34564 32076 34592
rect 32140 34632 33640 34660
rect 33873 34663 33931 34669
rect 31435 34561 31447 34564
rect 31389 34555 31447 34561
rect 31481 34527 31539 34533
rect 31481 34524 31493 34527
rect 30944 34496 31493 34524
rect 30837 34487 30895 34493
rect 31481 34493 31493 34496
rect 31527 34524 31539 34527
rect 32140 34524 32168 34632
rect 33873 34629 33885 34663
rect 33919 34660 33931 34663
rect 34054 34660 34060 34672
rect 33919 34632 34060 34660
rect 33919 34629 33931 34632
rect 33873 34623 33931 34629
rect 34054 34620 34060 34632
rect 34112 34620 34118 34672
rect 35084 34669 35112 34700
rect 35342 34688 35348 34700
rect 35400 34728 35406 34740
rect 38562 34728 38568 34740
rect 35400 34700 38568 34728
rect 35400 34688 35406 34700
rect 38562 34688 38568 34700
rect 38620 34728 38626 34740
rect 41969 34731 42027 34737
rect 41969 34728 41981 34731
rect 38620 34700 41981 34728
rect 38620 34688 38626 34700
rect 41969 34697 41981 34700
rect 42015 34697 42027 34731
rect 41969 34691 42027 34697
rect 42702 34688 42708 34740
rect 42760 34728 42766 34740
rect 43257 34731 43315 34737
rect 43257 34728 43269 34731
rect 42760 34700 43269 34728
rect 42760 34688 42766 34700
rect 43257 34697 43269 34700
rect 43303 34697 43315 34731
rect 43257 34691 43315 34697
rect 34609 34663 34667 34669
rect 34609 34629 34621 34663
rect 34655 34660 34667 34663
rect 35069 34663 35127 34669
rect 35069 34660 35081 34663
rect 34655 34632 35081 34660
rect 34655 34629 34667 34632
rect 34609 34623 34667 34629
rect 35069 34629 35081 34632
rect 35115 34629 35127 34663
rect 37829 34663 37887 34669
rect 37829 34660 37841 34663
rect 35069 34623 35127 34629
rect 36188 34632 37841 34660
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34592 32367 34595
rect 32766 34592 32772 34604
rect 32355 34564 32772 34592
rect 32355 34561 32367 34564
rect 32309 34555 32367 34561
rect 32766 34552 32772 34564
rect 32824 34592 32830 34604
rect 34624 34592 34652 34623
rect 36188 34604 36216 34632
rect 37829 34629 37841 34632
rect 37875 34660 37887 34663
rect 38102 34660 38108 34672
rect 37875 34632 38108 34660
rect 37875 34629 37887 34632
rect 37829 34623 37887 34629
rect 38102 34620 38108 34632
rect 38160 34620 38166 34672
rect 40310 34620 40316 34672
rect 40368 34620 40374 34672
rect 40494 34620 40500 34672
rect 40552 34660 40558 34672
rect 41417 34663 41475 34669
rect 41417 34660 41429 34663
rect 40552 34632 41429 34660
rect 40552 34620 40558 34632
rect 41417 34629 41429 34632
rect 41463 34629 41475 34663
rect 41417 34623 41475 34629
rect 36170 34592 36176 34604
rect 32824 34564 34652 34592
rect 35820 34564 36176 34592
rect 32824 34552 32830 34564
rect 31527 34496 32168 34524
rect 31527 34493 31539 34496
rect 31481 34487 31539 34493
rect 23676 34456 23704 34484
rect 28534 34456 28540 34468
rect 20772 34428 23428 34456
rect 23492 34428 28540 34456
rect 20772 34416 20778 34428
rect 13722 34348 13728 34400
rect 13780 34388 13786 34400
rect 20806 34388 20812 34400
rect 13780 34360 20812 34388
rect 13780 34348 13786 34360
rect 20806 34348 20812 34360
rect 20864 34348 20870 34400
rect 22554 34348 22560 34400
rect 22612 34348 22618 34400
rect 23290 34348 23296 34400
rect 23348 34388 23354 34400
rect 23492 34388 23520 34428
rect 28534 34416 28540 34428
rect 28592 34416 28598 34468
rect 30377 34459 30435 34465
rect 30377 34456 30389 34459
rect 29288 34428 30389 34456
rect 23348 34360 23520 34388
rect 23348 34348 23354 34360
rect 26510 34348 26516 34400
rect 26568 34348 26574 34400
rect 29288 34397 29316 34428
rect 30377 34425 30389 34428
rect 30423 34425 30435 34459
rect 30852 34456 30880 34487
rect 32214 34484 32220 34536
rect 32272 34524 32278 34536
rect 32272 34496 32996 34524
rect 32272 34484 32278 34496
rect 32674 34456 32680 34468
rect 30852 34428 32680 34456
rect 30377 34419 30435 34425
rect 32674 34416 32680 34428
rect 32732 34416 32738 34468
rect 32968 34456 32996 34496
rect 33042 34484 33048 34536
rect 33100 34484 33106 34536
rect 34238 34484 34244 34536
rect 34296 34524 34302 34536
rect 35820 34524 35848 34564
rect 36170 34552 36176 34564
rect 36228 34552 36234 34604
rect 36446 34552 36452 34604
rect 36504 34552 36510 34604
rect 36633 34595 36691 34601
rect 36633 34561 36645 34595
rect 36679 34592 36691 34595
rect 36722 34592 36728 34604
rect 36679 34564 36728 34592
rect 36679 34561 36691 34564
rect 36633 34555 36691 34561
rect 34296 34496 35848 34524
rect 35897 34527 35955 34533
rect 34296 34484 34302 34496
rect 35897 34493 35909 34527
rect 35943 34493 35955 34527
rect 35897 34487 35955 34493
rect 35912 34456 35940 34487
rect 36078 34484 36084 34536
rect 36136 34524 36142 34536
rect 36648 34524 36676 34555
rect 36722 34552 36728 34564
rect 36780 34552 36786 34604
rect 36814 34552 36820 34604
rect 36872 34592 36878 34604
rect 37550 34592 37556 34604
rect 36872 34564 37556 34592
rect 36872 34552 36878 34564
rect 37550 34552 37556 34564
rect 37608 34552 37614 34604
rect 37642 34552 37648 34604
rect 37700 34552 37706 34604
rect 37734 34552 37740 34604
rect 37792 34552 37798 34604
rect 37918 34552 37924 34604
rect 37976 34592 37982 34604
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 37976 34564 38025 34592
rect 37976 34552 37982 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 39022 34552 39028 34604
rect 39080 34592 39086 34604
rect 39586 34595 39644 34601
rect 39586 34592 39598 34595
rect 39080 34564 39598 34592
rect 39080 34552 39086 34564
rect 39586 34561 39598 34564
rect 39632 34561 39644 34595
rect 39586 34555 39644 34561
rect 40218 34552 40224 34604
rect 40276 34592 40282 34604
rect 40865 34595 40923 34601
rect 40865 34592 40877 34595
rect 40276 34564 40877 34592
rect 40276 34552 40282 34564
rect 40865 34561 40877 34564
rect 40911 34561 40923 34595
rect 40865 34555 40923 34561
rect 42794 34552 42800 34604
rect 42852 34552 42858 34604
rect 36136 34496 36676 34524
rect 36909 34527 36967 34533
rect 36136 34484 36142 34496
rect 36909 34493 36921 34527
rect 36955 34524 36967 34527
rect 38286 34524 38292 34536
rect 36955 34496 38292 34524
rect 36955 34493 36967 34496
rect 36909 34487 36967 34493
rect 38286 34484 38292 34496
rect 38344 34484 38350 34536
rect 39853 34527 39911 34533
rect 39853 34493 39865 34527
rect 39899 34493 39911 34527
rect 39853 34487 39911 34493
rect 38838 34456 38844 34468
rect 32968 34428 35848 34456
rect 35912 34428 38844 34456
rect 29273 34391 29331 34397
rect 29273 34357 29285 34391
rect 29319 34357 29331 34391
rect 29273 34351 29331 34357
rect 30834 34348 30840 34400
rect 30892 34388 30898 34400
rect 31389 34391 31447 34397
rect 31389 34388 31401 34391
rect 30892 34360 31401 34388
rect 30892 34348 30898 34360
rect 31389 34357 31401 34360
rect 31435 34388 31447 34391
rect 33686 34388 33692 34400
rect 31435 34360 33692 34388
rect 31435 34357 31447 34360
rect 31389 34351 31447 34357
rect 33686 34348 33692 34360
rect 33744 34348 33750 34400
rect 35820 34388 35848 34428
rect 38838 34416 38844 34428
rect 38896 34456 38902 34468
rect 38896 34428 38976 34456
rect 38896 34416 38902 34428
rect 37182 34388 37188 34400
rect 35820 34360 37188 34388
rect 37182 34348 37188 34360
rect 37240 34348 37246 34400
rect 37274 34348 37280 34400
rect 37332 34388 37338 34400
rect 37461 34391 37519 34397
rect 37461 34388 37473 34391
rect 37332 34360 37473 34388
rect 37332 34348 37338 34360
rect 37461 34357 37473 34360
rect 37507 34357 37519 34391
rect 37461 34351 37519 34357
rect 37550 34348 37556 34400
rect 37608 34388 37614 34400
rect 38470 34388 38476 34400
rect 37608 34360 38476 34388
rect 37608 34348 37614 34360
rect 38470 34348 38476 34360
rect 38528 34348 38534 34400
rect 38948 34388 38976 34428
rect 39868 34388 39896 34487
rect 40126 34484 40132 34536
rect 40184 34524 40190 34536
rect 40184 34496 42656 34524
rect 40184 34484 40190 34496
rect 42628 34456 42656 34496
rect 42702 34484 42708 34536
rect 42760 34484 42766 34536
rect 43070 34456 43076 34468
rect 42628 34428 43076 34456
rect 43070 34416 43076 34428
rect 43128 34416 43134 34468
rect 38948 34360 39896 34388
rect 40954 34348 40960 34400
rect 41012 34388 41018 34400
rect 42150 34388 42156 34400
rect 41012 34360 42156 34388
rect 41012 34348 41018 34360
rect 42150 34348 42156 34360
rect 42208 34348 42214 34400
rect 1104 34298 43884 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 43884 34298
rect 1104 34224 43884 34246
rect 13725 34187 13783 34193
rect 13725 34153 13737 34187
rect 13771 34184 13783 34187
rect 13814 34184 13820 34196
rect 13771 34156 13820 34184
rect 13771 34153 13783 34156
rect 13725 34147 13783 34153
rect 13814 34144 13820 34156
rect 13872 34144 13878 34196
rect 14458 34144 14464 34196
rect 14516 34144 14522 34196
rect 16850 34144 16856 34196
rect 16908 34144 16914 34196
rect 17310 34144 17316 34196
rect 17368 34184 17374 34196
rect 17773 34187 17831 34193
rect 17773 34184 17785 34187
rect 17368 34156 17785 34184
rect 17368 34144 17374 34156
rect 17773 34153 17785 34156
rect 17819 34153 17831 34187
rect 17773 34147 17831 34153
rect 22186 34144 22192 34196
rect 22244 34144 22250 34196
rect 24029 34187 24087 34193
rect 24029 34153 24041 34187
rect 24075 34184 24087 34187
rect 24210 34184 24216 34196
rect 24075 34156 24216 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 24210 34144 24216 34156
rect 24268 34144 24274 34196
rect 26786 34144 26792 34196
rect 26844 34184 26850 34196
rect 27062 34184 27068 34196
rect 26844 34156 27068 34184
rect 26844 34144 26850 34156
rect 27062 34144 27068 34156
rect 27120 34144 27126 34196
rect 29086 34144 29092 34196
rect 29144 34144 29150 34196
rect 29270 34144 29276 34196
rect 29328 34184 29334 34196
rect 29733 34187 29791 34193
rect 29733 34184 29745 34187
rect 29328 34156 29745 34184
rect 29328 34144 29334 34156
rect 29733 34153 29745 34156
rect 29779 34153 29791 34187
rect 29733 34147 29791 34153
rect 30742 34144 30748 34196
rect 30800 34184 30806 34196
rect 32214 34184 32220 34196
rect 30800 34156 32220 34184
rect 30800 34144 30806 34156
rect 32214 34144 32220 34156
rect 32272 34144 32278 34196
rect 32490 34144 32496 34196
rect 32548 34184 32554 34196
rect 32858 34184 32864 34196
rect 32548 34156 32864 34184
rect 32548 34144 32554 34156
rect 32858 34144 32864 34156
rect 32916 34184 32922 34196
rect 35986 34184 35992 34196
rect 32916 34156 35992 34184
rect 32916 34144 32922 34156
rect 35986 34144 35992 34156
rect 36044 34144 36050 34196
rect 38933 34187 38991 34193
rect 38933 34153 38945 34187
rect 38979 34184 38991 34187
rect 39022 34184 39028 34196
rect 38979 34156 39028 34184
rect 38979 34153 38991 34156
rect 38933 34147 38991 34153
rect 39022 34144 39028 34156
rect 39080 34144 39086 34196
rect 40954 34184 40960 34196
rect 39132 34156 40960 34184
rect 13262 34076 13268 34128
rect 13320 34116 13326 34128
rect 14369 34119 14427 34125
rect 14369 34116 14381 34119
rect 13320 34088 14381 34116
rect 13320 34076 13326 34088
rect 14369 34085 14381 34088
rect 14415 34085 14427 34119
rect 14369 34079 14427 34085
rect 20530 34076 20536 34128
rect 20588 34076 20594 34128
rect 22002 34076 22008 34128
rect 22060 34116 22066 34128
rect 25133 34119 25191 34125
rect 25133 34116 25145 34119
rect 22060 34088 25145 34116
rect 22060 34076 22066 34088
rect 25133 34085 25145 34088
rect 25179 34085 25191 34119
rect 26510 34116 26516 34128
rect 25133 34079 25191 34085
rect 25240 34088 26516 34116
rect 12713 34051 12771 34057
rect 12713 34017 12725 34051
rect 12759 34048 12771 34051
rect 17034 34048 17040 34060
rect 12759 34020 17040 34048
rect 12759 34017 12771 34020
rect 12713 34011 12771 34017
rect 17034 34008 17040 34020
rect 17092 34008 17098 34060
rect 18138 34008 18144 34060
rect 18196 34048 18202 34060
rect 18196 34020 18368 34048
rect 18196 34008 18202 34020
rect 18340 33992 18368 34020
rect 21082 34008 21088 34060
rect 21140 34048 21146 34060
rect 21140 34020 22876 34048
rect 21140 34008 21146 34020
rect 13170 33940 13176 33992
rect 13228 33940 13234 33992
rect 13262 33940 13268 33992
rect 13320 33940 13326 33992
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 13464 33844 13492 33943
rect 13538 33940 13544 33992
rect 13596 33940 13602 33992
rect 14274 33940 14280 33992
rect 14332 33940 14338 33992
rect 14553 33983 14611 33989
rect 14553 33949 14565 33983
rect 14599 33949 14611 33983
rect 14553 33943 14611 33949
rect 13556 33912 13584 33940
rect 14568 33912 14596 33943
rect 14642 33940 14648 33992
rect 14700 33940 14706 33992
rect 15930 33940 15936 33992
rect 15988 33980 15994 33992
rect 16666 33980 16672 33992
rect 15988 33952 16672 33980
rect 15988 33940 15994 33952
rect 16666 33940 16672 33952
rect 16724 33940 16730 33992
rect 16758 33940 16764 33992
rect 16816 33940 16822 33992
rect 17954 33940 17960 33992
rect 18012 33940 18018 33992
rect 18046 33940 18052 33992
rect 18104 33940 18110 33992
rect 18230 33940 18236 33992
rect 18288 33940 18294 33992
rect 18322 33940 18328 33992
rect 18380 33940 18386 33992
rect 18782 33940 18788 33992
rect 18840 33980 18846 33992
rect 18877 33983 18935 33989
rect 18877 33980 18889 33983
rect 18840 33952 18889 33980
rect 18840 33940 18846 33952
rect 18877 33949 18889 33952
rect 18923 33980 18935 33983
rect 21637 33983 21695 33989
rect 21637 33980 21649 33983
rect 18923 33952 21649 33980
rect 18923 33949 18935 33952
rect 18877 33943 18935 33949
rect 21637 33949 21649 33952
rect 21683 33949 21695 33983
rect 21637 33943 21695 33949
rect 22005 33983 22063 33989
rect 22005 33949 22017 33983
rect 22051 33980 22063 33983
rect 22848 33980 22876 34020
rect 22922 34008 22928 34060
rect 22980 34048 22986 34060
rect 23382 34048 23388 34060
rect 22980 34020 23388 34048
rect 22980 34008 22986 34020
rect 23382 34008 23388 34020
rect 23440 34048 23446 34060
rect 23845 34051 23903 34057
rect 23845 34048 23857 34051
rect 23440 34020 23857 34048
rect 23440 34008 23446 34020
rect 23845 34017 23857 34020
rect 23891 34048 23903 34051
rect 25240 34048 25268 34088
rect 26510 34076 26516 34088
rect 26568 34076 26574 34128
rect 26973 34119 27031 34125
rect 26973 34085 26985 34119
rect 27019 34116 27031 34119
rect 27525 34119 27583 34125
rect 27525 34116 27537 34119
rect 27019 34088 27537 34116
rect 27019 34085 27031 34088
rect 26973 34079 27031 34085
rect 27525 34085 27537 34088
rect 27571 34085 27583 34119
rect 27525 34079 27583 34085
rect 28166 34076 28172 34128
rect 28224 34116 28230 34128
rect 28224 34088 30021 34116
rect 28224 34076 28230 34088
rect 23891 34020 25268 34048
rect 23891 34017 23903 34020
rect 23845 34011 23903 34017
rect 25498 34008 25504 34060
rect 25556 34008 25562 34060
rect 26694 34048 26700 34060
rect 25792 34020 26700 34048
rect 23753 33983 23811 33989
rect 22051 33952 22784 33980
rect 22848 33952 23704 33980
rect 22051 33949 22063 33952
rect 22005 33943 22063 33949
rect 13556 33884 14596 33912
rect 13814 33844 13820 33856
rect 13464 33816 13820 33844
rect 13814 33804 13820 33816
rect 13872 33844 13878 33856
rect 14660 33844 14688 33940
rect 15102 33872 15108 33924
rect 15160 33912 15166 33924
rect 15381 33915 15439 33921
rect 15381 33912 15393 33915
rect 15160 33884 15393 33912
rect 15160 33872 15166 33884
rect 15381 33881 15393 33884
rect 15427 33912 15439 33915
rect 16025 33915 16083 33921
rect 16025 33912 16037 33915
rect 15427 33884 16037 33912
rect 15427 33881 15439 33884
rect 15381 33875 15439 33881
rect 16025 33881 16037 33884
rect 16071 33881 16083 33915
rect 16025 33875 16083 33881
rect 16209 33915 16267 33921
rect 16209 33881 16221 33915
rect 16255 33912 16267 33915
rect 16390 33912 16396 33924
rect 16255 33884 16396 33912
rect 16255 33881 16267 33884
rect 16209 33875 16267 33881
rect 13872 33816 14688 33844
rect 13872 33804 13878 33816
rect 15746 33804 15752 33856
rect 15804 33844 15810 33856
rect 15841 33847 15899 33853
rect 15841 33844 15853 33847
rect 15804 33816 15853 33844
rect 15804 33804 15810 33816
rect 15841 33813 15853 33816
rect 15887 33813 15899 33847
rect 16040 33844 16068 33875
rect 16390 33872 16396 33884
rect 16448 33872 16454 33924
rect 16574 33872 16580 33924
rect 16632 33912 16638 33924
rect 16945 33915 17003 33921
rect 16945 33912 16957 33915
rect 16632 33884 16957 33912
rect 16632 33872 16638 33884
rect 16945 33881 16957 33884
rect 16991 33881 17003 33915
rect 18248 33912 18276 33940
rect 19334 33912 19340 33924
rect 18248 33884 19340 33912
rect 16945 33875 17003 33881
rect 19334 33872 19340 33884
rect 19392 33872 19398 33924
rect 20898 33872 20904 33924
rect 20956 33872 20962 33924
rect 21821 33915 21879 33921
rect 21821 33881 21833 33915
rect 21867 33881 21879 33915
rect 21821 33875 21879 33881
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 22186 33912 22192 33924
rect 21959 33884 22192 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 16850 33844 16856 33856
rect 16040 33816 16856 33844
rect 15841 33807 15899 33813
rect 16850 33804 16856 33816
rect 16908 33804 16914 33856
rect 19978 33804 19984 33856
rect 20036 33804 20042 33856
rect 20438 33804 20444 33856
rect 20496 33804 20502 33856
rect 21836 33844 21864 33875
rect 22186 33872 22192 33884
rect 22244 33912 22250 33924
rect 22554 33912 22560 33924
rect 22244 33884 22560 33912
rect 22244 33872 22250 33884
rect 22554 33872 22560 33884
rect 22612 33872 22618 33924
rect 22756 33912 22784 33952
rect 23198 33912 23204 33924
rect 22756 33884 23204 33912
rect 23198 33872 23204 33884
rect 23256 33872 23262 33924
rect 23290 33872 23296 33924
rect 23348 33912 23354 33924
rect 23385 33915 23443 33921
rect 23385 33912 23397 33915
rect 23348 33884 23397 33912
rect 23348 33872 23354 33884
rect 23385 33881 23397 33884
rect 23431 33881 23443 33915
rect 23385 33875 23443 33881
rect 23477 33915 23535 33921
rect 23477 33881 23489 33915
rect 23523 33912 23535 33915
rect 23566 33912 23572 33924
rect 23523 33884 23572 33912
rect 23523 33881 23535 33884
rect 23477 33875 23535 33881
rect 23566 33872 23572 33884
rect 23624 33872 23630 33924
rect 23676 33912 23704 33952
rect 23753 33949 23765 33983
rect 23799 33980 23811 33983
rect 24394 33980 24400 33992
rect 23799 33952 24400 33980
rect 23799 33949 23811 33952
rect 23753 33943 23811 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 25314 33989 25320 33992
rect 25312 33980 25320 33989
rect 25275 33952 25320 33980
rect 25312 33943 25320 33952
rect 25314 33940 25320 33943
rect 25372 33940 25378 33992
rect 23676 33884 23796 33912
rect 23308 33844 23336 33872
rect 21836 33816 23336 33844
rect 23768 33844 23796 33884
rect 23842 33872 23848 33924
rect 23900 33912 23906 33924
rect 23900 33884 24716 33912
rect 23900 33872 23906 33884
rect 24394 33844 24400 33856
rect 23768 33816 24400 33844
rect 24394 33804 24400 33816
rect 24452 33844 24458 33856
rect 24581 33847 24639 33853
rect 24581 33844 24593 33847
rect 24452 33816 24593 33844
rect 24452 33804 24458 33816
rect 24581 33813 24593 33816
rect 24627 33813 24639 33847
rect 24688 33844 24716 33884
rect 25222 33872 25228 33924
rect 25280 33912 25286 33924
rect 25516 33921 25544 34008
rect 25792 33989 25820 34020
rect 26694 34008 26700 34020
rect 26752 34008 26758 34060
rect 27798 34048 27804 34060
rect 26896 34020 27804 34048
rect 25684 33983 25742 33989
rect 25684 33949 25696 33983
rect 25730 33949 25742 33983
rect 25684 33943 25742 33949
rect 25777 33983 25835 33989
rect 25777 33949 25789 33983
rect 25823 33949 25835 33983
rect 25777 33943 25835 33949
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 25280 33884 25421 33912
rect 25280 33872 25286 33884
rect 25409 33881 25421 33884
rect 25455 33881 25467 33915
rect 25409 33875 25467 33881
rect 25501 33915 25559 33921
rect 25501 33881 25513 33915
rect 25547 33881 25559 33915
rect 25501 33875 25559 33881
rect 25700 33912 25728 33943
rect 25866 33940 25872 33992
rect 25924 33980 25930 33992
rect 26543 33983 26601 33989
rect 26543 33980 26555 33983
rect 25924 33952 26555 33980
rect 25924 33940 25930 33952
rect 26543 33949 26555 33952
rect 26589 33980 26601 33983
rect 26896 33980 26924 34020
rect 27798 34008 27804 34020
rect 27856 34048 27862 34060
rect 27856 34020 28304 34048
rect 27856 34008 27862 34020
rect 26589 33952 26924 33980
rect 26589 33949 26601 33952
rect 26543 33943 26601 33949
rect 27062 33940 27068 33992
rect 27120 33940 27126 33992
rect 27706 33989 27712 33992
rect 27684 33983 27712 33989
rect 27684 33949 27696 33983
rect 27684 33943 27712 33949
rect 27706 33940 27712 33943
rect 27764 33940 27770 33992
rect 27890 33940 27896 33992
rect 27948 33940 27954 33992
rect 27982 33940 27988 33992
rect 28040 33989 28046 33992
rect 28040 33983 28079 33989
rect 28067 33949 28079 33983
rect 28040 33943 28079 33949
rect 28162 33983 28220 33989
rect 28162 33949 28174 33983
rect 28208 33979 28220 33983
rect 28276 33979 28304 34020
rect 28810 34008 28816 34060
rect 28868 34048 28874 34060
rect 28868 34020 28948 34048
rect 28868 34008 28874 34020
rect 28208 33951 28304 33979
rect 28920 33980 28948 34020
rect 29086 34008 29092 34060
rect 29144 34048 29150 34060
rect 29993 34048 30021 34088
rect 30098 34076 30104 34128
rect 30156 34116 30162 34128
rect 30156 34088 36768 34116
rect 30156 34076 30162 34088
rect 29144 34020 29960 34048
rect 29993 34020 33180 34048
rect 29144 34008 29150 34020
rect 29454 33980 29460 33992
rect 28920 33952 29460 33980
rect 28208 33949 28220 33951
rect 28162 33943 28220 33949
rect 28040 33940 28046 33943
rect 29454 33940 29460 33952
rect 29512 33940 29518 33992
rect 29546 33940 29552 33992
rect 29604 33980 29610 33992
rect 29932 33989 29960 34020
rect 29733 33983 29791 33989
rect 29733 33980 29745 33983
rect 29604 33952 29745 33980
rect 29604 33940 29610 33952
rect 29733 33949 29745 33952
rect 29779 33949 29791 33983
rect 29733 33943 29791 33949
rect 29917 33983 29975 33989
rect 29917 33949 29929 33983
rect 29963 33980 29975 33983
rect 30098 33980 30104 33992
rect 29963 33952 30104 33980
rect 29963 33949 29975 33952
rect 29917 33943 29975 33949
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 31478 33940 31484 33992
rect 31536 33980 31542 33992
rect 31573 33983 31631 33989
rect 31573 33980 31585 33983
rect 31536 33952 31585 33980
rect 31536 33940 31542 33952
rect 31573 33949 31585 33952
rect 31619 33949 31631 33983
rect 31573 33943 31631 33949
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33980 31815 33983
rect 31846 33980 31852 33992
rect 31803 33952 31852 33980
rect 31803 33949 31815 33952
rect 31757 33943 31815 33949
rect 31846 33940 31852 33952
rect 31904 33940 31910 33992
rect 32033 33983 32091 33989
rect 32033 33949 32045 33983
rect 32079 33980 32091 33983
rect 32582 33980 32588 33992
rect 32079 33952 32588 33980
rect 32079 33949 32091 33952
rect 32033 33943 32091 33949
rect 32582 33940 32588 33952
rect 32640 33940 32646 33992
rect 32858 33940 32864 33992
rect 32916 33980 32922 33992
rect 33152 33989 33180 34020
rect 33428 34020 36676 34048
rect 33428 33989 33456 34020
rect 33040 33983 33098 33989
rect 33040 33980 33052 33983
rect 32916 33952 33052 33980
rect 32916 33940 32922 33952
rect 33040 33949 33052 33952
rect 33086 33949 33098 33983
rect 33040 33943 33098 33949
rect 33137 33983 33195 33989
rect 33137 33949 33149 33983
rect 33183 33949 33195 33983
rect 33137 33943 33195 33949
rect 33412 33983 33470 33989
rect 33412 33949 33424 33983
rect 33458 33949 33470 33983
rect 33412 33943 33470 33949
rect 33505 33983 33563 33989
rect 33505 33949 33517 33983
rect 33551 33980 33563 33983
rect 34422 33980 34428 33992
rect 33551 33952 34428 33980
rect 33551 33949 33563 33952
rect 33505 33943 33563 33949
rect 34422 33940 34428 33952
rect 34480 33940 34486 33992
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 35802 33980 35808 33992
rect 34572 33952 35808 33980
rect 34572 33940 34578 33952
rect 35802 33940 35808 33952
rect 35860 33980 35866 33992
rect 35897 33983 35955 33989
rect 35897 33980 35909 33983
rect 35860 33952 35909 33980
rect 35860 33940 35866 33952
rect 35897 33949 35909 33952
rect 35943 33949 35955 33983
rect 35897 33943 35955 33949
rect 26050 33912 26056 33924
rect 25700 33884 26056 33912
rect 25700 33844 25728 33884
rect 26050 33872 26056 33884
rect 26108 33872 26114 33924
rect 27801 33915 27859 33921
rect 27801 33881 27813 33915
rect 27847 33912 27859 33915
rect 28718 33912 28724 33924
rect 27847 33884 28724 33912
rect 27847 33881 27859 33884
rect 27801 33875 27859 33881
rect 28718 33872 28724 33884
rect 28776 33872 28782 33924
rect 28810 33872 28816 33924
rect 28868 33872 28874 33924
rect 28902 33872 28908 33924
rect 28960 33912 28966 33924
rect 31389 33915 31447 33921
rect 31389 33912 31401 33915
rect 28960 33884 31401 33912
rect 28960 33872 28966 33884
rect 31389 33881 31401 33884
rect 31435 33881 31447 33915
rect 31864 33912 31892 33940
rect 32950 33912 32956 33924
rect 31864 33884 32956 33912
rect 31389 33875 31447 33881
rect 32950 33872 32956 33884
rect 33008 33912 33014 33924
rect 33229 33915 33287 33921
rect 33229 33912 33241 33915
rect 33008 33884 33241 33912
rect 33008 33872 33014 33884
rect 33229 33881 33241 33884
rect 33275 33881 33287 33915
rect 33229 33875 33287 33881
rect 33594 33872 33600 33924
rect 33652 33912 33658 33924
rect 33965 33915 34023 33921
rect 33965 33912 33977 33915
rect 33652 33884 33977 33912
rect 33652 33872 33658 33884
rect 33965 33881 33977 33884
rect 34011 33881 34023 33915
rect 33965 33875 34023 33881
rect 35161 33915 35219 33921
rect 35161 33881 35173 33915
rect 35207 33912 35219 33915
rect 35342 33912 35348 33924
rect 35207 33884 35348 33912
rect 35207 33881 35219 33884
rect 35161 33875 35219 33881
rect 24688 33816 25728 33844
rect 24581 33807 24639 33813
rect 26418 33804 26424 33856
rect 26476 33804 26482 33856
rect 26510 33804 26516 33856
rect 26568 33844 26574 33856
rect 26605 33847 26663 33853
rect 26605 33844 26617 33847
rect 26568 33816 26617 33844
rect 26568 33804 26574 33816
rect 26605 33813 26617 33816
rect 26651 33813 26663 33847
rect 26605 33807 26663 33813
rect 27614 33804 27620 33856
rect 27672 33844 27678 33856
rect 30006 33844 30012 33856
rect 27672 33816 30012 33844
rect 27672 33804 27678 33816
rect 30006 33804 30012 33816
rect 30064 33804 30070 33856
rect 30466 33804 30472 33856
rect 30524 33844 30530 33856
rect 30926 33844 30932 33856
rect 30524 33816 30932 33844
rect 30524 33804 30530 33816
rect 30926 33804 30932 33816
rect 30984 33804 30990 33856
rect 32861 33847 32919 33853
rect 32861 33813 32873 33847
rect 32907 33844 32919 33847
rect 33502 33844 33508 33856
rect 32907 33816 33508 33844
rect 32907 33813 32919 33816
rect 32861 33807 32919 33813
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 33980 33844 34008 33875
rect 35342 33872 35348 33884
rect 35400 33872 35406 33924
rect 36648 33912 36676 34020
rect 36740 33989 36768 34088
rect 37182 34076 37188 34128
rect 37240 34116 37246 34128
rect 38010 34116 38016 34128
rect 37240 34088 38016 34116
rect 37240 34076 37246 34088
rect 38010 34076 38016 34088
rect 38068 34076 38074 34128
rect 37461 34051 37519 34057
rect 37461 34017 37473 34051
rect 37507 34048 37519 34051
rect 39132 34048 39160 34156
rect 40954 34144 40960 34156
rect 41012 34144 41018 34196
rect 41046 34144 41052 34196
rect 41104 34184 41110 34196
rect 41104 34156 41414 34184
rect 41104 34144 41110 34156
rect 41386 34128 41414 34156
rect 41386 34088 41420 34128
rect 41414 34076 41420 34088
rect 41472 34076 41478 34128
rect 37507 34020 39160 34048
rect 37507 34017 37519 34020
rect 37461 34011 37519 34017
rect 36725 33983 36783 33989
rect 36725 33949 36737 33983
rect 36771 33949 36783 33983
rect 36725 33943 36783 33949
rect 36906 33940 36912 33992
rect 36964 33980 36970 33992
rect 37185 33983 37243 33989
rect 37185 33980 37197 33983
rect 36964 33952 37197 33980
rect 36964 33940 36970 33952
rect 37185 33949 37197 33952
rect 37231 33949 37243 33983
rect 37185 33943 37243 33949
rect 37642 33940 37648 33992
rect 37700 33980 37706 33992
rect 38105 33983 38163 33989
rect 38105 33980 38117 33983
rect 37700 33952 38117 33980
rect 37700 33940 37706 33952
rect 38105 33949 38117 33952
rect 38151 33949 38163 33983
rect 38105 33943 38163 33949
rect 38378 33940 38384 33992
rect 38436 33980 38442 33992
rect 38473 33983 38531 33989
rect 38473 33980 38485 33983
rect 38436 33952 38485 33980
rect 38436 33940 38442 33952
rect 38473 33949 38485 33952
rect 38519 33949 38531 33983
rect 38473 33943 38531 33949
rect 39114 33940 39120 33992
rect 39172 33940 39178 33992
rect 39393 33983 39451 33989
rect 39393 33949 39405 33983
rect 39439 33980 39451 33983
rect 39758 33980 39764 33992
rect 39439 33952 39764 33980
rect 39439 33949 39451 33952
rect 39393 33943 39451 33949
rect 39758 33940 39764 33952
rect 39816 33940 39822 33992
rect 40034 33940 40040 33992
rect 40092 33980 40098 33992
rect 41322 33980 41328 33992
rect 40092 33952 41328 33980
rect 40092 33940 40098 33952
rect 41322 33940 41328 33952
rect 41380 33980 41386 33992
rect 43162 33980 43168 33992
rect 41380 33952 43168 33980
rect 41380 33940 41386 33952
rect 43162 33940 43168 33952
rect 43220 33980 43226 33992
rect 43257 33983 43315 33989
rect 43257 33980 43269 33983
rect 43220 33952 43269 33980
rect 43220 33940 43226 33952
rect 43257 33949 43269 33952
rect 43303 33949 43315 33983
rect 43257 33943 43315 33949
rect 37090 33912 37096 33924
rect 36648 33884 37096 33912
rect 37090 33872 37096 33884
rect 37148 33872 37154 33924
rect 36446 33844 36452 33856
rect 33980 33816 36452 33844
rect 36446 33804 36452 33816
rect 36504 33804 36510 33856
rect 37182 33804 37188 33856
rect 37240 33844 37246 33856
rect 37660 33844 37688 33940
rect 38010 33872 38016 33924
rect 38068 33912 38074 33924
rect 38197 33915 38255 33921
rect 38197 33912 38209 33915
rect 38068 33884 38209 33912
rect 38068 33872 38074 33884
rect 38197 33881 38209 33884
rect 38243 33881 38255 33915
rect 38197 33875 38255 33881
rect 38289 33915 38347 33921
rect 38289 33881 38301 33915
rect 38335 33881 38347 33915
rect 38289 33875 38347 33881
rect 37240 33816 37688 33844
rect 37240 33804 37246 33816
rect 37918 33804 37924 33856
rect 37976 33804 37982 33856
rect 38102 33804 38108 33856
rect 38160 33844 38166 33856
rect 38304 33844 38332 33875
rect 38930 33872 38936 33924
rect 38988 33912 38994 33924
rect 40282 33915 40340 33921
rect 40282 33912 40294 33915
rect 38988 33884 40294 33912
rect 38988 33872 38994 33884
rect 40282 33881 40294 33884
rect 40328 33881 40340 33915
rect 42150 33912 42156 33924
rect 40282 33875 40340 33881
rect 41386 33884 42156 33912
rect 38378 33844 38384 33856
rect 38160 33816 38384 33844
rect 38160 33804 38166 33816
rect 38378 33804 38384 33816
rect 38436 33804 38442 33856
rect 38470 33804 38476 33856
rect 38528 33844 38534 33856
rect 39301 33847 39359 33853
rect 39301 33844 39313 33847
rect 38528 33816 39313 33844
rect 38528 33804 38534 33816
rect 39301 33813 39313 33816
rect 39347 33813 39359 33847
rect 39301 33807 39359 33813
rect 39390 33804 39396 33856
rect 39448 33844 39454 33856
rect 41386 33844 41414 33884
rect 42150 33872 42156 33884
rect 42208 33912 42214 33924
rect 42794 33912 42800 33924
rect 42208 33884 42800 33912
rect 42208 33872 42214 33884
rect 42794 33872 42800 33884
rect 42852 33872 42858 33924
rect 42978 33872 42984 33924
rect 43036 33921 43042 33924
rect 43036 33912 43048 33921
rect 43036 33884 43081 33912
rect 43036 33875 43048 33884
rect 43036 33872 43042 33875
rect 39448 33816 41414 33844
rect 39448 33804 39454 33816
rect 41874 33804 41880 33856
rect 41932 33804 41938 33856
rect 1104 33754 43884 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 43884 33754
rect 1104 33680 43884 33702
rect 12989 33643 13047 33649
rect 12989 33609 13001 33643
rect 13035 33640 13047 33643
rect 13538 33640 13544 33652
rect 13035 33612 13544 33640
rect 13035 33609 13047 33612
rect 12989 33603 13047 33609
rect 13538 33600 13544 33612
rect 13596 33600 13602 33652
rect 13633 33643 13691 33649
rect 13633 33609 13645 33643
rect 13679 33640 13691 33643
rect 13814 33640 13820 33652
rect 13679 33612 13820 33640
rect 13679 33609 13691 33612
rect 13633 33603 13691 33609
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 15102 33600 15108 33652
rect 15160 33600 15166 33652
rect 15562 33600 15568 33652
rect 15620 33600 15626 33652
rect 15930 33600 15936 33652
rect 15988 33640 15994 33652
rect 16209 33643 16267 33649
rect 16209 33640 16221 33643
rect 15988 33612 16221 33640
rect 15988 33600 15994 33612
rect 16209 33609 16221 33612
rect 16255 33609 16267 33643
rect 16209 33603 16267 33609
rect 16574 33600 16580 33652
rect 16632 33640 16638 33652
rect 17957 33643 18015 33649
rect 17957 33640 17969 33643
rect 16632 33612 17969 33640
rect 16632 33600 16638 33612
rect 17957 33609 17969 33612
rect 18003 33609 18015 33643
rect 17957 33603 18015 33609
rect 19978 33600 19984 33652
rect 20036 33640 20042 33652
rect 23566 33640 23572 33652
rect 20036 33612 23572 33640
rect 20036 33600 20042 33612
rect 23566 33600 23572 33612
rect 23624 33640 23630 33652
rect 24210 33640 24216 33652
rect 23624 33612 24216 33640
rect 23624 33600 23630 33612
rect 24210 33600 24216 33612
rect 24268 33600 24274 33652
rect 24489 33643 24547 33649
rect 24489 33609 24501 33643
rect 24535 33640 24547 33643
rect 24854 33640 24860 33652
rect 24535 33612 24860 33640
rect 24535 33609 24547 33612
rect 24489 33603 24547 33609
rect 24854 33600 24860 33612
rect 24912 33600 24918 33652
rect 24949 33643 25007 33649
rect 24949 33609 24961 33643
rect 24995 33640 25007 33643
rect 25682 33640 25688 33652
rect 24995 33612 25688 33640
rect 24995 33609 25007 33612
rect 24949 33603 25007 33609
rect 25682 33600 25688 33612
rect 25740 33600 25746 33652
rect 28258 33600 28264 33652
rect 28316 33640 28322 33652
rect 28445 33643 28503 33649
rect 28445 33640 28457 33643
rect 28316 33612 28457 33640
rect 28316 33600 28322 33612
rect 28445 33609 28457 33612
rect 28491 33609 28503 33643
rect 28445 33603 28503 33609
rect 28534 33600 28540 33652
rect 28592 33640 28598 33652
rect 31202 33640 31208 33652
rect 28592 33612 31208 33640
rect 28592 33600 28598 33612
rect 31202 33600 31208 33612
rect 31260 33600 31266 33652
rect 31294 33600 31300 33652
rect 31352 33640 31358 33652
rect 31352 33612 31892 33640
rect 31352 33600 31358 33612
rect 15120 33572 15148 33600
rect 12728 33544 15148 33572
rect 17405 33575 17463 33581
rect 12728 33513 12756 33544
rect 17405 33541 17417 33575
rect 17451 33541 17463 33575
rect 24762 33572 24768 33584
rect 17405 33535 17463 33541
rect 19628 33544 24768 33572
rect 12253 33507 12311 33513
rect 12253 33473 12265 33507
rect 12299 33504 12311 33507
rect 12713 33507 12771 33513
rect 12713 33504 12725 33507
rect 12299 33476 12725 33504
rect 12299 33473 12311 33476
rect 12253 33467 12311 33473
rect 12713 33473 12725 33476
rect 12759 33473 12771 33507
rect 12713 33467 12771 33473
rect 12897 33507 12955 33513
rect 12897 33473 12909 33507
rect 12943 33473 12955 33507
rect 12897 33467 12955 33473
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 12912 33368 12940 33467
rect 13173 33439 13231 33445
rect 13173 33405 13185 33439
rect 13219 33436 13231 33439
rect 14108 33436 14136 33467
rect 15746 33464 15752 33516
rect 15804 33464 15810 33516
rect 16942 33464 16948 33516
rect 17000 33504 17006 33516
rect 17129 33507 17187 33513
rect 17129 33504 17141 33507
rect 17000 33476 17141 33504
rect 17000 33464 17006 33476
rect 17129 33473 17141 33476
rect 17175 33473 17187 33507
rect 17420 33504 17448 33535
rect 17865 33507 17923 33513
rect 17865 33504 17877 33507
rect 17420 33476 17877 33504
rect 17129 33467 17187 33473
rect 17865 33473 17877 33476
rect 17911 33473 17923 33507
rect 17865 33467 17923 33473
rect 18046 33464 18052 33516
rect 18104 33464 18110 33516
rect 19628 33448 19656 33544
rect 20162 33464 20168 33516
rect 20220 33504 20226 33516
rect 21100 33513 21128 33544
rect 24762 33532 24768 33544
rect 24820 33532 24826 33584
rect 25866 33572 25872 33584
rect 25056 33544 25872 33572
rect 20349 33507 20407 33513
rect 20349 33504 20361 33507
rect 20220 33476 20361 33504
rect 20220 33464 20226 33476
rect 20349 33473 20361 33476
rect 20395 33473 20407 33507
rect 20349 33467 20407 33473
rect 21085 33507 21143 33513
rect 21085 33473 21097 33507
rect 21131 33473 21143 33507
rect 21085 33467 21143 33473
rect 21266 33464 21272 33516
rect 21324 33464 21330 33516
rect 22554 33464 22560 33516
rect 22612 33504 22618 33516
rect 23385 33507 23443 33513
rect 23385 33504 23397 33507
rect 22612 33476 23397 33504
rect 22612 33464 22618 33476
rect 23385 33473 23397 33476
rect 23431 33473 23443 33507
rect 23385 33467 23443 33473
rect 23566 33464 23572 33516
rect 23624 33464 23630 33516
rect 24302 33464 24308 33516
rect 24360 33464 24366 33516
rect 24489 33507 24547 33513
rect 24489 33473 24501 33507
rect 24535 33504 24547 33507
rect 25056 33504 25084 33544
rect 25866 33532 25872 33544
rect 25924 33532 25930 33584
rect 27522 33532 27528 33584
rect 27580 33572 27586 33584
rect 29546 33572 29552 33584
rect 27580 33544 29552 33572
rect 27580 33532 27586 33544
rect 29546 33532 29552 33544
rect 29604 33532 29610 33584
rect 29733 33575 29791 33581
rect 29733 33541 29745 33575
rect 29779 33572 29791 33575
rect 30742 33572 30748 33584
rect 29779 33544 30748 33572
rect 29779 33541 29791 33544
rect 29733 33535 29791 33541
rect 30742 33532 30748 33544
rect 30800 33532 30806 33584
rect 30929 33575 30987 33581
rect 30929 33541 30941 33575
rect 30975 33572 30987 33575
rect 31018 33572 31024 33584
rect 30975 33544 31024 33572
rect 30975 33541 30987 33544
rect 30929 33535 30987 33541
rect 31018 33532 31024 33544
rect 31076 33532 31082 33584
rect 31113 33575 31171 33581
rect 31113 33541 31125 33575
rect 31159 33572 31171 33575
rect 31754 33572 31760 33584
rect 31159 33544 31760 33572
rect 31159 33541 31171 33544
rect 31113 33535 31171 33541
rect 31754 33532 31760 33544
rect 31812 33532 31818 33584
rect 31864 33572 31892 33612
rect 32398 33600 32404 33652
rect 32456 33600 32462 33652
rect 33686 33640 33692 33652
rect 32600 33612 33692 33640
rect 32600 33572 32628 33612
rect 33686 33600 33692 33612
rect 33744 33600 33750 33652
rect 33778 33600 33784 33652
rect 33836 33640 33842 33652
rect 37734 33640 37740 33652
rect 33836 33612 37740 33640
rect 33836 33600 33842 33612
rect 37734 33600 37740 33612
rect 37792 33600 37798 33652
rect 38930 33600 38936 33652
rect 38988 33600 38994 33652
rect 39022 33600 39028 33652
rect 39080 33640 39086 33652
rect 41598 33640 41604 33652
rect 39080 33612 41604 33640
rect 39080 33600 39086 33612
rect 41598 33600 41604 33612
rect 41656 33600 41662 33652
rect 43070 33600 43076 33652
rect 43128 33640 43134 33652
rect 43257 33643 43315 33649
rect 43257 33640 43269 33643
rect 43128 33612 43269 33640
rect 43128 33600 43134 33612
rect 43257 33609 43269 33612
rect 43303 33609 43315 33643
rect 43257 33603 43315 33609
rect 37461 33575 37519 33581
rect 37461 33572 37473 33575
rect 31864 33544 32628 33572
rect 32692 33544 37473 33572
rect 24535 33476 25084 33504
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 25130 33464 25136 33516
rect 25188 33464 25194 33516
rect 25225 33507 25283 33513
rect 25225 33473 25237 33507
rect 25271 33473 25283 33507
rect 25225 33467 25283 33473
rect 13219 33408 14136 33436
rect 13219 33405 13231 33408
rect 13173 33399 13231 33405
rect 14108 33368 14136 33408
rect 15841 33439 15899 33445
rect 15841 33405 15853 33439
rect 15887 33436 15899 33439
rect 16482 33436 16488 33448
rect 15887 33408 16488 33436
rect 15887 33405 15899 33408
rect 15841 33399 15899 33405
rect 16482 33396 16488 33408
rect 16540 33396 16546 33448
rect 17405 33439 17463 33445
rect 17405 33405 17417 33439
rect 17451 33436 17463 33439
rect 17678 33436 17684 33448
rect 17451 33408 17684 33436
rect 17451 33405 17463 33408
rect 17405 33399 17463 33405
rect 17678 33396 17684 33408
rect 17736 33396 17742 33448
rect 18690 33396 18696 33448
rect 18748 33436 18754 33448
rect 19153 33439 19211 33445
rect 19153 33436 19165 33439
rect 18748 33408 19165 33436
rect 18748 33396 18754 33408
rect 19153 33405 19165 33408
rect 19199 33405 19211 33439
rect 19153 33399 19211 33405
rect 19242 33396 19248 33448
rect 19300 33396 19306 33448
rect 19610 33396 19616 33448
rect 19668 33396 19674 33448
rect 20254 33396 20260 33448
rect 20312 33396 20318 33448
rect 20441 33439 20499 33445
rect 20441 33405 20453 33439
rect 20487 33405 20499 33439
rect 20441 33399 20499 33405
rect 20533 33439 20591 33445
rect 20533 33405 20545 33439
rect 20579 33436 20591 33439
rect 21177 33439 21235 33445
rect 21177 33436 21189 33439
rect 20579 33408 21189 33436
rect 20579 33405 20591 33408
rect 20533 33399 20591 33405
rect 21177 33405 21189 33408
rect 21223 33405 21235 33439
rect 22281 33439 22339 33445
rect 22281 33436 22293 33439
rect 21177 33399 21235 33405
rect 22066 33408 22293 33436
rect 20073 33371 20131 33377
rect 20073 33368 20085 33371
rect 12912 33340 13860 33368
rect 14108 33340 20085 33368
rect 13832 33309 13860 33340
rect 20073 33337 20085 33340
rect 20119 33337 20131 33371
rect 20073 33331 20131 33337
rect 13817 33303 13875 33309
rect 13817 33269 13829 33303
rect 13863 33300 13875 33303
rect 14366 33300 14372 33312
rect 13863 33272 14372 33300
rect 13863 33269 13875 33272
rect 13817 33263 13875 33269
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 17218 33260 17224 33312
rect 17276 33260 17282 33312
rect 18969 33303 19027 33309
rect 18969 33269 18981 33303
rect 19015 33300 19027 33303
rect 19150 33300 19156 33312
rect 19015 33272 19156 33300
rect 19015 33269 19027 33272
rect 18969 33263 19027 33269
rect 19150 33260 19156 33272
rect 19208 33260 19214 33312
rect 19334 33260 19340 33312
rect 19392 33300 19398 33312
rect 20346 33300 20352 33312
rect 19392 33272 20352 33300
rect 19392 33260 19398 33272
rect 20346 33260 20352 33272
rect 20404 33300 20410 33312
rect 20456 33300 20484 33399
rect 20714 33328 20720 33380
rect 20772 33368 20778 33380
rect 22066 33368 22094 33408
rect 22281 33405 22293 33408
rect 22327 33405 22339 33439
rect 22281 33399 22339 33405
rect 23750 33396 23756 33448
rect 23808 33436 23814 33448
rect 23845 33439 23903 33445
rect 23845 33436 23857 33439
rect 23808 33408 23857 33436
rect 23808 33396 23814 33408
rect 23845 33405 23857 33408
rect 23891 33405 23903 33439
rect 23845 33399 23903 33405
rect 24578 33396 24584 33448
rect 24636 33436 24642 33448
rect 24946 33436 24952 33448
rect 24636 33408 24952 33436
rect 24636 33396 24642 33408
rect 24946 33396 24952 33408
rect 25004 33436 25010 33448
rect 25240 33436 25268 33467
rect 25314 33464 25320 33516
rect 25372 33464 25378 33516
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33473 25559 33507
rect 25501 33467 25559 33473
rect 25004 33408 25268 33436
rect 25004 33396 25010 33408
rect 20772 33340 22094 33368
rect 22373 33371 22431 33377
rect 20772 33328 20778 33340
rect 22373 33337 22385 33371
rect 22419 33368 22431 33371
rect 22646 33368 22652 33380
rect 22419 33340 22652 33368
rect 22419 33337 22431 33340
rect 22373 33331 22431 33337
rect 22646 33328 22652 33340
rect 22704 33328 22710 33380
rect 23474 33328 23480 33380
rect 23532 33368 23538 33380
rect 23532 33340 24256 33368
rect 23532 33328 23538 33340
rect 21266 33300 21272 33312
rect 20404 33272 21272 33300
rect 20404 33260 20410 33272
rect 21266 33260 21272 33272
rect 21324 33260 21330 33312
rect 22462 33260 22468 33312
rect 22520 33260 22526 33312
rect 23382 33260 23388 33312
rect 23440 33300 23446 33312
rect 23753 33303 23811 33309
rect 23753 33300 23765 33303
rect 23440 33272 23765 33300
rect 23440 33260 23446 33272
rect 23753 33269 23765 33272
rect 23799 33269 23811 33303
rect 24228 33300 24256 33340
rect 24486 33328 24492 33380
rect 24544 33368 24550 33380
rect 25038 33368 25044 33380
rect 24544 33340 25044 33368
rect 24544 33328 24550 33340
rect 25038 33328 25044 33340
rect 25096 33328 25102 33380
rect 25516 33368 25544 33467
rect 26510 33464 26516 33516
rect 26568 33504 26574 33516
rect 28169 33507 28227 33513
rect 26568 33476 28120 33504
rect 26568 33464 26574 33476
rect 26605 33439 26663 33445
rect 26605 33405 26617 33439
rect 26651 33436 26663 33439
rect 27706 33436 27712 33448
rect 26651 33408 27712 33436
rect 26651 33405 26663 33408
rect 26605 33399 26663 33405
rect 27706 33396 27712 33408
rect 27764 33436 27770 33448
rect 27801 33439 27859 33445
rect 27801 33436 27813 33439
rect 27764 33408 27813 33436
rect 27764 33396 27770 33408
rect 27801 33405 27813 33408
rect 27847 33405 27859 33439
rect 27801 33399 27859 33405
rect 27893 33439 27951 33445
rect 27893 33405 27905 33439
rect 27939 33436 27951 33439
rect 27982 33436 27988 33448
rect 27939 33408 27988 33436
rect 27939 33405 27951 33408
rect 27893 33399 27951 33405
rect 27982 33396 27988 33408
rect 28040 33396 28046 33448
rect 28092 33436 28120 33476
rect 28169 33473 28181 33507
rect 28215 33504 28227 33507
rect 28902 33504 28908 33516
rect 28215 33476 28908 33504
rect 28215 33473 28227 33476
rect 28169 33467 28227 33473
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 29638 33513 29644 33516
rect 29636 33504 29644 33513
rect 29599 33476 29644 33504
rect 29636 33467 29644 33476
rect 29638 33464 29644 33467
rect 29696 33464 29702 33516
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 30006 33504 30012 33516
rect 29967 33476 30012 33504
rect 29825 33467 29883 33473
rect 28258 33436 28264 33448
rect 28092 33408 28264 33436
rect 28258 33396 28264 33408
rect 28316 33436 28322 33448
rect 29730 33436 29736 33448
rect 28316 33408 29736 33436
rect 28316 33396 28322 33408
rect 29730 33396 29736 33408
rect 29788 33396 29794 33448
rect 29840 33436 29868 33467
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 30098 33464 30104 33516
rect 30156 33464 30162 33516
rect 30282 33464 30288 33516
rect 30340 33504 30346 33516
rect 30837 33507 30895 33513
rect 30837 33504 30849 33507
rect 30340 33476 30849 33504
rect 30340 33464 30346 33476
rect 30837 33473 30849 33476
rect 30883 33473 30895 33507
rect 31573 33507 31631 33513
rect 30837 33467 30895 33473
rect 30944 33502 31524 33504
rect 31573 33502 31585 33507
rect 30944 33476 31585 33502
rect 30300 33436 30328 33464
rect 29840 33408 30328 33436
rect 30944 33368 30972 33476
rect 31496 33474 31585 33476
rect 31573 33473 31585 33474
rect 31619 33473 31631 33507
rect 32692 33504 32720 33544
rect 37461 33541 37473 33544
rect 37507 33541 37519 33575
rect 37461 33535 37519 33541
rect 37642 33532 37648 33584
rect 37700 33572 37706 33584
rect 38562 33572 38568 33584
rect 37700 33544 38568 33572
rect 37700 33532 37706 33544
rect 38562 33532 38568 33544
rect 38620 33572 38626 33584
rect 41046 33572 41052 33584
rect 38620 33544 41052 33572
rect 38620 33532 38626 33544
rect 41046 33532 41052 33544
rect 41104 33532 41110 33584
rect 42978 33572 42984 33584
rect 42076 33544 42984 33572
rect 31573 33467 31631 33473
rect 31680 33476 32720 33504
rect 31202 33396 31208 33448
rect 31260 33436 31266 33448
rect 31680 33436 31708 33476
rect 32766 33464 32772 33516
rect 32824 33464 32830 33516
rect 33229 33507 33287 33513
rect 33229 33473 33241 33507
rect 33275 33504 33287 33507
rect 33870 33504 33876 33516
rect 33275 33476 33876 33504
rect 33275 33473 33287 33476
rect 33229 33467 33287 33473
rect 33870 33464 33876 33476
rect 33928 33464 33934 33516
rect 34054 33464 34060 33516
rect 34112 33464 34118 33516
rect 34517 33507 34575 33513
rect 34517 33473 34529 33507
rect 34563 33504 34575 33507
rect 34698 33504 34704 33516
rect 34563 33476 34704 33504
rect 34563 33473 34575 33476
rect 34517 33467 34575 33473
rect 31260 33408 31708 33436
rect 31260 33396 31266 33408
rect 32582 33396 32588 33448
rect 32640 33436 32646 33448
rect 32677 33439 32735 33445
rect 32677 33436 32689 33439
rect 32640 33408 32689 33436
rect 32640 33396 32646 33408
rect 32677 33405 32689 33408
rect 32723 33436 32735 33439
rect 32858 33436 32864 33448
rect 32723 33408 32864 33436
rect 32723 33405 32735 33408
rect 32677 33399 32735 33405
rect 32858 33396 32864 33408
rect 32916 33396 32922 33448
rect 33594 33396 33600 33448
rect 33652 33436 33658 33448
rect 34532 33436 34560 33467
rect 34698 33464 34704 33476
rect 34756 33464 34762 33516
rect 35345 33507 35403 33513
rect 35345 33473 35357 33507
rect 35391 33473 35403 33507
rect 35989 33507 36047 33513
rect 35989 33504 36001 33507
rect 35345 33467 35403 33473
rect 35728 33476 36001 33504
rect 33652 33408 34560 33436
rect 33652 33396 33658 33408
rect 35250 33396 35256 33448
rect 35308 33396 35314 33448
rect 31018 33368 31024 33380
rect 25516 33340 31024 33368
rect 31018 33328 31024 33340
rect 31076 33328 31082 33380
rect 31665 33371 31723 33377
rect 31665 33337 31677 33371
rect 31711 33368 31723 33371
rect 35360 33368 35388 33467
rect 31711 33340 35388 33368
rect 31711 33337 31723 33340
rect 31665 33331 31723 33337
rect 25406 33300 25412 33312
rect 24228 33272 25412 33300
rect 23753 33263 23811 33269
rect 25406 33260 25412 33272
rect 25464 33300 25470 33312
rect 25961 33303 26019 33309
rect 25961 33300 25973 33303
rect 25464 33272 25973 33300
rect 25464 33260 25470 33272
rect 25961 33269 25973 33272
rect 26007 33300 26019 33303
rect 26326 33300 26332 33312
rect 26007 33272 26332 33300
rect 26007 33269 26019 33272
rect 25961 33263 26019 33269
rect 26326 33260 26332 33272
rect 26384 33260 26390 33312
rect 27249 33303 27307 33309
rect 27249 33269 27261 33303
rect 27295 33300 27307 33303
rect 27338 33300 27344 33312
rect 27295 33272 27344 33300
rect 27295 33269 27307 33272
rect 27249 33263 27307 33269
rect 27338 33260 27344 33272
rect 27396 33260 27402 33312
rect 27706 33260 27712 33312
rect 27764 33300 27770 33312
rect 28534 33300 28540 33312
rect 27764 33272 28540 33300
rect 27764 33260 27770 33272
rect 28534 33260 28540 33272
rect 28592 33260 28598 33312
rect 28994 33260 29000 33312
rect 29052 33260 29058 33312
rect 29454 33260 29460 33312
rect 29512 33260 29518 33312
rect 29730 33260 29736 33312
rect 29788 33300 29794 33312
rect 30926 33300 30932 33312
rect 29788 33272 30932 33300
rect 29788 33260 29794 33272
rect 30926 33260 30932 33272
rect 30984 33260 30990 33312
rect 31110 33260 31116 33312
rect 31168 33260 31174 33312
rect 31478 33260 31484 33312
rect 31536 33300 31542 33312
rect 32674 33300 32680 33312
rect 31536 33272 32680 33300
rect 31536 33260 31542 33272
rect 32674 33260 32680 33272
rect 32732 33260 32738 33312
rect 32769 33303 32827 33309
rect 32769 33269 32781 33303
rect 32815 33300 32827 33303
rect 32950 33300 32956 33312
rect 32815 33272 32956 33300
rect 32815 33269 32827 33272
rect 32769 33263 32827 33269
rect 32950 33260 32956 33272
rect 33008 33260 33014 33312
rect 33134 33260 33140 33312
rect 33192 33300 33198 33312
rect 33413 33303 33471 33309
rect 33413 33300 33425 33303
rect 33192 33272 33425 33300
rect 33192 33260 33198 33272
rect 33413 33269 33425 33272
rect 33459 33269 33471 33303
rect 33413 33263 33471 33269
rect 33962 33260 33968 33312
rect 34020 33300 34026 33312
rect 35728 33300 35756 33476
rect 35989 33473 36001 33476
rect 36035 33473 36047 33507
rect 35989 33467 36047 33473
rect 36630 33464 36636 33516
rect 36688 33504 36694 33516
rect 36725 33507 36783 33513
rect 36725 33504 36737 33507
rect 36688 33476 36737 33504
rect 36688 33464 36694 33476
rect 36725 33473 36737 33476
rect 36771 33473 36783 33507
rect 36725 33467 36783 33473
rect 36909 33507 36967 33513
rect 36909 33473 36921 33507
rect 36955 33504 36967 33507
rect 36998 33504 37004 33516
rect 36955 33476 37004 33504
rect 36955 33473 36967 33476
rect 36909 33467 36967 33473
rect 36998 33464 37004 33476
rect 37056 33464 37062 33516
rect 37550 33464 37556 33516
rect 37608 33504 37614 33516
rect 38197 33507 38255 33513
rect 38197 33504 38209 33507
rect 37608 33476 38209 33504
rect 37608 33464 37614 33476
rect 38197 33473 38209 33476
rect 38243 33473 38255 33507
rect 38197 33467 38255 33473
rect 38286 33464 38292 33516
rect 38344 33504 38350 33516
rect 38657 33507 38715 33513
rect 38657 33504 38669 33507
rect 38344 33476 38669 33504
rect 38344 33464 38350 33476
rect 38657 33473 38669 33476
rect 38703 33473 38715 33507
rect 38657 33467 38715 33473
rect 38764 33476 39068 33504
rect 35894 33396 35900 33448
rect 35952 33436 35958 33448
rect 36541 33439 36599 33445
rect 36541 33436 36553 33439
rect 35952 33408 36553 33436
rect 35952 33396 35958 33408
rect 36541 33405 36553 33408
rect 36587 33405 36599 33439
rect 36541 33399 36599 33405
rect 37829 33439 37887 33445
rect 37829 33405 37841 33439
rect 37875 33436 37887 33439
rect 38764 33436 38792 33476
rect 37875 33408 38792 33436
rect 38933 33439 38991 33445
rect 37875 33405 37887 33408
rect 37829 33399 37887 33405
rect 38933 33405 38945 33439
rect 38979 33405 38991 33439
rect 39040 33436 39068 33476
rect 39390 33464 39396 33516
rect 39448 33504 39454 33516
rect 39942 33504 39948 33516
rect 39448 33476 39948 33504
rect 39448 33464 39454 33476
rect 39942 33464 39948 33476
rect 40000 33464 40006 33516
rect 40037 33507 40095 33513
rect 40037 33473 40049 33507
rect 40083 33504 40095 33507
rect 40770 33504 40776 33516
rect 40083 33476 40776 33504
rect 40083 33473 40095 33476
rect 40037 33467 40095 33473
rect 40770 33464 40776 33476
rect 40828 33464 40834 33516
rect 40862 33464 40868 33516
rect 40920 33464 40926 33516
rect 41414 33464 41420 33516
rect 41472 33504 41478 33516
rect 42076 33513 42104 33544
rect 42978 33532 42984 33544
rect 43036 33532 43042 33584
rect 41693 33507 41751 33513
rect 41693 33504 41705 33507
rect 41472 33476 41705 33504
rect 41472 33464 41478 33476
rect 41693 33473 41705 33476
rect 41739 33473 41751 33507
rect 41693 33467 41751 33473
rect 42061 33507 42119 33513
rect 42061 33473 42073 33507
rect 42107 33473 42119 33507
rect 42061 33467 42119 33473
rect 42794 33464 42800 33516
rect 42852 33464 42858 33516
rect 39482 33436 39488 33448
rect 39040 33408 39488 33436
rect 38933 33399 38991 33405
rect 35805 33371 35863 33377
rect 35805 33337 35817 33371
rect 35851 33368 35863 33371
rect 36078 33368 36084 33380
rect 35851 33340 36084 33368
rect 35851 33337 35863 33340
rect 35805 33331 35863 33337
rect 36078 33328 36084 33340
rect 36136 33368 36142 33380
rect 37458 33368 37464 33380
rect 36136 33340 37464 33368
rect 36136 33328 36142 33340
rect 37458 33328 37464 33340
rect 37516 33328 37522 33380
rect 37734 33328 37740 33380
rect 37792 33368 37798 33380
rect 37921 33371 37979 33377
rect 37921 33368 37933 33371
rect 37792 33340 37933 33368
rect 37792 33328 37798 33340
rect 37921 33337 37933 33340
rect 37967 33337 37979 33371
rect 38948 33368 38976 33399
rect 39482 33396 39488 33408
rect 39540 33396 39546 33448
rect 41049 33371 41107 33377
rect 38948 33340 40172 33368
rect 37921 33331 37979 33337
rect 37642 33300 37648 33312
rect 34020 33272 37648 33300
rect 34020 33260 34026 33272
rect 37642 33260 37648 33272
rect 37700 33260 37706 33312
rect 38059 33303 38117 33309
rect 38059 33269 38071 33303
rect 38105 33300 38117 33303
rect 38470 33300 38476 33312
rect 38105 33272 38476 33300
rect 38105 33269 38117 33272
rect 38059 33263 38117 33269
rect 38470 33260 38476 33272
rect 38528 33260 38534 33312
rect 38746 33260 38752 33312
rect 38804 33300 38810 33312
rect 39022 33300 39028 33312
rect 38804 33272 39028 33300
rect 38804 33260 38810 33272
rect 39022 33260 39028 33272
rect 39080 33260 39086 33312
rect 40144 33300 40172 33340
rect 41049 33337 41061 33371
rect 41095 33368 41107 33371
rect 41598 33368 41604 33380
rect 41095 33340 41604 33368
rect 41095 33337 41107 33340
rect 41049 33331 41107 33337
rect 41598 33328 41604 33340
rect 41656 33328 41662 33380
rect 41509 33303 41567 33309
rect 41509 33300 41521 33303
rect 40144 33272 41521 33300
rect 41509 33269 41521 33272
rect 41555 33269 41567 33303
rect 41509 33263 41567 33269
rect 41874 33260 41880 33312
rect 41932 33260 41938 33312
rect 42426 33260 42432 33312
rect 42484 33300 42490 33312
rect 42705 33303 42763 33309
rect 42705 33300 42717 33303
rect 42484 33272 42717 33300
rect 42484 33260 42490 33272
rect 42705 33269 42717 33272
rect 42751 33269 42763 33303
rect 42705 33263 42763 33269
rect 1104 33210 43884 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 43884 33210
rect 1104 33136 43884 33158
rect 12618 33056 12624 33108
rect 12676 33056 12682 33108
rect 13081 33099 13139 33105
rect 13081 33065 13093 33099
rect 13127 33096 13139 33099
rect 13262 33096 13268 33108
rect 13127 33068 13268 33096
rect 13127 33065 13139 33068
rect 13081 33059 13139 33065
rect 13096 32960 13124 33059
rect 13262 33056 13268 33068
rect 13320 33056 13326 33108
rect 14366 33056 14372 33108
rect 14424 33056 14430 33108
rect 16482 33056 16488 33108
rect 16540 33056 16546 33108
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 16761 33099 16819 33105
rect 16761 33096 16773 33099
rect 16724 33068 16773 33096
rect 16724 33056 16730 33068
rect 16761 33065 16773 33068
rect 16807 33065 16819 33099
rect 16761 33059 16819 33065
rect 17865 33099 17923 33105
rect 17865 33065 17877 33099
rect 17911 33096 17923 33099
rect 18046 33096 18052 33108
rect 17911 33068 18052 33096
rect 17911 33065 17923 33068
rect 17865 33059 17923 33065
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 18322 33056 18328 33108
rect 18380 33096 18386 33108
rect 19889 33099 19947 33105
rect 18380 33068 18828 33096
rect 18380 33056 18386 33068
rect 18690 32988 18696 33040
rect 18748 32988 18754 33040
rect 18800 33028 18828 33068
rect 19889 33065 19901 33099
rect 19935 33096 19947 33099
rect 20254 33096 20260 33108
rect 19935 33068 20260 33096
rect 19935 33065 19947 33068
rect 19889 33059 19947 33065
rect 20254 33056 20260 33068
rect 20312 33056 20318 33108
rect 23477 33099 23535 33105
rect 23477 33096 23489 33099
rect 20732 33068 23489 33096
rect 20732 33028 20760 33068
rect 23477 33065 23489 33068
rect 23523 33065 23535 33099
rect 23477 33059 23535 33065
rect 23845 33099 23903 33105
rect 23845 33065 23857 33099
rect 23891 33096 23903 33099
rect 24118 33096 24124 33108
rect 23891 33068 24124 33096
rect 23891 33065 23903 33068
rect 23845 33059 23903 33065
rect 24118 33056 24124 33068
rect 24176 33096 24182 33108
rect 24302 33096 24308 33108
rect 24176 33068 24308 33096
rect 24176 33056 24182 33068
rect 24302 33056 24308 33068
rect 24360 33056 24366 33108
rect 25222 33056 25228 33108
rect 25280 33096 25286 33108
rect 25869 33099 25927 33105
rect 25869 33096 25881 33099
rect 25280 33068 25881 33096
rect 25280 33056 25286 33068
rect 25869 33065 25881 33068
rect 25915 33065 25927 33099
rect 25869 33059 25927 33065
rect 27062 33056 27068 33108
rect 27120 33056 27126 33108
rect 28810 33056 28816 33108
rect 28868 33056 28874 33108
rect 30374 33056 30380 33108
rect 30432 33096 30438 33108
rect 30745 33099 30803 33105
rect 30745 33096 30757 33099
rect 30432 33068 30757 33096
rect 30432 33056 30438 33068
rect 30745 33065 30757 33068
rect 30791 33065 30803 33099
rect 30745 33059 30803 33065
rect 30926 33056 30932 33108
rect 30984 33096 30990 33108
rect 34330 33096 34336 33108
rect 30984 33068 34336 33096
rect 30984 33056 30990 33068
rect 34330 33056 34336 33068
rect 34388 33056 34394 33108
rect 35710 33056 35716 33108
rect 35768 33096 35774 33108
rect 36541 33099 36599 33105
rect 36541 33096 36553 33099
rect 35768 33068 36553 33096
rect 35768 33056 35774 33068
rect 36541 33065 36553 33068
rect 36587 33065 36599 33099
rect 36541 33059 36599 33065
rect 36725 33099 36783 33105
rect 36725 33065 36737 33099
rect 36771 33065 36783 33099
rect 36725 33059 36783 33065
rect 21085 33031 21143 33037
rect 21085 33028 21097 33031
rect 18800 33000 20760 33028
rect 20824 33000 21097 33028
rect 12452 32932 13124 32960
rect 15841 32963 15899 32969
rect 12452 32901 12480 32932
rect 15841 32929 15853 32963
rect 15887 32960 15899 32963
rect 16206 32960 16212 32972
rect 15887 32932 16212 32960
rect 15887 32929 15899 32932
rect 15841 32923 15899 32929
rect 16206 32920 16212 32932
rect 16264 32920 16270 32972
rect 16298 32920 16304 32972
rect 16356 32960 16362 32972
rect 16485 32963 16543 32969
rect 16485 32960 16497 32963
rect 16356 32932 16497 32960
rect 16356 32920 16362 32932
rect 16485 32929 16497 32932
rect 16531 32929 16543 32963
rect 16485 32923 16543 32929
rect 18417 32963 18475 32969
rect 18417 32929 18429 32963
rect 18463 32960 18475 32963
rect 19610 32960 19616 32972
rect 18463 32932 19616 32960
rect 18463 32929 18475 32932
rect 18417 32923 18475 32929
rect 19610 32920 19616 32932
rect 19668 32920 19674 32972
rect 20438 32920 20444 32972
rect 20496 32920 20502 32972
rect 12437 32895 12495 32901
rect 12437 32861 12449 32895
rect 12483 32861 12495 32895
rect 12437 32855 12495 32861
rect 12618 32852 12624 32904
rect 12676 32852 12682 32904
rect 13354 32852 13360 32904
rect 13412 32852 13418 32904
rect 13906 32852 13912 32904
rect 13964 32892 13970 32904
rect 14737 32895 14795 32901
rect 13964 32864 14688 32892
rect 13964 32852 13970 32864
rect 13078 32784 13084 32836
rect 13136 32784 13142 32836
rect 14550 32784 14556 32836
rect 14608 32784 14614 32836
rect 14660 32824 14688 32864
rect 14737 32861 14749 32895
rect 14783 32892 14795 32895
rect 16316 32892 16344 32920
rect 14783 32864 16344 32892
rect 14783 32861 14795 32864
rect 14737 32855 14795 32861
rect 16390 32852 16396 32904
rect 16448 32852 16454 32904
rect 17218 32852 17224 32904
rect 17276 32892 17282 32904
rect 17497 32895 17555 32901
rect 17497 32892 17509 32895
rect 17276 32864 17509 32892
rect 17276 32852 17282 32864
rect 17497 32861 17509 32864
rect 17543 32861 17555 32895
rect 17497 32855 17555 32861
rect 20257 32895 20315 32901
rect 20257 32861 20269 32895
rect 20303 32892 20315 32895
rect 20714 32892 20720 32904
rect 20303 32864 20720 32892
rect 20303 32861 20315 32864
rect 20257 32855 20315 32861
rect 20714 32852 20720 32864
rect 20772 32852 20778 32904
rect 14660 32796 16068 32824
rect 13262 32716 13268 32768
rect 13320 32716 13326 32768
rect 14090 32716 14096 32768
rect 14148 32756 14154 32768
rect 15197 32759 15255 32765
rect 15197 32756 15209 32759
rect 14148 32728 15209 32756
rect 14148 32716 14154 32728
rect 15197 32725 15209 32728
rect 15243 32725 15255 32759
rect 15197 32719 15255 32725
rect 15378 32716 15384 32768
rect 15436 32756 15442 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 15436 32728 15577 32756
rect 15436 32716 15442 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 15565 32719 15623 32725
rect 15657 32759 15715 32765
rect 15657 32725 15669 32759
rect 15703 32756 15715 32759
rect 15930 32756 15936 32768
rect 15703 32728 15936 32756
rect 15703 32725 15715 32728
rect 15657 32719 15715 32725
rect 15930 32716 15936 32728
rect 15988 32716 15994 32768
rect 16040 32756 16068 32796
rect 17678 32784 17684 32836
rect 17736 32784 17742 32836
rect 20824 32824 20852 33000
rect 21085 32997 21097 33000
rect 21131 32997 21143 33031
rect 21085 32991 21143 32997
rect 21910 32988 21916 33040
rect 21968 33028 21974 33040
rect 29733 33031 29791 33037
rect 29733 33028 29745 33031
rect 21968 33000 29745 33028
rect 21968 32988 21974 33000
rect 29733 32997 29745 33000
rect 29779 32997 29791 33031
rect 29733 32991 29791 32997
rect 29914 32988 29920 33040
rect 29972 32988 29978 33040
rect 31754 32988 31760 33040
rect 31812 32988 31818 33040
rect 32950 32988 32956 33040
rect 33008 32988 33014 33040
rect 34149 33031 34207 33037
rect 34149 32997 34161 33031
rect 34195 33028 34207 33031
rect 34606 33028 34612 33040
rect 34195 33000 34612 33028
rect 34195 32997 34207 33000
rect 34149 32991 34207 32997
rect 34606 32988 34612 33000
rect 34664 32988 34670 33040
rect 35894 32988 35900 33040
rect 35952 33028 35958 33040
rect 36740 33028 36768 33059
rect 36814 33056 36820 33108
rect 36872 33096 36878 33108
rect 37369 33099 37427 33105
rect 37369 33096 37381 33099
rect 36872 33068 37381 33096
rect 36872 33056 36878 33068
rect 37369 33065 37381 33068
rect 37415 33096 37427 33099
rect 37642 33096 37648 33108
rect 37415 33068 37648 33096
rect 37415 33065 37427 33068
rect 37369 33059 37427 33065
rect 37642 33056 37648 33068
rect 37700 33056 37706 33108
rect 37734 33056 37740 33108
rect 37792 33056 37798 33108
rect 40954 33028 40960 33040
rect 35952 33000 40960 33028
rect 35952 32988 35958 33000
rect 40954 32988 40960 33000
rect 41012 32988 41018 33040
rect 21266 32920 21272 32972
rect 21324 32960 21330 32972
rect 21634 32960 21640 32972
rect 21324 32932 21640 32960
rect 21324 32920 21330 32932
rect 21634 32920 21640 32932
rect 21692 32920 21698 32972
rect 23750 32920 23756 32972
rect 23808 32960 23814 32972
rect 23937 32963 23995 32969
rect 23937 32960 23949 32963
rect 23808 32932 23949 32960
rect 23808 32920 23814 32932
rect 23937 32929 23949 32932
rect 23983 32929 23995 32963
rect 25130 32960 25136 32972
rect 23937 32923 23995 32929
rect 25056 32932 25136 32960
rect 22094 32852 22100 32904
rect 22152 32892 22158 32904
rect 22462 32892 22468 32904
rect 22152 32864 22468 32892
rect 22152 32852 22158 32864
rect 22462 32852 22468 32864
rect 22520 32852 22526 32904
rect 22554 32852 22560 32904
rect 22612 32852 22618 32904
rect 22646 32852 22652 32904
rect 22704 32852 22710 32904
rect 22830 32852 22836 32904
rect 22888 32852 22894 32904
rect 23661 32895 23719 32901
rect 23661 32861 23673 32895
rect 23707 32892 23719 32895
rect 23842 32892 23848 32904
rect 23707 32864 23848 32892
rect 23707 32861 23719 32864
rect 23661 32855 23719 32861
rect 23842 32852 23848 32864
rect 23900 32852 23906 32904
rect 25056 32901 25084 32932
rect 25130 32920 25136 32932
rect 25188 32960 25194 32972
rect 26142 32960 26148 32972
rect 25188 32932 26148 32960
rect 25188 32920 25194 32932
rect 26142 32920 26148 32932
rect 26200 32960 26206 32972
rect 27617 32963 27675 32969
rect 26200 32932 26924 32960
rect 26200 32920 26206 32932
rect 25041 32895 25099 32901
rect 25041 32861 25053 32895
rect 25087 32861 25099 32895
rect 25041 32855 25099 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32892 25467 32895
rect 25682 32892 25688 32904
rect 25455 32864 25688 32892
rect 25455 32861 25467 32864
rect 25409 32855 25467 32861
rect 25682 32852 25688 32864
rect 25740 32852 25746 32904
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26896 32901 26924 32932
rect 27617 32929 27629 32963
rect 27663 32960 27675 32963
rect 27798 32960 27804 32972
rect 27663 32932 27804 32960
rect 27663 32929 27675 32932
rect 27617 32923 27675 32929
rect 27798 32920 27804 32932
rect 27856 32920 27862 32972
rect 27982 32920 27988 32972
rect 28040 32960 28046 32972
rect 28534 32960 28540 32972
rect 28040 32932 28540 32960
rect 28040 32920 28046 32932
rect 28534 32920 28540 32932
rect 28592 32920 28598 32972
rect 29932 32960 29960 32988
rect 34057 32963 34115 32969
rect 28966 32932 29960 32960
rect 30024 32932 31984 32960
rect 26513 32895 26571 32901
rect 26513 32892 26525 32895
rect 26384 32864 26525 32892
rect 26384 32852 26390 32864
rect 26513 32861 26525 32864
rect 26559 32861 26571 32895
rect 26513 32855 26571 32861
rect 26881 32895 26939 32901
rect 26881 32861 26893 32895
rect 26927 32892 26939 32895
rect 26927 32864 27568 32892
rect 26927 32861 26939 32864
rect 26881 32855 26939 32861
rect 17788 32796 20852 32824
rect 17788 32756 17816 32796
rect 20898 32784 20904 32836
rect 20956 32824 20962 32836
rect 21453 32827 21511 32833
rect 21453 32824 21465 32827
rect 20956 32796 21465 32824
rect 20956 32784 20962 32796
rect 21453 32793 21465 32796
rect 21499 32824 21511 32827
rect 21726 32824 21732 32836
rect 21499 32796 21732 32824
rect 21499 32793 21511 32796
rect 21453 32787 21511 32793
rect 21726 32784 21732 32796
rect 21784 32784 21790 32836
rect 25133 32827 25191 32833
rect 25133 32824 25145 32827
rect 25056 32796 25145 32824
rect 25056 32768 25084 32796
rect 25133 32793 25145 32796
rect 25179 32793 25191 32827
rect 25133 32787 25191 32793
rect 25225 32827 25283 32833
rect 25225 32793 25237 32827
rect 25271 32824 25283 32827
rect 25314 32824 25320 32836
rect 25271 32796 25320 32824
rect 25271 32793 25283 32796
rect 25225 32787 25283 32793
rect 25314 32784 25320 32796
rect 25372 32824 25378 32836
rect 26697 32827 26755 32833
rect 26697 32824 26709 32827
rect 25372 32796 26709 32824
rect 25372 32784 25378 32796
rect 26697 32793 26709 32796
rect 26743 32793 26755 32827
rect 26697 32787 26755 32793
rect 16040 32728 17816 32756
rect 18877 32759 18935 32765
rect 18877 32725 18889 32759
rect 18923 32756 18935 32759
rect 19978 32756 19984 32768
rect 18923 32728 19984 32756
rect 18923 32725 18935 32728
rect 18877 32719 18935 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20346 32716 20352 32768
rect 20404 32716 20410 32768
rect 21545 32759 21603 32765
rect 21545 32725 21557 32759
rect 21591 32756 21603 32759
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 21591 32728 22293 32756
rect 21591 32725 21603 32728
rect 21545 32719 21603 32725
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 22281 32719 22339 32725
rect 22370 32716 22376 32768
rect 22428 32756 22434 32768
rect 24857 32759 24915 32765
rect 24857 32756 24869 32759
rect 22428 32728 24869 32756
rect 22428 32716 22434 32728
rect 24857 32725 24869 32728
rect 24903 32725 24915 32759
rect 24857 32719 24915 32725
rect 25038 32716 25044 32768
rect 25096 32716 25102 32768
rect 26712 32756 26740 32787
rect 26786 32784 26792 32836
rect 26844 32784 26850 32836
rect 27430 32756 27436 32768
rect 26712 32728 27436 32756
rect 27430 32716 27436 32728
rect 27488 32716 27494 32768
rect 27540 32756 27568 32864
rect 27706 32852 27712 32904
rect 27764 32852 27770 32904
rect 27893 32895 27951 32901
rect 27893 32861 27905 32895
rect 27939 32892 27951 32895
rect 27939 32864 28672 32892
rect 27939 32861 27951 32864
rect 27893 32855 27951 32861
rect 27724 32824 27752 32852
rect 28644 32833 28672 32864
rect 28445 32827 28503 32833
rect 28445 32824 28457 32827
rect 27724 32796 28457 32824
rect 28445 32793 28457 32796
rect 28491 32793 28503 32827
rect 28445 32787 28503 32793
rect 28629 32827 28687 32833
rect 28629 32793 28641 32827
rect 28675 32824 28687 32827
rect 28810 32824 28816 32836
rect 28675 32796 28816 32824
rect 28675 32793 28687 32796
rect 28629 32787 28687 32793
rect 28810 32784 28816 32796
rect 28868 32784 28874 32836
rect 28966 32824 28994 32932
rect 29454 32852 29460 32904
rect 29512 32892 29518 32904
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 29512 32864 29745 32892
rect 29512 32852 29518 32864
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29914 32852 29920 32904
rect 29972 32892 29978 32904
rect 30024 32901 30052 32932
rect 31956 32904 31984 32932
rect 34057 32929 34069 32963
rect 34103 32960 34115 32963
rect 35342 32960 35348 32972
rect 34103 32932 35348 32960
rect 34103 32929 34115 32932
rect 34057 32923 34115 32929
rect 35342 32920 35348 32932
rect 35400 32920 35406 32972
rect 35618 32920 35624 32972
rect 35676 32920 35682 32972
rect 35986 32920 35992 32972
rect 36044 32960 36050 32972
rect 37461 32963 37519 32969
rect 37461 32960 37473 32963
rect 36044 32932 37473 32960
rect 36044 32920 36050 32932
rect 37461 32929 37473 32932
rect 37507 32929 37519 32963
rect 37461 32923 37519 32929
rect 37642 32920 37648 32972
rect 37700 32960 37706 32972
rect 41046 32960 41052 32972
rect 37700 32932 41052 32960
rect 37700 32920 37706 32932
rect 41046 32920 41052 32932
rect 41104 32920 41110 32972
rect 41322 32920 41328 32972
rect 41380 32920 41386 32972
rect 41598 32920 41604 32972
rect 41656 32920 41662 32972
rect 42794 32920 42800 32972
rect 42852 32960 42858 32972
rect 43349 32963 43407 32969
rect 43349 32960 43361 32963
rect 42852 32932 43361 32960
rect 42852 32920 42858 32932
rect 43349 32929 43361 32932
rect 43395 32929 43407 32963
rect 43349 32923 43407 32929
rect 30009 32895 30067 32901
rect 30009 32892 30021 32895
rect 29972 32864 30021 32892
rect 29972 32852 29978 32864
rect 30009 32861 30021 32864
rect 30055 32861 30067 32895
rect 30282 32892 30288 32904
rect 30009 32855 30067 32861
rect 30116 32864 30288 32892
rect 28920 32796 28994 32824
rect 28920 32756 28948 32796
rect 29270 32784 29276 32836
rect 29328 32824 29334 32836
rect 30116 32824 30144 32864
rect 30282 32852 30288 32864
rect 30340 32892 30346 32904
rect 30469 32895 30527 32901
rect 30469 32892 30481 32895
rect 30340 32864 30481 32892
rect 30340 32852 30346 32864
rect 30469 32861 30481 32864
rect 30515 32861 30527 32895
rect 30469 32855 30527 32861
rect 30558 32852 30564 32904
rect 30616 32852 30622 32904
rect 30742 32852 30748 32904
rect 30800 32852 30806 32904
rect 31938 32852 31944 32904
rect 31996 32852 32002 32904
rect 32030 32852 32036 32904
rect 32088 32892 32094 32904
rect 32214 32892 32220 32904
rect 32088 32864 32220 32892
rect 32088 32852 32094 32864
rect 32214 32852 32220 32864
rect 32272 32852 32278 32904
rect 32306 32852 32312 32904
rect 32364 32852 32370 32904
rect 32674 32852 32680 32904
rect 32732 32892 32738 32904
rect 32769 32895 32827 32901
rect 32769 32892 32781 32895
rect 32732 32864 32781 32892
rect 32732 32852 32738 32864
rect 32769 32861 32781 32864
rect 32815 32861 32827 32895
rect 32769 32855 32827 32861
rect 33962 32852 33968 32904
rect 34020 32852 34026 32904
rect 34241 32895 34299 32901
rect 34241 32861 34253 32895
rect 34287 32861 34299 32895
rect 34241 32855 34299 32861
rect 35529 32895 35587 32901
rect 35529 32861 35541 32895
rect 35575 32892 35587 32895
rect 35802 32892 35808 32904
rect 35575 32864 35808 32892
rect 35575 32861 35587 32864
rect 35529 32855 35587 32861
rect 29328 32796 30144 32824
rect 29328 32784 29334 32796
rect 30190 32784 30196 32836
rect 30248 32824 30254 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 30248 32796 32137 32824
rect 30248 32784 30254 32796
rect 32125 32793 32137 32796
rect 32171 32824 32183 32827
rect 32398 32824 32404 32836
rect 32171 32796 32404 32824
rect 32171 32793 32183 32796
rect 32125 32787 32183 32793
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 33778 32784 33784 32836
rect 33836 32784 33842 32836
rect 34256 32824 34284 32855
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 36078 32852 36084 32904
rect 36136 32852 36142 32904
rect 37366 32852 37372 32904
rect 37424 32852 37430 32904
rect 39209 32895 39267 32901
rect 39209 32861 39221 32895
rect 39255 32861 39267 32895
rect 39209 32855 39267 32861
rect 36909 32827 36967 32833
rect 36909 32824 36921 32827
rect 33980 32796 34284 32824
rect 34992 32796 36921 32824
rect 33980 32768 34008 32796
rect 27540 32728 28948 32756
rect 28994 32716 29000 32768
rect 29052 32756 29058 32768
rect 29917 32759 29975 32765
rect 29917 32756 29929 32759
rect 29052 32728 29929 32756
rect 29052 32716 29058 32728
rect 29917 32725 29929 32728
rect 29963 32725 29975 32759
rect 29917 32719 29975 32725
rect 31202 32716 31208 32768
rect 31260 32716 31266 32768
rect 33962 32716 33968 32768
rect 34020 32716 34026 32768
rect 34054 32716 34060 32768
rect 34112 32756 34118 32768
rect 34992 32756 35020 32796
rect 36909 32793 36921 32796
rect 36955 32793 36967 32827
rect 39224 32824 39252 32855
rect 39390 32852 39396 32904
rect 39448 32852 39454 32904
rect 40034 32852 40040 32904
rect 40092 32852 40098 32904
rect 40221 32895 40279 32901
rect 40221 32861 40233 32895
rect 40267 32861 40279 32895
rect 40221 32855 40279 32861
rect 40681 32895 40739 32901
rect 40681 32861 40693 32895
rect 40727 32892 40739 32895
rect 40770 32892 40776 32904
rect 40727 32864 40776 32892
rect 40727 32861 40739 32864
rect 40681 32855 40739 32861
rect 39942 32824 39948 32836
rect 39224 32796 39948 32824
rect 36909 32787 36967 32793
rect 39942 32784 39948 32796
rect 40000 32824 40006 32836
rect 40129 32827 40187 32833
rect 40129 32824 40141 32827
rect 40000 32796 40141 32824
rect 40000 32784 40006 32796
rect 40129 32793 40141 32796
rect 40175 32793 40187 32827
rect 40236 32824 40264 32855
rect 40770 32852 40776 32864
rect 40828 32852 40834 32904
rect 40862 32852 40868 32904
rect 40920 32852 40926 32904
rect 42702 32852 42708 32904
rect 42760 32852 42766 32904
rect 41138 32824 41144 32836
rect 40236 32796 41144 32824
rect 40129 32787 40187 32793
rect 34112 32728 35020 32756
rect 36709 32759 36767 32765
rect 34112 32716 34118 32728
rect 36709 32725 36721 32759
rect 36755 32756 36767 32759
rect 37642 32756 37648 32768
rect 36755 32728 37648 32756
rect 36755 32725 36767 32728
rect 36709 32719 36767 32725
rect 37642 32716 37648 32728
rect 37700 32716 37706 32768
rect 38194 32716 38200 32768
rect 38252 32716 38258 32768
rect 39298 32716 39304 32768
rect 39356 32716 39362 32768
rect 40144 32756 40172 32787
rect 41138 32784 41144 32796
rect 41196 32784 41202 32836
rect 40494 32756 40500 32768
rect 40144 32728 40500 32756
rect 40494 32716 40500 32728
rect 40552 32716 40558 32768
rect 40678 32716 40684 32768
rect 40736 32756 40742 32768
rect 40773 32759 40831 32765
rect 40773 32756 40785 32759
rect 40736 32728 40785 32756
rect 40736 32716 40742 32728
rect 40773 32725 40785 32728
rect 40819 32725 40831 32759
rect 40773 32719 40831 32725
rect 1104 32666 43884 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 43884 32666
rect 1104 32592 43884 32614
rect 15194 32512 15200 32564
rect 15252 32552 15258 32564
rect 15933 32555 15991 32561
rect 15933 32552 15945 32555
rect 15252 32524 15945 32552
rect 15252 32512 15258 32524
rect 15933 32521 15945 32524
rect 15979 32521 15991 32555
rect 15933 32515 15991 32521
rect 16301 32555 16359 32561
rect 16301 32521 16313 32555
rect 16347 32552 16359 32555
rect 16390 32552 16396 32564
rect 16347 32524 16396 32552
rect 16347 32521 16359 32524
rect 16301 32515 16359 32521
rect 16390 32512 16396 32524
rect 16448 32512 16454 32564
rect 18598 32552 18604 32564
rect 16500 32524 18604 32552
rect 13081 32487 13139 32493
rect 13081 32453 13093 32487
rect 13127 32484 13139 32487
rect 13170 32484 13176 32496
rect 13127 32456 13176 32484
rect 13127 32453 13139 32456
rect 13081 32447 13139 32453
rect 13170 32444 13176 32456
rect 13228 32484 13234 32496
rect 14274 32484 14280 32496
rect 13228 32456 14280 32484
rect 13228 32444 13234 32456
rect 14274 32444 14280 32456
rect 14332 32444 14338 32496
rect 16500 32484 16528 32524
rect 18598 32512 18604 32524
rect 18656 32512 18662 32564
rect 20162 32512 20168 32564
rect 20220 32512 20226 32564
rect 20809 32555 20867 32561
rect 20809 32521 20821 32555
rect 20855 32552 20867 32555
rect 20898 32552 20904 32564
rect 20855 32524 20904 32552
rect 20855 32521 20867 32524
rect 20809 32515 20867 32521
rect 20898 32512 20904 32524
rect 20956 32512 20962 32564
rect 21453 32555 21511 32561
rect 21453 32521 21465 32555
rect 21499 32552 21511 32555
rect 22094 32552 22100 32564
rect 21499 32524 22100 32552
rect 21499 32521 21511 32524
rect 21453 32515 21511 32521
rect 22094 32512 22100 32524
rect 22152 32512 22158 32564
rect 22189 32555 22247 32561
rect 22189 32521 22201 32555
rect 22235 32552 22247 32555
rect 22830 32552 22836 32564
rect 22235 32524 22836 32552
rect 22235 32521 22247 32524
rect 22189 32515 22247 32521
rect 22830 32512 22836 32524
rect 22888 32512 22894 32564
rect 24854 32552 24860 32564
rect 24044 32524 24860 32552
rect 15764 32456 16528 32484
rect 18049 32487 18107 32493
rect 13265 32419 13323 32425
rect 13265 32385 13277 32419
rect 13311 32416 13323 32419
rect 13725 32419 13783 32425
rect 13725 32416 13737 32419
rect 13311 32388 13737 32416
rect 13311 32385 13323 32388
rect 13265 32379 13323 32385
rect 13725 32385 13737 32388
rect 13771 32385 13783 32419
rect 13725 32379 13783 32385
rect 13906 32376 13912 32428
rect 13964 32376 13970 32428
rect 14090 32376 14096 32428
rect 14148 32376 14154 32428
rect 14185 32419 14243 32425
rect 14185 32385 14197 32419
rect 14231 32416 14243 32419
rect 14921 32419 14979 32425
rect 14921 32416 14933 32419
rect 14231 32388 14933 32416
rect 14231 32385 14243 32388
rect 14185 32379 14243 32385
rect 14921 32385 14933 32388
rect 14967 32416 14979 32419
rect 15010 32416 15016 32428
rect 14967 32388 15016 32416
rect 14967 32385 14979 32388
rect 14921 32379 14979 32385
rect 15010 32376 15016 32388
rect 15068 32376 15074 32428
rect 15105 32419 15163 32425
rect 15105 32385 15117 32419
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 13924 32280 13952 32376
rect 14458 32280 14464 32292
rect 13924 32252 14464 32280
rect 14458 32240 14464 32252
rect 14516 32240 14522 32292
rect 15120 32280 15148 32379
rect 15764 32357 15792 32456
rect 18049 32453 18061 32487
rect 18095 32484 18107 32487
rect 18693 32487 18751 32493
rect 18693 32484 18705 32487
rect 18095 32456 18705 32484
rect 18095 32453 18107 32456
rect 18049 32447 18107 32453
rect 18693 32453 18705 32456
rect 18739 32453 18751 32487
rect 24044 32484 24072 32524
rect 24854 32512 24860 32524
rect 24912 32512 24918 32564
rect 24946 32512 24952 32564
rect 25004 32552 25010 32564
rect 25777 32555 25835 32561
rect 25777 32552 25789 32555
rect 25004 32524 25789 32552
rect 25004 32512 25010 32524
rect 25777 32521 25789 32524
rect 25823 32521 25835 32555
rect 25777 32515 25835 32521
rect 26234 32512 26240 32564
rect 26292 32552 26298 32564
rect 27154 32552 27160 32564
rect 26292 32524 27160 32552
rect 26292 32512 26298 32524
rect 27154 32512 27160 32524
rect 27212 32512 27218 32564
rect 28994 32552 29000 32564
rect 28092 32524 29000 32552
rect 18693 32447 18751 32453
rect 21284 32456 22094 32484
rect 17770 32376 17776 32428
rect 17828 32376 17834 32428
rect 17862 32376 17868 32428
rect 17920 32376 17926 32428
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 18598 32416 18604 32428
rect 18380 32388 18604 32416
rect 18380 32376 18386 32388
rect 18598 32376 18604 32388
rect 18656 32376 18662 32428
rect 18966 32376 18972 32428
rect 19024 32376 19030 32428
rect 19058 32376 19064 32428
rect 19116 32376 19122 32428
rect 19150 32376 19156 32428
rect 19208 32376 19214 32428
rect 19334 32376 19340 32428
rect 19392 32376 19398 32428
rect 21284 32425 21312 32456
rect 21269 32419 21327 32425
rect 21269 32416 21281 32419
rect 19720 32388 21281 32416
rect 15749 32351 15807 32357
rect 15749 32317 15761 32351
rect 15795 32317 15807 32351
rect 15749 32311 15807 32317
rect 15841 32351 15899 32357
rect 15841 32317 15853 32351
rect 15887 32348 15899 32351
rect 15930 32348 15936 32360
rect 15887 32320 15936 32348
rect 15887 32317 15899 32320
rect 15841 32311 15899 32317
rect 15856 32280 15884 32311
rect 15930 32308 15936 32320
rect 15988 32308 15994 32360
rect 16206 32308 16212 32360
rect 16264 32348 16270 32360
rect 19720 32348 19748 32388
rect 21269 32385 21281 32388
rect 21315 32385 21327 32419
rect 21269 32379 21327 32385
rect 21453 32419 21511 32425
rect 21453 32385 21465 32419
rect 21499 32385 21511 32419
rect 22066 32416 22094 32456
rect 23952 32456 24072 32484
rect 24121 32487 24179 32493
rect 23952 32428 23980 32456
rect 24121 32453 24133 32487
rect 24167 32484 24179 32487
rect 24670 32484 24676 32496
rect 24167 32456 24676 32484
rect 24167 32453 24179 32456
rect 24121 32447 24179 32453
rect 24670 32444 24676 32456
rect 24728 32484 24734 32496
rect 25133 32487 25191 32493
rect 25133 32484 25145 32487
rect 24728 32456 25145 32484
rect 24728 32444 24734 32456
rect 25133 32453 25145 32456
rect 25179 32484 25191 32487
rect 26145 32487 26203 32493
rect 26145 32484 26157 32487
rect 25179 32456 26157 32484
rect 25179 32453 25191 32456
rect 25133 32447 25191 32453
rect 26145 32453 26157 32456
rect 26191 32453 26203 32487
rect 27246 32484 27252 32496
rect 26145 32447 26203 32453
rect 26252 32456 27252 32484
rect 22741 32419 22799 32425
rect 22741 32416 22753 32419
rect 22066 32388 22753 32416
rect 21453 32379 21511 32385
rect 22741 32385 22753 32388
rect 22787 32385 22799 32419
rect 22741 32379 22799 32385
rect 16264 32320 19748 32348
rect 20349 32351 20407 32357
rect 16264 32308 16270 32320
rect 20349 32317 20361 32351
rect 20395 32317 20407 32351
rect 20349 32311 20407 32317
rect 20441 32351 20499 32357
rect 20441 32317 20453 32351
rect 20487 32348 20499 32351
rect 20530 32348 20536 32360
rect 20487 32320 20536 32348
rect 20487 32317 20499 32320
rect 20441 32311 20499 32317
rect 15120 32252 15884 32280
rect 16482 32240 16488 32292
rect 16540 32280 16546 32292
rect 18049 32283 18107 32289
rect 18049 32280 18061 32283
rect 16540 32252 18061 32280
rect 16540 32240 16546 32252
rect 18049 32249 18061 32252
rect 18095 32249 18107 32283
rect 18049 32243 18107 32249
rect 19242 32240 19248 32292
rect 19300 32280 19306 32292
rect 20254 32280 20260 32292
rect 19300 32252 20260 32280
rect 19300 32240 19306 32252
rect 20254 32240 20260 32252
rect 20312 32280 20318 32292
rect 20364 32280 20392 32311
rect 20530 32308 20536 32320
rect 20588 32308 20594 32360
rect 21468 32280 21496 32379
rect 22462 32308 22468 32360
rect 22520 32308 22526 32360
rect 22756 32348 22784 32379
rect 23934 32376 23940 32428
rect 23992 32376 23998 32428
rect 24026 32376 24032 32428
rect 24084 32376 24090 32428
rect 24302 32376 24308 32428
rect 24360 32376 24366 32428
rect 24578 32376 24584 32428
rect 24636 32416 24642 32428
rect 24636 32388 24900 32416
rect 24636 32376 24642 32388
rect 24872 32348 24900 32388
rect 24946 32376 24952 32428
rect 25004 32376 25010 32428
rect 25041 32419 25099 32425
rect 25041 32385 25053 32419
rect 25087 32416 25099 32419
rect 25222 32416 25228 32428
rect 25087 32388 25228 32416
rect 25087 32385 25099 32388
rect 25041 32379 25099 32385
rect 25222 32376 25228 32388
rect 25280 32376 25286 32428
rect 25314 32376 25320 32428
rect 25372 32376 25378 32428
rect 25866 32376 25872 32428
rect 25924 32416 25930 32428
rect 25961 32419 26019 32425
rect 25961 32416 25973 32419
rect 25924 32388 25973 32416
rect 25924 32376 25930 32388
rect 25961 32385 25973 32388
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 26053 32419 26111 32425
rect 26053 32385 26065 32419
rect 26099 32416 26111 32419
rect 26252 32416 26280 32456
rect 27246 32444 27252 32456
rect 27304 32444 27310 32496
rect 26099 32388 26280 32416
rect 26329 32419 26387 32425
rect 26099 32385 26111 32388
rect 26053 32379 26111 32385
rect 26329 32385 26341 32419
rect 26375 32416 26387 32419
rect 26970 32416 26976 32428
rect 26375 32388 26976 32416
rect 26375 32385 26387 32388
rect 26329 32379 26387 32385
rect 26970 32376 26976 32388
rect 27028 32416 27034 32428
rect 28092 32416 28120 32524
rect 28994 32512 29000 32524
rect 29052 32512 29058 32564
rect 29270 32552 29276 32564
rect 29196 32524 29276 32552
rect 28258 32444 28264 32496
rect 28316 32444 28322 32496
rect 28534 32444 28540 32496
rect 28592 32484 28598 32496
rect 29196 32493 29224 32524
rect 29270 32512 29276 32524
rect 29328 32512 29334 32564
rect 29546 32512 29552 32564
rect 29604 32552 29610 32564
rect 29604 32524 30236 32552
rect 29604 32512 29610 32524
rect 29181 32487 29239 32493
rect 28592 32456 29040 32484
rect 28592 32444 28598 32456
rect 27028 32388 28120 32416
rect 28169 32419 28227 32425
rect 27028 32376 27034 32388
rect 28169 32385 28181 32419
rect 28215 32385 28227 32419
rect 28276 32416 28304 32444
rect 29012 32425 29040 32456
rect 29181 32453 29193 32487
rect 29227 32453 29239 32487
rect 29181 32447 29239 32453
rect 28353 32419 28411 32425
rect 28353 32416 28365 32419
rect 28276 32388 28365 32416
rect 28169 32379 28227 32385
rect 28353 32385 28365 32388
rect 28399 32385 28411 32419
rect 28353 32379 28411 32385
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 28998 32419 29056 32425
rect 28998 32385 29010 32419
rect 29044 32385 29056 32419
rect 28998 32379 29056 32385
rect 28184 32348 28212 32379
rect 22756 32320 24808 32348
rect 24872 32320 28212 32348
rect 24780 32289 24808 32320
rect 24765 32283 24823 32289
rect 20312 32252 21496 32280
rect 22066 32252 23888 32280
rect 20312 32240 20318 32252
rect 12897 32215 12955 32221
rect 12897 32181 12909 32215
rect 12943 32212 12955 32215
rect 13078 32212 13084 32224
rect 12943 32184 13084 32212
rect 12943 32181 12955 32184
rect 12897 32175 12955 32181
rect 13078 32172 13084 32184
rect 13136 32212 13142 32224
rect 13446 32212 13452 32224
rect 13136 32184 13452 32212
rect 13136 32172 13142 32184
rect 13446 32172 13452 32184
rect 13504 32172 13510 32224
rect 14921 32215 14979 32221
rect 14921 32181 14933 32215
rect 14967 32212 14979 32215
rect 15194 32212 15200 32224
rect 14967 32184 15200 32212
rect 14967 32181 14979 32184
rect 14921 32175 14979 32181
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 16942 32172 16948 32224
rect 17000 32212 17006 32224
rect 17221 32215 17279 32221
rect 17221 32212 17233 32215
rect 17000 32184 17233 32212
rect 17000 32172 17006 32184
rect 17221 32181 17233 32184
rect 17267 32181 17279 32215
rect 17221 32175 17279 32181
rect 18690 32172 18696 32224
rect 18748 32212 18754 32224
rect 22066 32212 22094 32252
rect 18748 32184 22094 32212
rect 18748 32172 18754 32184
rect 22554 32172 22560 32224
rect 22612 32172 22618 32224
rect 23290 32172 23296 32224
rect 23348 32172 23354 32224
rect 23750 32172 23756 32224
rect 23808 32172 23814 32224
rect 23860 32212 23888 32252
rect 24765 32249 24777 32283
rect 24811 32249 24823 32283
rect 24765 32243 24823 32249
rect 24946 32240 24952 32292
rect 25004 32280 25010 32292
rect 25866 32280 25872 32292
rect 25004 32252 25872 32280
rect 25004 32240 25010 32252
rect 25866 32240 25872 32252
rect 25924 32240 25930 32292
rect 26234 32240 26240 32292
rect 26292 32280 26298 32292
rect 26786 32280 26792 32292
rect 26292 32252 26792 32280
rect 26292 32240 26298 32252
rect 26786 32240 26792 32252
rect 26844 32240 26850 32292
rect 27062 32240 27068 32292
rect 27120 32280 27126 32292
rect 27246 32280 27252 32292
rect 27120 32252 27252 32280
rect 27120 32240 27126 32252
rect 27246 32240 27252 32252
rect 27304 32240 27310 32292
rect 28184 32280 28212 32320
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32348 28319 32351
rect 28920 32348 28948 32379
rect 29270 32376 29276 32428
rect 29328 32376 29334 32428
rect 29411 32419 29469 32425
rect 29411 32385 29423 32419
rect 29457 32416 29469 32419
rect 29638 32416 29644 32428
rect 29457 32388 29644 32416
rect 29457 32385 29469 32388
rect 29411 32379 29469 32385
rect 29638 32376 29644 32388
rect 29696 32416 29702 32428
rect 29696 32388 29960 32416
rect 29696 32376 29702 32388
rect 28307 32320 28948 32348
rect 29932 32348 29960 32388
rect 30006 32376 30012 32428
rect 30064 32376 30070 32428
rect 30208 32425 30236 32524
rect 30374 32512 30380 32564
rect 30432 32552 30438 32564
rect 31938 32552 31944 32564
rect 30432 32524 31944 32552
rect 30432 32512 30438 32524
rect 31938 32512 31944 32524
rect 31996 32512 32002 32564
rect 32030 32512 32036 32564
rect 32088 32552 32094 32564
rect 32398 32552 32404 32564
rect 32088 32524 32404 32552
rect 32088 32512 32094 32524
rect 32398 32512 32404 32524
rect 32456 32552 32462 32564
rect 33603 32555 33661 32561
rect 32456 32524 33456 32552
rect 32456 32512 32462 32524
rect 30466 32444 30472 32496
rect 30524 32484 30530 32496
rect 30929 32487 30987 32493
rect 30929 32484 30941 32487
rect 30524 32456 30941 32484
rect 30524 32444 30530 32456
rect 30929 32453 30941 32456
rect 30975 32453 30987 32487
rect 30929 32447 30987 32453
rect 31113 32487 31171 32493
rect 31113 32453 31125 32487
rect 31159 32484 31171 32487
rect 31159 32456 31708 32484
rect 31159 32453 31171 32456
rect 31113 32447 31171 32453
rect 30193 32419 30251 32425
rect 30193 32385 30205 32419
rect 30239 32385 30251 32419
rect 30193 32379 30251 32385
rect 30282 32376 30288 32428
rect 30340 32416 30346 32428
rect 30837 32419 30895 32425
rect 30837 32416 30849 32419
rect 30340 32388 30849 32416
rect 30340 32376 30346 32388
rect 30837 32385 30849 32388
rect 30883 32416 30895 32419
rect 31573 32419 31631 32425
rect 30883 32388 30972 32416
rect 30883 32385 30895 32388
rect 30837 32379 30895 32385
rect 30944 32360 30972 32388
rect 31573 32385 31585 32419
rect 31619 32385 31631 32419
rect 31573 32379 31631 32385
rect 30374 32348 30380 32360
rect 29932 32320 30380 32348
rect 28307 32317 28319 32320
rect 28261 32311 28319 32317
rect 30374 32308 30380 32320
rect 30432 32308 30438 32360
rect 30926 32308 30932 32360
rect 30984 32308 30990 32360
rect 29638 32280 29644 32292
rect 28184 32252 29644 32280
rect 29638 32240 29644 32252
rect 29696 32280 29702 32292
rect 30006 32280 30012 32292
rect 29696 32252 30012 32280
rect 29696 32240 29702 32252
rect 30006 32240 30012 32252
rect 30064 32240 30070 32292
rect 30098 32240 30104 32292
rect 30156 32280 30162 32292
rect 30193 32283 30251 32289
rect 30193 32280 30205 32283
rect 30156 32252 30205 32280
rect 30156 32240 30162 32252
rect 30193 32249 30205 32252
rect 30239 32249 30251 32283
rect 31588 32280 31616 32379
rect 31680 32348 31708 32456
rect 32122 32444 32128 32496
rect 32180 32484 32186 32496
rect 32685 32487 32743 32493
rect 32685 32484 32697 32487
rect 32180 32456 32697 32484
rect 32180 32444 32186 32456
rect 32685 32453 32697 32456
rect 32731 32453 32743 32487
rect 32685 32447 32743 32453
rect 31757 32419 31815 32425
rect 31757 32385 31769 32419
rect 31803 32416 31815 32419
rect 32030 32416 32036 32428
rect 31803 32388 32036 32416
rect 31803 32385 31815 32388
rect 31757 32379 31815 32385
rect 32030 32376 32036 32388
rect 32088 32376 32094 32428
rect 32398 32376 32404 32428
rect 32456 32422 32462 32428
rect 32561 32422 32619 32425
rect 32456 32419 32628 32422
rect 32456 32394 32573 32419
rect 32456 32376 32462 32394
rect 32561 32385 32573 32394
rect 32607 32388 32628 32419
rect 32769 32419 32827 32425
rect 32607 32385 32619 32388
rect 32561 32379 32619 32385
rect 32769 32385 32781 32419
rect 32815 32416 32827 32419
rect 32858 32416 32864 32428
rect 32815 32388 32864 32416
rect 32815 32385 32827 32388
rect 32769 32379 32827 32385
rect 32858 32376 32864 32388
rect 32916 32376 32922 32428
rect 32953 32419 33011 32425
rect 32953 32385 32965 32419
rect 32999 32416 33011 32419
rect 33226 32416 33232 32428
rect 32999 32388 33232 32416
rect 32999 32385 33011 32388
rect 32953 32379 33011 32385
rect 33226 32376 33232 32388
rect 33284 32376 33290 32428
rect 33428 32416 33456 32524
rect 33603 32521 33615 32555
rect 33649 32552 33661 32555
rect 33962 32552 33968 32564
rect 33649 32524 33968 32552
rect 33649 32521 33661 32524
rect 33603 32515 33661 32521
rect 33962 32512 33968 32524
rect 34020 32512 34026 32564
rect 34330 32512 34336 32564
rect 34388 32512 34394 32564
rect 37458 32512 37464 32564
rect 37516 32512 37522 32564
rect 39850 32552 39856 32564
rect 37752 32524 39856 32552
rect 33502 32444 33508 32496
rect 33560 32444 33566 32496
rect 37182 32484 37188 32496
rect 33612 32456 37188 32484
rect 33612 32416 33640 32456
rect 33428 32388 33640 32416
rect 33686 32376 33692 32428
rect 33744 32376 33750 32428
rect 33778 32376 33784 32428
rect 33836 32376 33842 32428
rect 35084 32425 35112 32456
rect 37182 32444 37188 32456
rect 37240 32444 37246 32496
rect 35069 32419 35127 32425
rect 35069 32385 35081 32419
rect 35115 32385 35127 32419
rect 35069 32379 35127 32385
rect 35158 32376 35164 32428
rect 35216 32376 35222 32428
rect 35253 32419 35311 32425
rect 35253 32385 35265 32419
rect 35299 32385 35311 32419
rect 35253 32379 35311 32385
rect 35268 32348 35296 32379
rect 35434 32376 35440 32428
rect 35492 32376 35498 32428
rect 35989 32419 36047 32425
rect 35989 32385 36001 32419
rect 36035 32385 36047 32419
rect 35989 32379 36047 32385
rect 31680 32320 34928 32348
rect 34422 32280 34428 32292
rect 31588 32252 34428 32280
rect 30193 32243 30251 32249
rect 34422 32240 34428 32252
rect 34480 32240 34486 32292
rect 34900 32289 34928 32320
rect 35176 32320 35296 32348
rect 36004 32348 36032 32379
rect 36078 32376 36084 32428
rect 36136 32376 36142 32428
rect 36170 32376 36176 32428
rect 36228 32416 36234 32428
rect 37752 32425 37780 32524
rect 39850 32512 39856 32524
rect 39908 32512 39914 32564
rect 40954 32512 40960 32564
rect 41012 32552 41018 32564
rect 42058 32552 42064 32564
rect 41012 32524 42064 32552
rect 41012 32512 41018 32524
rect 42058 32512 42064 32524
rect 42116 32512 42122 32564
rect 43070 32512 43076 32564
rect 43128 32552 43134 32564
rect 43257 32555 43315 32561
rect 43257 32552 43269 32555
rect 43128 32524 43269 32552
rect 43128 32512 43134 32524
rect 43257 32521 43269 32524
rect 43303 32552 43315 32555
rect 43346 32552 43352 32564
rect 43303 32524 43352 32552
rect 43303 32521 43315 32524
rect 43257 32515 43315 32521
rect 43346 32512 43352 32524
rect 43404 32512 43410 32564
rect 38286 32484 38292 32496
rect 37936 32456 38292 32484
rect 36265 32419 36323 32425
rect 36265 32416 36277 32419
rect 36228 32388 36277 32416
rect 36228 32376 36234 32388
rect 36265 32385 36277 32388
rect 36311 32385 36323 32419
rect 36265 32379 36323 32385
rect 37737 32419 37795 32425
rect 37737 32385 37749 32419
rect 37783 32385 37795 32419
rect 37737 32379 37795 32385
rect 37826 32376 37832 32428
rect 37884 32376 37890 32428
rect 37936 32425 37964 32456
rect 38286 32444 38292 32456
rect 38344 32484 38350 32496
rect 39298 32484 39304 32496
rect 38344 32456 39304 32484
rect 38344 32444 38350 32456
rect 39298 32444 39304 32456
rect 39356 32444 39362 32496
rect 39390 32444 39396 32496
rect 39448 32484 39454 32496
rect 41230 32484 41236 32496
rect 39448 32456 41236 32484
rect 39448 32444 39454 32456
rect 37921 32419 37979 32425
rect 37921 32385 37933 32419
rect 37967 32385 37979 32419
rect 37921 32379 37979 32385
rect 38105 32419 38163 32425
rect 38105 32385 38117 32419
rect 38151 32385 38163 32419
rect 38105 32379 38163 32385
rect 36354 32348 36360 32360
rect 36004 32320 36360 32348
rect 34885 32283 34943 32289
rect 34885 32249 34897 32283
rect 34931 32249 34943 32283
rect 34885 32243 34943 32249
rect 25590 32212 25596 32224
rect 23860 32184 25596 32212
rect 25590 32172 25596 32184
rect 25648 32172 25654 32224
rect 26804 32212 26832 32240
rect 28442 32212 28448 32224
rect 26804 32184 28448 32212
rect 28442 32172 28448 32184
rect 28500 32172 28506 32224
rect 28718 32172 28724 32224
rect 28776 32212 28782 32224
rect 29549 32215 29607 32221
rect 29549 32212 29561 32215
rect 28776 32184 29561 32212
rect 28776 32172 28782 32184
rect 29549 32181 29561 32184
rect 29595 32181 29607 32215
rect 29549 32175 29607 32181
rect 30374 32172 30380 32224
rect 30432 32212 30438 32224
rect 31113 32215 31171 32221
rect 31113 32212 31125 32215
rect 30432 32184 31125 32212
rect 30432 32172 30438 32184
rect 31113 32181 31125 32184
rect 31159 32181 31171 32215
rect 31113 32175 31171 32181
rect 31573 32215 31631 32221
rect 31573 32181 31585 32215
rect 31619 32212 31631 32215
rect 32306 32212 32312 32224
rect 31619 32184 32312 32212
rect 31619 32181 31631 32184
rect 31573 32175 31631 32181
rect 32306 32172 32312 32184
rect 32364 32172 32370 32224
rect 32398 32172 32404 32224
rect 32456 32172 32462 32224
rect 32766 32172 32772 32224
rect 32824 32212 32830 32224
rect 33134 32212 33140 32224
rect 32824 32184 33140 32212
rect 32824 32172 32830 32184
rect 33134 32172 33140 32184
rect 33192 32212 33198 32224
rect 33778 32212 33784 32224
rect 33192 32184 33784 32212
rect 33192 32172 33198 32184
rect 33778 32172 33784 32184
rect 33836 32172 33842 32224
rect 34238 32172 34244 32224
rect 34296 32212 34302 32224
rect 35176 32212 35204 32320
rect 36354 32308 36360 32320
rect 36412 32308 36418 32360
rect 36446 32308 36452 32360
rect 36504 32348 36510 32360
rect 36725 32351 36783 32357
rect 36725 32348 36737 32351
rect 36504 32320 36737 32348
rect 36504 32308 36510 32320
rect 36725 32317 36737 32320
rect 36771 32317 36783 32351
rect 36725 32311 36783 32317
rect 37090 32308 37096 32360
rect 37148 32348 37154 32360
rect 38120 32348 38148 32379
rect 39114 32376 39120 32428
rect 39172 32376 39178 32428
rect 40328 32425 40356 32456
rect 41230 32444 41236 32456
rect 41288 32484 41294 32496
rect 41509 32487 41567 32493
rect 41509 32484 41521 32487
rect 41288 32456 41521 32484
rect 41288 32444 41294 32456
rect 41509 32453 41521 32456
rect 41555 32453 41567 32487
rect 41509 32447 41567 32453
rect 39485 32419 39543 32425
rect 39485 32385 39497 32419
rect 39531 32416 39543 32419
rect 40221 32419 40279 32425
rect 40221 32416 40233 32419
rect 39531 32388 40233 32416
rect 39531 32385 39543 32388
rect 39485 32379 39543 32385
rect 40221 32385 40233 32388
rect 40267 32385 40279 32419
rect 40221 32379 40279 32385
rect 40313 32419 40371 32425
rect 40313 32385 40325 32419
rect 40359 32385 40371 32419
rect 40313 32379 40371 32385
rect 40586 32376 40592 32428
rect 40644 32376 40650 32428
rect 40770 32376 40776 32428
rect 40828 32416 40834 32428
rect 41417 32419 41475 32425
rect 41417 32416 41429 32419
rect 40828 32388 41429 32416
rect 40828 32376 40834 32388
rect 41417 32385 41429 32388
rect 41463 32385 41475 32419
rect 41417 32379 41475 32385
rect 41598 32376 41604 32428
rect 41656 32376 41662 32428
rect 42797 32419 42855 32425
rect 42797 32385 42809 32419
rect 42843 32416 42855 32419
rect 43254 32416 43260 32428
rect 42843 32388 43260 32416
rect 42843 32385 42855 32388
rect 42797 32379 42855 32385
rect 43254 32376 43260 32388
rect 43312 32376 43318 32428
rect 37148 32320 38148 32348
rect 38749 32351 38807 32357
rect 37148 32308 37154 32320
rect 38749 32317 38761 32351
rect 38795 32348 38807 32351
rect 40034 32348 40040 32360
rect 38795 32320 40040 32348
rect 38795 32317 38807 32320
rect 38749 32311 38807 32317
rect 40034 32308 40040 32320
rect 40092 32308 40098 32360
rect 40129 32351 40187 32357
rect 40129 32317 40141 32351
rect 40175 32317 40187 32351
rect 40129 32311 40187 32317
rect 35802 32240 35808 32292
rect 35860 32280 35866 32292
rect 39022 32280 39028 32292
rect 35860 32252 39028 32280
rect 35860 32240 35866 32252
rect 39022 32240 39028 32252
rect 39080 32280 39086 32292
rect 39390 32280 39396 32292
rect 39080 32252 39396 32280
rect 39080 32240 39086 32252
rect 39390 32240 39396 32252
rect 39448 32240 39454 32292
rect 39482 32240 39488 32292
rect 39540 32240 39546 32292
rect 34296 32184 35204 32212
rect 34296 32172 34302 32184
rect 35434 32172 35440 32224
rect 35492 32212 35498 32224
rect 40144 32212 40172 32311
rect 40494 32308 40500 32360
rect 40552 32348 40558 32360
rect 40957 32351 41015 32357
rect 40957 32348 40969 32351
rect 40552 32320 40969 32348
rect 40552 32308 40558 32320
rect 40957 32317 40969 32320
rect 41003 32317 41015 32351
rect 40957 32311 41015 32317
rect 35492 32184 40172 32212
rect 42613 32215 42671 32221
rect 35492 32172 35498 32184
rect 42613 32181 42625 32215
rect 42659 32212 42671 32215
rect 42886 32212 42892 32224
rect 42659 32184 42892 32212
rect 42659 32181 42671 32184
rect 42613 32175 42671 32181
rect 42886 32172 42892 32184
rect 42944 32172 42950 32224
rect 1104 32122 43884 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 43884 32122
rect 1104 32048 43884 32070
rect 12618 31968 12624 32020
rect 12676 32008 12682 32020
rect 13081 32011 13139 32017
rect 13081 32008 13093 32011
rect 12676 31980 13093 32008
rect 12676 31968 12682 31980
rect 13081 31977 13093 31980
rect 13127 31977 13139 32011
rect 13081 31971 13139 31977
rect 13262 31968 13268 32020
rect 13320 31968 13326 32020
rect 14274 31968 14280 32020
rect 14332 31968 14338 32020
rect 14550 31968 14556 32020
rect 14608 32008 14614 32020
rect 15841 32011 15899 32017
rect 15841 32008 15853 32011
rect 14608 31980 15853 32008
rect 14608 31968 14614 31980
rect 15841 31977 15853 31980
rect 15887 31977 15899 32011
rect 15841 31971 15899 31977
rect 17034 31968 17040 32020
rect 17092 32008 17098 32020
rect 20714 32008 20720 32020
rect 17092 31980 20720 32008
rect 17092 31968 17098 31980
rect 20714 31968 20720 31980
rect 20772 31968 20778 32020
rect 26697 32011 26755 32017
rect 26697 32008 26709 32011
rect 20824 31980 26709 32008
rect 12710 31900 12716 31952
rect 12768 31940 12774 31952
rect 13280 31940 13308 31968
rect 12768 31912 13308 31940
rect 12768 31900 12774 31912
rect 14090 31900 14096 31952
rect 14148 31940 14154 31952
rect 14148 31912 14412 31940
rect 14148 31900 14154 31912
rect 12529 31875 12587 31881
rect 12529 31841 12541 31875
rect 12575 31872 12587 31875
rect 14182 31872 14188 31884
rect 12575 31844 14188 31872
rect 12575 31841 12587 31844
rect 12529 31835 12587 31841
rect 14182 31832 14188 31844
rect 14240 31832 14246 31884
rect 12437 31807 12495 31813
rect 12437 31773 12449 31807
rect 12483 31804 12495 31807
rect 12483 31776 12572 31804
rect 12483 31773 12495 31776
rect 12437 31767 12495 31773
rect 12544 31736 12572 31776
rect 12618 31764 12624 31816
rect 12676 31764 12682 31816
rect 13354 31804 13360 31816
rect 12728 31776 13360 31804
rect 12728 31736 12756 31776
rect 13280 31745 13308 31776
rect 13354 31764 13360 31776
rect 13412 31764 13418 31816
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31806 14335 31807
rect 14384 31806 14412 31912
rect 15378 31900 15384 31952
rect 15436 31900 15442 31952
rect 17218 31900 17224 31952
rect 17276 31940 17282 31952
rect 17589 31943 17647 31949
rect 17589 31940 17601 31943
rect 17276 31912 17601 31940
rect 17276 31900 17282 31912
rect 17589 31909 17601 31912
rect 17635 31909 17647 31943
rect 17589 31903 17647 31909
rect 19058 31900 19064 31952
rect 19116 31940 19122 31952
rect 19429 31943 19487 31949
rect 19429 31940 19441 31943
rect 19116 31912 19441 31940
rect 19116 31900 19122 31912
rect 19429 31909 19441 31912
rect 19475 31909 19487 31943
rect 19429 31903 19487 31909
rect 20622 31900 20628 31952
rect 20680 31940 20686 31952
rect 20824 31940 20852 31980
rect 26697 31977 26709 31980
rect 26743 31977 26755 32011
rect 26697 31971 26755 31977
rect 26970 31968 26976 32020
rect 27028 32008 27034 32020
rect 29822 32008 29828 32020
rect 27028 31980 29828 32008
rect 27028 31968 27034 31980
rect 29822 31968 29828 31980
rect 29880 31968 29886 32020
rect 30193 32011 30251 32017
rect 30193 31977 30205 32011
rect 30239 32008 30251 32011
rect 30282 32008 30288 32020
rect 30239 31980 30288 32008
rect 30239 31977 30251 31980
rect 30193 31971 30251 31977
rect 30282 31968 30288 31980
rect 30340 31968 30346 32020
rect 31849 32011 31907 32017
rect 31849 32008 31861 32011
rect 31726 31980 31861 32008
rect 20680 31912 20852 31940
rect 20680 31900 20686 31912
rect 24762 31900 24768 31952
rect 24820 31940 24826 31952
rect 28721 31943 28779 31949
rect 28721 31940 28733 31943
rect 24820 31912 28733 31940
rect 24820 31900 24826 31912
rect 28721 31909 28733 31912
rect 28767 31909 28779 31943
rect 28721 31903 28779 31909
rect 28810 31900 28816 31952
rect 28868 31940 28874 31952
rect 31726 31940 31754 31980
rect 31849 31977 31861 31980
rect 31895 31977 31907 32011
rect 31849 31971 31907 31977
rect 32306 31968 32312 32020
rect 32364 32008 32370 32020
rect 32766 32008 32772 32020
rect 32364 31980 32772 32008
rect 32364 31968 32370 31980
rect 32766 31968 32772 31980
rect 32824 31968 32830 32020
rect 34238 32008 34244 32020
rect 32876 31980 34244 32008
rect 28868 31912 31754 31940
rect 28868 31900 28874 31912
rect 31938 31900 31944 31952
rect 31996 31940 32002 31952
rect 32876 31940 32904 31980
rect 34238 31968 34244 31980
rect 34296 31968 34302 32020
rect 34606 31968 34612 32020
rect 34664 32008 34670 32020
rect 34885 32011 34943 32017
rect 34885 32008 34897 32011
rect 34664 31980 34897 32008
rect 34664 31968 34670 31980
rect 34885 31977 34897 31980
rect 34931 31977 34943 32011
rect 34885 31971 34943 31977
rect 36541 32011 36599 32017
rect 36541 31977 36553 32011
rect 36587 32008 36599 32011
rect 37090 32008 37096 32020
rect 36587 31980 37096 32008
rect 36587 31977 36599 31980
rect 36541 31971 36599 31977
rect 37090 31968 37096 31980
rect 37148 31968 37154 32020
rect 37642 31968 37648 32020
rect 37700 31968 37706 32020
rect 37826 31968 37832 32020
rect 37884 31968 37890 32020
rect 38197 32011 38255 32017
rect 38197 31977 38209 32011
rect 38243 32008 38255 32011
rect 39206 32008 39212 32020
rect 38243 31980 39212 32008
rect 38243 31977 38255 31980
rect 38197 31971 38255 31977
rect 39206 31968 39212 31980
rect 39264 31968 39270 32020
rect 39850 31968 39856 32020
rect 39908 32008 39914 32020
rect 40586 32008 40592 32020
rect 39908 31980 40592 32008
rect 39908 31968 39914 31980
rect 31996 31912 32904 31940
rect 32953 31943 33011 31949
rect 31996 31900 32002 31912
rect 32953 31909 32965 31943
rect 32999 31940 33011 31943
rect 34149 31943 34207 31949
rect 32999 31912 34100 31940
rect 32999 31909 33011 31912
rect 32953 31903 33011 31909
rect 16298 31872 16304 31884
rect 15028 31844 16304 31872
rect 14323 31778 14412 31806
rect 14323 31773 14335 31778
rect 14277 31767 14335 31773
rect 14458 31764 14464 31816
rect 14516 31764 14522 31816
rect 15028 31813 15056 31844
rect 16298 31832 16304 31844
rect 16356 31832 16362 31884
rect 16485 31875 16543 31881
rect 16485 31841 16497 31875
rect 16531 31872 16543 31875
rect 18233 31875 18291 31881
rect 16531 31844 18184 31872
rect 16531 31841 16543 31844
rect 16485 31835 16543 31841
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31773 15071 31807
rect 15013 31767 15071 31773
rect 15194 31764 15200 31816
rect 15252 31804 15258 31816
rect 16209 31807 16267 31813
rect 16209 31804 16221 31807
rect 15252 31776 16221 31804
rect 15252 31764 15258 31776
rect 16209 31773 16221 31776
rect 16255 31773 16267 31807
rect 18046 31804 18052 31816
rect 16209 31767 16267 31773
rect 16592 31776 18052 31804
rect 12544 31708 12756 31736
rect 13249 31739 13308 31745
rect 13249 31705 13261 31739
rect 13295 31708 13308 31739
rect 13295 31705 13307 31708
rect 13249 31699 13307 31705
rect 13446 31696 13452 31748
rect 13504 31696 13510 31748
rect 16592 31736 16620 31776
rect 18046 31764 18052 31776
rect 18104 31764 18110 31816
rect 18156 31804 18184 31844
rect 18233 31841 18245 31875
rect 18279 31872 18291 31875
rect 18279 31844 19104 31872
rect 18279 31841 18291 31844
rect 18233 31835 18291 31841
rect 19076 31816 19104 31844
rect 19978 31832 19984 31884
rect 20036 31832 20042 31884
rect 20346 31832 20352 31884
rect 20404 31872 20410 31884
rect 20717 31875 20775 31881
rect 20717 31872 20729 31875
rect 20404 31844 20729 31872
rect 20404 31832 20410 31844
rect 20717 31841 20729 31844
rect 20763 31841 20775 31875
rect 20717 31835 20775 31841
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 20956 31844 21864 31872
rect 20956 31832 20962 31844
rect 18156 31776 18828 31804
rect 16500 31708 16620 31736
rect 15930 31628 15936 31680
rect 15988 31668 15994 31680
rect 16301 31671 16359 31677
rect 16301 31668 16313 31671
rect 15988 31640 16313 31668
rect 15988 31628 15994 31640
rect 16301 31637 16313 31640
rect 16347 31668 16359 31671
rect 16500 31668 16528 31708
rect 17862 31696 17868 31748
rect 17920 31736 17926 31748
rect 18800 31736 18828 31776
rect 18874 31764 18880 31816
rect 18932 31764 18938 31816
rect 19058 31764 19064 31816
rect 19116 31764 19122 31816
rect 20530 31804 20536 31816
rect 19168 31776 20536 31804
rect 19168 31736 19196 31776
rect 20530 31764 20536 31776
rect 20588 31764 20594 31816
rect 20809 31807 20867 31813
rect 20809 31773 20821 31807
rect 20855 31804 20867 31807
rect 21082 31804 21088 31816
rect 20855 31776 21088 31804
rect 20855 31773 20867 31776
rect 20809 31767 20867 31773
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 21358 31764 21364 31816
rect 21416 31804 21422 31816
rect 21729 31807 21787 31813
rect 21729 31804 21741 31807
rect 21416 31776 21741 31804
rect 21416 31764 21422 31776
rect 21729 31773 21741 31776
rect 21775 31773 21787 31807
rect 21836 31804 21864 31844
rect 21910 31832 21916 31884
rect 21968 31872 21974 31884
rect 23109 31875 23167 31881
rect 23109 31872 23121 31875
rect 21968 31844 23121 31872
rect 21968 31832 21974 31844
rect 23109 31841 23121 31844
rect 23155 31841 23167 31875
rect 25038 31872 25044 31884
rect 23109 31835 23167 31841
rect 23952 31844 25044 31872
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21836 31776 22017 31804
rect 21729 31767 21787 31773
rect 22005 31773 22017 31776
rect 22051 31804 22063 31807
rect 23014 31804 23020 31816
rect 22051 31776 23020 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 23290 31764 23296 31816
rect 23348 31804 23354 31816
rect 23952 31813 23980 31844
rect 25038 31832 25044 31844
rect 25096 31832 25102 31884
rect 30098 31872 30104 31884
rect 25884 31844 30104 31872
rect 25884 31816 25912 31844
rect 23937 31807 23995 31813
rect 23937 31804 23949 31807
rect 23348 31776 23949 31804
rect 23348 31764 23354 31776
rect 23937 31773 23949 31776
rect 23983 31773 23995 31807
rect 23937 31767 23995 31773
rect 24210 31764 24216 31816
rect 24268 31804 24274 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 24268 31776 24777 31804
rect 24268 31764 24274 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 24946 31764 24952 31816
rect 25004 31764 25010 31816
rect 25130 31764 25136 31816
rect 25188 31764 25194 31816
rect 25225 31807 25283 31813
rect 25225 31773 25237 31807
rect 25271 31804 25283 31807
rect 25866 31804 25872 31816
rect 25271 31776 25305 31804
rect 25827 31776 25872 31804
rect 25271 31773 25283 31776
rect 25225 31767 25283 31773
rect 20898 31736 20904 31748
rect 17920 31708 18092 31736
rect 18800 31708 19196 31736
rect 19260 31708 20904 31736
rect 17920 31696 17926 31708
rect 16347 31640 16528 31668
rect 16347 31637 16359 31640
rect 16301 31631 16359 31637
rect 17954 31628 17960 31680
rect 18012 31628 18018 31680
rect 18064 31668 18092 31708
rect 19260 31680 19288 31708
rect 20898 31696 20904 31708
rect 20956 31696 20962 31748
rect 21821 31739 21879 31745
rect 21821 31705 21833 31739
rect 21867 31736 21879 31739
rect 22370 31736 22376 31748
rect 21867 31708 22376 31736
rect 21867 31705 21879 31708
rect 21821 31699 21879 31705
rect 22370 31696 22376 31708
rect 22428 31696 22434 31748
rect 23658 31696 23664 31748
rect 23716 31736 23722 31748
rect 24578 31736 24584 31748
rect 23716 31708 24584 31736
rect 23716 31696 23722 31708
rect 24578 31696 24584 31708
rect 24636 31736 24642 31748
rect 25240 31736 25268 31767
rect 25866 31764 25872 31776
rect 25924 31764 25930 31816
rect 26237 31807 26295 31813
rect 26237 31773 26249 31807
rect 26283 31804 26295 31807
rect 26786 31804 26792 31816
rect 26283 31776 26792 31804
rect 26283 31773 26295 31776
rect 26237 31767 26295 31773
rect 26786 31764 26792 31776
rect 26844 31764 26850 31816
rect 26896 31813 26924 31844
rect 30098 31832 30104 31844
rect 30156 31832 30162 31884
rect 32125 31875 32183 31881
rect 32125 31841 32137 31875
rect 32171 31872 32183 31875
rect 33134 31872 33140 31884
rect 32171 31844 33140 31872
rect 32171 31841 32183 31844
rect 32125 31835 32183 31841
rect 33134 31832 33140 31844
rect 33192 31832 33198 31884
rect 33226 31832 33232 31884
rect 33284 31832 33290 31884
rect 26881 31807 26939 31813
rect 26881 31773 26893 31807
rect 26927 31773 26939 31807
rect 26881 31767 26939 31773
rect 26970 31764 26976 31816
rect 27028 31764 27034 31816
rect 27065 31807 27123 31813
rect 27065 31773 27077 31807
rect 27111 31773 27123 31807
rect 27065 31767 27123 31773
rect 24636 31708 25268 31736
rect 25961 31739 26019 31745
rect 24636 31696 24642 31708
rect 25961 31705 25973 31739
rect 26007 31705 26019 31739
rect 25961 31699 26019 31705
rect 18230 31668 18236 31680
rect 18064 31640 18236 31668
rect 18230 31628 18236 31640
rect 18288 31668 18294 31680
rect 19242 31668 19248 31680
rect 18288 31640 19248 31668
rect 18288 31628 18294 31640
rect 19242 31628 19248 31640
rect 19300 31628 19306 31680
rect 19794 31628 19800 31680
rect 19852 31628 19858 31680
rect 19889 31671 19947 31677
rect 19889 31637 19901 31671
rect 19935 31668 19947 31671
rect 20070 31668 20076 31680
rect 19935 31640 20076 31668
rect 19935 31637 19947 31640
rect 19889 31631 19947 31637
rect 20070 31628 20076 31640
rect 20128 31628 20134 31680
rect 22189 31671 22247 31677
rect 22189 31637 22201 31671
rect 22235 31668 22247 31671
rect 22278 31668 22284 31680
rect 22235 31640 22284 31668
rect 22235 31637 22247 31640
rect 22189 31631 22247 31637
rect 22278 31628 22284 31640
rect 22336 31628 22342 31680
rect 22922 31628 22928 31680
rect 22980 31668 22986 31680
rect 24670 31668 24676 31680
rect 22980 31640 24676 31668
rect 22980 31628 22986 31640
rect 24670 31628 24676 31640
rect 24728 31628 24734 31680
rect 24762 31628 24768 31680
rect 24820 31668 24826 31680
rect 25222 31668 25228 31680
rect 24820 31640 25228 31668
rect 24820 31628 24826 31640
rect 25222 31628 25228 31640
rect 25280 31628 25286 31680
rect 25590 31628 25596 31680
rect 25648 31668 25654 31680
rect 25685 31671 25743 31677
rect 25685 31668 25697 31671
rect 25648 31640 25697 31668
rect 25648 31628 25654 31640
rect 25685 31637 25697 31640
rect 25731 31637 25743 31671
rect 25976 31668 26004 31699
rect 26050 31696 26056 31748
rect 26108 31736 26114 31748
rect 27080 31736 27108 31767
rect 27246 31764 27252 31816
rect 27304 31764 27310 31816
rect 27798 31764 27804 31816
rect 27856 31804 27862 31816
rect 27856 31776 28672 31804
rect 27856 31764 27862 31776
rect 26108 31708 27108 31736
rect 27264 31736 27292 31764
rect 28534 31736 28540 31748
rect 27264 31708 28540 31736
rect 26108 31696 26114 31708
rect 26234 31668 26240 31680
rect 25976 31640 26240 31668
rect 25685 31631 25743 31637
rect 26234 31628 26240 31640
rect 26292 31628 26298 31680
rect 27080 31668 27108 31708
rect 28534 31696 28540 31708
rect 28592 31696 28598 31748
rect 28644 31736 28672 31776
rect 28718 31764 28724 31816
rect 28776 31764 28782 31816
rect 28902 31764 28908 31816
rect 28960 31764 28966 31816
rect 28997 31807 29055 31813
rect 28997 31773 29009 31807
rect 29043 31804 29055 31807
rect 29914 31804 29920 31816
rect 29043 31776 29920 31804
rect 29043 31773 29055 31776
rect 28997 31767 29055 31773
rect 29914 31764 29920 31776
rect 29972 31764 29978 31816
rect 30009 31807 30067 31813
rect 30009 31773 30021 31807
rect 30055 31804 30067 31807
rect 30190 31804 30196 31816
rect 30055 31776 30196 31804
rect 30055 31773 30067 31776
rect 30009 31767 30067 31773
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 31297 31807 31355 31813
rect 30300 31776 31248 31804
rect 30300 31736 30328 31776
rect 28644 31708 30328 31736
rect 31220 31736 31248 31776
rect 31297 31773 31309 31807
rect 31343 31804 31355 31807
rect 32030 31804 32036 31816
rect 31343 31776 32036 31804
rect 31343 31773 31355 31776
rect 31297 31767 31355 31773
rect 32030 31764 32036 31776
rect 32088 31764 32094 31816
rect 32214 31764 32220 31816
rect 32272 31804 32278 31816
rect 32309 31807 32367 31813
rect 32309 31804 32321 31807
rect 32272 31776 32321 31804
rect 32272 31764 32278 31776
rect 32309 31773 32321 31776
rect 32355 31804 32367 31807
rect 32674 31804 32680 31816
rect 32355 31776 32680 31804
rect 32355 31773 32367 31776
rect 32309 31767 32367 31773
rect 32674 31764 32680 31776
rect 32732 31764 32738 31816
rect 32766 31764 32772 31816
rect 32824 31764 32830 31816
rect 33244 31804 33272 31832
rect 33965 31807 34023 31813
rect 33965 31804 33977 31807
rect 32876 31776 33977 31804
rect 32876 31736 32904 31776
rect 33965 31773 33977 31776
rect 34011 31773 34023 31807
rect 33965 31767 34023 31773
rect 31220 31708 32904 31736
rect 34072 31736 34100 31912
rect 34149 31909 34161 31943
rect 34195 31940 34207 31943
rect 34698 31940 34704 31952
rect 34195 31912 34704 31940
rect 34195 31909 34207 31912
rect 34149 31903 34207 31909
rect 34698 31900 34704 31912
rect 34756 31940 34762 31952
rect 35434 31940 35440 31952
rect 34756 31912 35440 31940
rect 34756 31900 34762 31912
rect 35434 31900 35440 31912
rect 35492 31900 35498 31952
rect 37182 31900 37188 31952
rect 37240 31940 37246 31952
rect 37844 31940 37872 31968
rect 40310 31940 40316 31952
rect 37240 31912 40316 31940
rect 37240 31900 37246 31912
rect 34238 31832 34244 31884
rect 34296 31832 34302 31884
rect 37734 31872 37740 31884
rect 35360 31844 36308 31872
rect 34422 31764 34428 31816
rect 34480 31804 34486 31816
rect 35253 31807 35311 31813
rect 35253 31804 35265 31807
rect 34480 31776 35265 31804
rect 34480 31764 34486 31776
rect 35253 31773 35265 31776
rect 35299 31773 35311 31807
rect 35253 31767 35311 31773
rect 34606 31736 34612 31748
rect 34072 31708 34612 31736
rect 34606 31696 34612 31708
rect 34664 31696 34670 31748
rect 35066 31696 35072 31748
rect 35124 31736 35130 31748
rect 35360 31736 35388 31844
rect 35897 31807 35955 31813
rect 35897 31773 35909 31807
rect 35943 31804 35955 31807
rect 35986 31804 35992 31816
rect 35943 31776 35992 31804
rect 35943 31773 35955 31776
rect 35897 31767 35955 31773
rect 35986 31764 35992 31776
rect 36044 31764 36050 31816
rect 36078 31764 36084 31816
rect 36136 31764 36142 31816
rect 36280 31813 36308 31844
rect 36372 31844 37740 31872
rect 36173 31807 36231 31813
rect 36173 31773 36185 31807
rect 36219 31773 36231 31807
rect 36173 31767 36231 31773
rect 36265 31807 36323 31813
rect 36265 31773 36277 31807
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 35124 31708 35388 31736
rect 35124 31696 35130 31708
rect 35434 31696 35440 31748
rect 35492 31736 35498 31748
rect 35710 31736 35716 31748
rect 35492 31708 35716 31736
rect 35492 31696 35498 31708
rect 35710 31696 35716 31708
rect 35768 31696 35774 31748
rect 36188 31736 36216 31767
rect 36372 31736 36400 31844
rect 37734 31832 37740 31844
rect 37792 31832 37798 31884
rect 37844 31844 39252 31872
rect 36998 31764 37004 31816
rect 37056 31764 37062 31816
rect 37844 31813 37872 31844
rect 37829 31807 37887 31813
rect 37829 31773 37841 31807
rect 37875 31773 37887 31807
rect 37829 31767 37887 31773
rect 38010 31764 38016 31816
rect 38068 31764 38074 31816
rect 38286 31764 38292 31816
rect 38344 31764 38350 31816
rect 36188 31708 36400 31736
rect 39224 31736 39252 31844
rect 39316 31813 39344 31912
rect 40310 31900 40316 31912
rect 40368 31900 40374 31952
rect 40126 31872 40132 31884
rect 39408 31844 40132 31872
rect 39301 31807 39359 31813
rect 39301 31773 39313 31807
rect 39347 31773 39359 31807
rect 39301 31767 39359 31773
rect 39408 31736 39436 31844
rect 40126 31832 40132 31844
rect 40184 31832 40190 31884
rect 40420 31872 40448 31980
rect 40586 31968 40592 31980
rect 40644 32008 40650 32020
rect 41874 32008 41880 32020
rect 40644 31980 41880 32008
rect 40644 31968 40650 31980
rect 41874 31968 41880 31980
rect 41932 31968 41938 32020
rect 41230 31872 41236 31884
rect 40420 31844 40507 31872
rect 39485 31807 39543 31813
rect 39485 31773 39497 31807
rect 39531 31804 39543 31807
rect 40218 31804 40224 31816
rect 39531 31776 40224 31804
rect 39531 31773 39543 31776
rect 39485 31767 39543 31773
rect 40218 31764 40224 31776
rect 40276 31764 40282 31816
rect 40479 31813 40507 31844
rect 40605 31844 41236 31872
rect 40605 31813 40633 31844
rect 41230 31832 41236 31844
rect 41288 31832 41294 31884
rect 42886 31832 42892 31884
rect 42944 31832 42950 31884
rect 43162 31832 43168 31884
rect 43220 31832 43226 31884
rect 40313 31807 40371 31813
rect 40313 31773 40325 31807
rect 40359 31804 40371 31807
rect 40464 31807 40522 31813
rect 40359 31776 40393 31804
rect 40359 31773 40371 31776
rect 40313 31767 40371 31773
rect 40464 31773 40476 31807
rect 40510 31773 40522 31807
rect 40464 31767 40522 31773
rect 40589 31807 40647 31813
rect 40589 31773 40601 31807
rect 40635 31773 40647 31807
rect 40589 31767 40647 31773
rect 39224 31708 39436 31736
rect 39942 31696 39948 31748
rect 40000 31736 40006 31748
rect 40328 31736 40356 31767
rect 40678 31764 40684 31816
rect 40736 31764 40742 31816
rect 40000 31708 40356 31736
rect 40000 31696 40006 31708
rect 42426 31696 42432 31748
rect 42484 31696 42490 31748
rect 29270 31668 29276 31680
rect 27080 31640 29276 31668
rect 29270 31628 29276 31640
rect 29328 31628 29334 31680
rect 31113 31671 31171 31677
rect 31113 31637 31125 31671
rect 31159 31668 31171 31671
rect 32490 31668 32496 31680
rect 31159 31640 32496 31668
rect 31159 31637 31171 31640
rect 31113 31631 31171 31637
rect 32490 31628 32496 31640
rect 32548 31628 32554 31680
rect 33778 31628 33784 31680
rect 33836 31628 33842 31680
rect 39117 31671 39175 31677
rect 39117 31637 39129 31671
rect 39163 31668 39175 31671
rect 39390 31668 39396 31680
rect 39163 31640 39396 31668
rect 39163 31637 39175 31640
rect 39117 31631 39175 31637
rect 39390 31628 39396 31640
rect 39448 31628 39454 31680
rect 40129 31671 40187 31677
rect 40129 31637 40141 31671
rect 40175 31668 40187 31671
rect 40402 31668 40408 31680
rect 40175 31640 40408 31668
rect 40175 31637 40187 31640
rect 40129 31631 40187 31637
rect 40402 31628 40408 31640
rect 40460 31628 40466 31680
rect 41414 31628 41420 31680
rect 41472 31628 41478 31680
rect 1104 31578 43884 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 43884 31578
rect 1104 31504 43884 31526
rect 12069 31467 12127 31473
rect 12069 31433 12081 31467
rect 12115 31464 12127 31467
rect 13081 31467 13139 31473
rect 13081 31464 13093 31467
rect 12115 31436 13093 31464
rect 12115 31433 12127 31436
rect 12069 31427 12127 31433
rect 13081 31433 13093 31436
rect 13127 31433 13139 31467
rect 15289 31467 15347 31473
rect 15289 31464 15301 31467
rect 13081 31427 13139 31433
rect 14292 31436 15301 31464
rect 13262 31396 13268 31408
rect 12268 31368 13268 31396
rect 12268 31337 12296 31368
rect 13262 31356 13268 31368
rect 13320 31396 13326 31408
rect 14292 31405 14320 31436
rect 15289 31433 15301 31436
rect 15335 31433 15347 31467
rect 15289 31427 15347 31433
rect 15378 31424 15384 31476
rect 15436 31464 15442 31476
rect 15654 31464 15660 31476
rect 15436 31436 15660 31464
rect 15436 31424 15442 31436
rect 15654 31424 15660 31436
rect 15712 31464 15718 31476
rect 17954 31464 17960 31476
rect 15712 31436 17960 31464
rect 15712 31424 15718 31436
rect 17954 31424 17960 31436
rect 18012 31424 18018 31476
rect 18233 31467 18291 31473
rect 18233 31433 18245 31467
rect 18279 31464 18291 31467
rect 18506 31464 18512 31476
rect 18279 31436 18512 31464
rect 18279 31433 18291 31436
rect 18233 31427 18291 31433
rect 18506 31424 18512 31436
rect 18564 31424 18570 31476
rect 18874 31424 18880 31476
rect 18932 31464 18938 31476
rect 19150 31464 19156 31476
rect 18932 31436 19156 31464
rect 18932 31424 18938 31436
rect 19150 31424 19156 31436
rect 19208 31424 19214 31476
rect 21082 31464 21088 31476
rect 19812 31436 21088 31464
rect 14277 31399 14335 31405
rect 14277 31396 14289 31399
rect 13320 31368 14289 31396
rect 13320 31356 13326 31368
rect 14277 31365 14289 31368
rect 14323 31365 14335 31399
rect 14277 31359 14335 31365
rect 14829 31399 14887 31405
rect 14829 31365 14841 31399
rect 14875 31396 14887 31399
rect 15010 31396 15016 31408
rect 14875 31368 15016 31396
rect 14875 31365 14887 31368
rect 14829 31359 14887 31365
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31297 12311 31331
rect 12253 31291 12311 31297
rect 13173 31331 13231 31337
rect 13173 31297 13185 31331
rect 13219 31328 13231 31331
rect 13909 31331 13967 31337
rect 13909 31328 13921 31331
rect 13219 31300 13921 31328
rect 13219 31297 13231 31300
rect 13173 31291 13231 31297
rect 13909 31297 13921 31300
rect 13955 31297 13967 31331
rect 13909 31291 13967 31297
rect 14093 31331 14151 31337
rect 14093 31297 14105 31331
rect 14139 31328 14151 31331
rect 14844 31328 14872 31359
rect 15010 31356 15016 31368
rect 15068 31356 15074 31408
rect 17218 31356 17224 31408
rect 17276 31356 17282 31408
rect 17770 31356 17776 31408
rect 17828 31396 17834 31408
rect 17828 31368 19748 31396
rect 17828 31356 17834 31368
rect 14139 31300 14872 31328
rect 15749 31331 15807 31337
rect 14139 31297 14151 31300
rect 14093 31291 14151 31297
rect 15749 31297 15761 31331
rect 15795 31328 15807 31331
rect 15930 31328 15936 31340
rect 15795 31300 15936 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 15930 31288 15936 31300
rect 15988 31288 15994 31340
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 13357 31263 13415 31269
rect 13357 31229 13369 31263
rect 13403 31229 13415 31263
rect 13357 31223 13415 31229
rect 13372 31192 13400 31223
rect 15838 31220 15844 31272
rect 15896 31220 15902 31272
rect 16960 31260 16988 31291
rect 17034 31288 17040 31340
rect 17092 31288 17098 31340
rect 18230 31328 18236 31340
rect 18191 31300 18236 31328
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 18598 31288 18604 31340
rect 18656 31328 18662 31340
rect 19518 31328 19524 31340
rect 18656 31300 19524 31328
rect 18656 31288 18662 31300
rect 19518 31288 19524 31300
rect 19576 31288 19582 31340
rect 17678 31260 17684 31272
rect 16960 31232 17684 31260
rect 17678 31220 17684 31232
rect 17736 31260 17742 31272
rect 17736 31232 18092 31260
rect 17736 31220 17742 31232
rect 13446 31192 13452 31204
rect 13372 31164 13452 31192
rect 13446 31152 13452 31164
rect 13504 31192 13510 31204
rect 18064 31201 18092 31232
rect 18690 31220 18696 31272
rect 18748 31220 18754 31272
rect 18874 31220 18880 31272
rect 18932 31260 18938 31272
rect 19058 31260 19064 31272
rect 18932 31232 19064 31260
rect 18932 31220 18938 31232
rect 19058 31220 19064 31232
rect 19116 31260 19122 31272
rect 19720 31269 19748 31368
rect 19812 31337 19840 31436
rect 21082 31424 21088 31436
rect 21140 31424 21146 31476
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 26142 31464 26148 31476
rect 25096 31436 26148 31464
rect 25096 31424 25102 31436
rect 19978 31356 19984 31408
rect 20036 31396 20042 31408
rect 20254 31396 20260 31408
rect 20036 31368 20260 31396
rect 20036 31356 20042 31368
rect 20254 31356 20260 31368
rect 20312 31356 20318 31408
rect 20441 31399 20499 31405
rect 20441 31365 20453 31399
rect 20487 31365 20499 31399
rect 22370 31396 22376 31408
rect 20441 31359 20499 31365
rect 21468 31368 22376 31396
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 20456 31328 20484 31359
rect 19935 31300 20484 31328
rect 20717 31331 20775 31337
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 20717 31297 20729 31331
rect 20763 31297 20775 31331
rect 20717 31291 20775 31297
rect 19613 31263 19671 31269
rect 19613 31260 19625 31263
rect 19116 31232 19625 31260
rect 19116 31220 19122 31232
rect 19613 31229 19625 31232
rect 19659 31229 19671 31263
rect 19613 31223 19671 31229
rect 19705 31263 19763 31269
rect 19705 31229 19717 31263
rect 19751 31260 19763 31263
rect 19978 31260 19984 31272
rect 19751 31232 19984 31260
rect 19751 31229 19763 31232
rect 19705 31223 19763 31229
rect 18049 31195 18107 31201
rect 13504 31164 17356 31192
rect 13504 31152 13510 31164
rect 12713 31127 12771 31133
rect 12713 31093 12725 31127
rect 12759 31124 12771 31127
rect 12894 31124 12900 31136
rect 12759 31096 12900 31124
rect 12759 31093 12771 31096
rect 12713 31087 12771 31093
rect 12894 31084 12900 31096
rect 12952 31084 12958 31136
rect 17218 31084 17224 31136
rect 17276 31084 17282 31136
rect 17328 31124 17356 31164
rect 18049 31161 18061 31195
rect 18095 31161 18107 31195
rect 19628 31192 19656 31223
rect 19978 31220 19984 31232
rect 20036 31220 20042 31272
rect 20438 31220 20444 31272
rect 20496 31220 20502 31272
rect 20732 31260 20760 31291
rect 21358 31288 21364 31340
rect 21416 31288 21422 31340
rect 21468 31337 21496 31368
rect 22370 31356 22376 31368
rect 22428 31396 22434 31408
rect 23017 31399 23075 31405
rect 23017 31396 23029 31399
rect 22428 31368 23029 31396
rect 22428 31356 22434 31368
rect 23017 31365 23029 31368
rect 23063 31365 23075 31399
rect 23017 31359 23075 31365
rect 23934 31356 23940 31408
rect 23992 31396 23998 31408
rect 23992 31368 24348 31396
rect 23992 31356 23998 31368
rect 21453 31331 21511 31337
rect 21453 31297 21465 31331
rect 21499 31297 21511 31331
rect 21453 31291 21511 31297
rect 21910 31288 21916 31340
rect 21968 31328 21974 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21968 31300 22201 31328
rect 21968 31288 21974 31300
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22189 31291 22247 31297
rect 22278 31288 22284 31340
rect 22336 31288 22342 31340
rect 24320 31337 24348 31368
rect 24394 31356 24400 31408
rect 24452 31356 24458 31408
rect 24489 31399 24547 31405
rect 24489 31365 24501 31399
rect 24535 31396 24547 31399
rect 24762 31396 24768 31408
rect 24535 31368 24768 31396
rect 24535 31365 24547 31368
rect 24489 31359 24547 31365
rect 24762 31356 24768 31368
rect 24820 31356 24826 31408
rect 25424 31405 25452 31436
rect 26142 31424 26148 31436
rect 26200 31424 26206 31476
rect 37274 31464 37280 31476
rect 29196 31436 37280 31464
rect 25409 31399 25467 31405
rect 25409 31365 25421 31399
rect 25455 31396 25467 31399
rect 25455 31368 25489 31396
rect 25455 31365 25467 31368
rect 25409 31359 25467 31365
rect 25590 31356 25596 31408
rect 25648 31396 25654 31408
rect 26050 31396 26056 31408
rect 25648 31368 26056 31396
rect 25648 31356 25654 31368
rect 26050 31356 26056 31368
rect 26108 31356 26114 31408
rect 28626 31356 28632 31408
rect 28684 31396 28690 31408
rect 28684 31368 28948 31396
rect 28684 31356 28690 31368
rect 28920 31340 28948 31368
rect 22557 31331 22615 31337
rect 22557 31297 22569 31331
rect 22603 31297 22615 31331
rect 22557 31291 22615 31297
rect 23201 31331 23259 31337
rect 23201 31297 23213 31331
rect 23247 31328 23259 31331
rect 24305 31331 24363 31337
rect 23247 31300 24256 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 20806 31260 20812 31272
rect 20732 31232 20812 31260
rect 20806 31220 20812 31232
rect 20864 31260 20870 31272
rect 21177 31263 21235 31269
rect 21177 31260 21189 31263
rect 20864 31232 21189 31260
rect 20864 31220 20870 31232
rect 21177 31229 21189 31232
rect 21223 31260 21235 31263
rect 21266 31260 21272 31272
rect 21223 31232 21272 31260
rect 21223 31229 21235 31232
rect 21177 31223 21235 31229
rect 21266 31220 21272 31232
rect 21324 31220 21330 31272
rect 21634 31220 21640 31272
rect 21692 31260 21698 31272
rect 22572 31260 22600 31291
rect 22646 31260 22652 31272
rect 21692 31232 22652 31260
rect 21692 31220 21698 31232
rect 22646 31220 22652 31232
rect 22704 31220 22710 31272
rect 23106 31220 23112 31272
rect 23164 31260 23170 31272
rect 23382 31260 23388 31272
rect 23164 31232 23388 31260
rect 23164 31220 23170 31232
rect 23382 31220 23388 31232
rect 23440 31220 23446 31272
rect 23477 31263 23535 31269
rect 23477 31229 23489 31263
rect 23523 31260 23535 31263
rect 23566 31260 23572 31272
rect 23523 31232 23572 31260
rect 23523 31229 23535 31232
rect 23477 31223 23535 31229
rect 23566 31220 23572 31232
rect 23624 31220 23630 31272
rect 20622 31192 20628 31204
rect 18049 31155 18107 31161
rect 18156 31164 19564 31192
rect 19628 31164 20628 31192
rect 18156 31124 18184 31164
rect 17328 31096 18184 31124
rect 18601 31127 18659 31133
rect 18601 31093 18613 31127
rect 18647 31124 18659 31127
rect 19429 31127 19487 31133
rect 19429 31124 19441 31127
rect 18647 31096 19441 31124
rect 18647 31093 18659 31096
rect 18601 31087 18659 31093
rect 19429 31093 19441 31096
rect 19475 31093 19487 31127
rect 19536 31124 19564 31164
rect 20622 31152 20628 31164
rect 20680 31152 20686 31204
rect 22005 31195 22063 31201
rect 22005 31192 22017 31195
rect 20732 31164 22017 31192
rect 20732 31124 20760 31164
rect 22005 31161 22017 31164
rect 22051 31161 22063 31195
rect 22005 31155 22063 31161
rect 22465 31195 22523 31201
rect 22465 31161 22477 31195
rect 22511 31192 22523 31195
rect 22554 31192 22560 31204
rect 22511 31164 22560 31192
rect 22511 31161 22523 31164
rect 22465 31155 22523 31161
rect 22554 31152 22560 31164
rect 22612 31152 22618 31204
rect 24228 31192 24256 31300
rect 24305 31297 24317 31331
rect 24351 31328 24363 31331
rect 24578 31328 24584 31340
rect 24351 31300 24584 31328
rect 24351 31297 24363 31300
rect 24305 31291 24363 31297
rect 24578 31288 24584 31300
rect 24636 31288 24642 31340
rect 24670 31288 24676 31340
rect 24728 31288 24734 31340
rect 25038 31288 25044 31340
rect 25096 31328 25102 31340
rect 27709 31331 27767 31337
rect 27709 31328 27721 31331
rect 25096 31300 27721 31328
rect 25096 31288 25102 31300
rect 27709 31297 27721 31300
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 28813 31331 28871 31337
rect 28813 31297 28825 31331
rect 28859 31297 28871 31331
rect 28813 31291 28871 31297
rect 26142 31220 26148 31272
rect 26200 31220 26206 31272
rect 27985 31263 28043 31269
rect 27985 31229 27997 31263
rect 28031 31260 28043 31263
rect 28629 31263 28687 31269
rect 28629 31260 28641 31263
rect 28031 31232 28641 31260
rect 28031 31229 28043 31232
rect 27985 31223 28043 31229
rect 28629 31229 28641 31232
rect 28675 31229 28687 31263
rect 28828 31260 28856 31291
rect 28902 31288 28908 31340
rect 28960 31288 28966 31340
rect 29086 31288 29092 31340
rect 29144 31288 29150 31340
rect 29196 31337 29224 31436
rect 37274 31424 37280 31436
rect 37332 31424 37338 31476
rect 37384 31436 39988 31464
rect 29546 31356 29552 31408
rect 29604 31396 29610 31408
rect 30193 31399 30251 31405
rect 30193 31396 30205 31399
rect 29604 31368 30205 31396
rect 29604 31356 29610 31368
rect 30193 31365 30205 31368
rect 30239 31365 30251 31399
rect 30193 31359 30251 31365
rect 30282 31356 30288 31408
rect 30340 31356 30346 31408
rect 31205 31399 31263 31405
rect 30484 31368 31156 31396
rect 29181 31331 29239 31337
rect 29181 31297 29193 31331
rect 29227 31297 29239 31331
rect 29181 31291 29239 31297
rect 29914 31288 29920 31340
rect 29972 31328 29978 31340
rect 30484 31337 30512 31368
rect 30101 31331 30159 31337
rect 30101 31328 30113 31331
rect 29972 31300 30113 31328
rect 29972 31288 29978 31300
rect 30101 31297 30113 31300
rect 30147 31297 30159 31331
rect 30101 31291 30159 31297
rect 30469 31331 30527 31337
rect 30469 31297 30481 31331
rect 30515 31297 30527 31331
rect 30469 31291 30527 31297
rect 30926 31288 30932 31340
rect 30984 31288 30990 31340
rect 31021 31331 31079 31337
rect 31021 31297 31033 31331
rect 31067 31297 31079 31331
rect 31128 31328 31156 31368
rect 31205 31365 31217 31399
rect 31251 31396 31263 31399
rect 32398 31396 32404 31408
rect 31251 31368 32404 31396
rect 31251 31365 31263 31368
rect 31205 31359 31263 31365
rect 32398 31356 32404 31368
rect 32456 31356 32462 31408
rect 33226 31356 33232 31408
rect 33284 31396 33290 31408
rect 33962 31396 33968 31408
rect 33284 31368 33968 31396
rect 33284 31356 33290 31368
rect 33962 31356 33968 31368
rect 34020 31356 34026 31408
rect 34793 31399 34851 31405
rect 34793 31365 34805 31399
rect 34839 31396 34851 31399
rect 35526 31396 35532 31408
rect 34839 31368 35532 31396
rect 34839 31365 34851 31368
rect 34793 31359 34851 31365
rect 35526 31356 35532 31368
rect 35584 31356 35590 31408
rect 35986 31356 35992 31408
rect 36044 31396 36050 31408
rect 36044 31368 36860 31396
rect 36044 31356 36050 31368
rect 31570 31328 31576 31340
rect 31128 31300 31576 31328
rect 31021 31291 31079 31297
rect 30944 31260 30972 31288
rect 28828 31232 30972 31260
rect 31036 31260 31064 31291
rect 31570 31288 31576 31300
rect 31628 31288 31634 31340
rect 31665 31331 31723 31337
rect 31665 31297 31677 31331
rect 31711 31328 31723 31331
rect 31846 31328 31852 31340
rect 31711 31300 31852 31328
rect 31711 31297 31723 31300
rect 31665 31291 31723 31297
rect 31846 31288 31852 31300
rect 31904 31288 31910 31340
rect 32490 31288 32496 31340
rect 32548 31288 32554 31340
rect 32858 31288 32864 31340
rect 32916 31288 32922 31340
rect 34333 31331 34391 31337
rect 34333 31297 34345 31331
rect 34379 31328 34391 31331
rect 34698 31328 34704 31340
rect 34379 31300 34704 31328
rect 34379 31297 34391 31300
rect 34333 31291 34391 31297
rect 34698 31288 34704 31300
rect 34756 31328 34762 31340
rect 34885 31331 34943 31337
rect 34885 31328 34897 31331
rect 34756 31300 34897 31328
rect 34756 31288 34762 31300
rect 34885 31297 34897 31300
rect 34931 31328 34943 31331
rect 34974 31328 34980 31340
rect 34931 31300 34980 31328
rect 34931 31297 34943 31300
rect 34885 31291 34943 31297
rect 34974 31288 34980 31300
rect 35032 31288 35038 31340
rect 35069 31331 35127 31337
rect 35069 31297 35081 31331
rect 35115 31328 35127 31331
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 35115 31300 35817 31328
rect 35115 31297 35127 31300
rect 35069 31291 35127 31297
rect 35805 31297 35817 31300
rect 35851 31328 35863 31331
rect 35851 31300 36584 31328
rect 35851 31297 35863 31300
rect 35805 31291 35863 31297
rect 31754 31260 31760 31272
rect 31036 31232 31760 31260
rect 28629 31223 28687 31229
rect 31754 31220 31760 31232
rect 31812 31220 31818 31272
rect 33686 31220 33692 31272
rect 33744 31260 33750 31272
rect 35084 31260 35112 31291
rect 35710 31260 35716 31272
rect 33744 31232 35112 31260
rect 35176 31232 35716 31260
rect 33744 31220 33750 31232
rect 30374 31192 30380 31204
rect 24228 31164 30380 31192
rect 30374 31152 30380 31164
rect 30432 31152 30438 31204
rect 33594 31152 33600 31204
rect 33652 31192 33658 31204
rect 35176 31192 35204 31232
rect 35710 31220 35716 31232
rect 35768 31220 35774 31272
rect 35897 31263 35955 31269
rect 35897 31229 35909 31263
rect 35943 31229 35955 31263
rect 35897 31223 35955 31229
rect 35989 31263 36047 31269
rect 35989 31229 36001 31263
rect 36035 31260 36047 31263
rect 36446 31260 36452 31272
rect 36035 31232 36452 31260
rect 36035 31229 36047 31232
rect 35989 31223 36047 31229
rect 35912 31192 35940 31223
rect 36446 31220 36452 31232
rect 36504 31220 36510 31272
rect 36556 31260 36584 31300
rect 36630 31288 36636 31340
rect 36688 31288 36694 31340
rect 36832 31337 36860 31368
rect 36998 31356 37004 31408
rect 37056 31396 37062 31408
rect 37384 31396 37412 31436
rect 37056 31368 37412 31396
rect 37056 31356 37062 31368
rect 38746 31356 38752 31408
rect 38804 31356 38810 31408
rect 36817 31331 36875 31337
rect 36817 31297 36829 31331
rect 36863 31328 36875 31331
rect 37461 31331 37519 31337
rect 37461 31328 37473 31331
rect 36863 31300 37473 31328
rect 36863 31297 36875 31300
rect 36817 31291 36875 31297
rect 37461 31297 37473 31300
rect 37507 31297 37519 31331
rect 37461 31291 37519 31297
rect 38286 31288 38292 31340
rect 38344 31328 38350 31340
rect 38565 31331 38623 31337
rect 38565 31328 38577 31331
rect 38344 31300 38577 31328
rect 38344 31288 38350 31300
rect 38565 31297 38577 31300
rect 38611 31297 38623 31331
rect 38565 31291 38623 31297
rect 39114 31288 39120 31340
rect 39172 31328 39178 31340
rect 39209 31331 39267 31337
rect 39209 31328 39221 31331
rect 39172 31300 39221 31328
rect 39172 31288 39178 31300
rect 39209 31297 39221 31300
rect 39255 31297 39267 31331
rect 39209 31291 39267 31297
rect 37366 31260 37372 31272
rect 36556 31232 37372 31260
rect 37366 31220 37372 31232
rect 37424 31220 37430 31272
rect 38378 31260 38384 31272
rect 37844 31232 38384 31260
rect 33652 31164 35204 31192
rect 35728 31164 35940 31192
rect 33652 31152 33658 31164
rect 35728 31136 35756 31164
rect 36078 31152 36084 31204
rect 36136 31192 36142 31204
rect 36136 31164 36768 31192
rect 36136 31152 36142 31164
rect 36740 31136 36768 31164
rect 37274 31152 37280 31204
rect 37332 31192 37338 31204
rect 37844 31201 37872 31232
rect 38378 31220 38384 31232
rect 38436 31220 38442 31272
rect 39224 31260 39252 31291
rect 39390 31288 39396 31340
rect 39448 31288 39454 31340
rect 39960 31328 39988 31436
rect 41874 31424 41880 31476
rect 41932 31424 41938 31476
rect 40034 31356 40040 31408
rect 40092 31396 40098 31408
rect 40310 31396 40316 31408
rect 40092 31368 40316 31396
rect 40092 31356 40098 31368
rect 40310 31356 40316 31368
rect 40368 31396 40374 31408
rect 41049 31399 41107 31405
rect 41049 31396 41061 31399
rect 40368 31368 41061 31396
rect 40368 31356 40374 31368
rect 41049 31365 41061 31368
rect 41095 31365 41107 31399
rect 41049 31359 41107 31365
rect 40405 31331 40463 31337
rect 40405 31328 40417 31331
rect 39960 31300 40417 31328
rect 40405 31297 40417 31300
rect 40451 31328 40463 31331
rect 40494 31328 40500 31340
rect 40451 31300 40500 31328
rect 40451 31297 40463 31300
rect 40405 31291 40463 31297
rect 40494 31288 40500 31300
rect 40552 31288 40558 31340
rect 40954 31288 40960 31340
rect 41012 31328 41018 31340
rect 41233 31331 41291 31337
rect 41233 31328 41245 31331
rect 41012 31300 41245 31328
rect 41012 31288 41018 31300
rect 41233 31297 41245 31300
rect 41279 31297 41291 31331
rect 41233 31291 41291 31297
rect 41322 31288 41328 31340
rect 41380 31288 41386 31340
rect 41414 31288 41420 31340
rect 41472 31328 41478 31340
rect 42061 31331 42119 31337
rect 42061 31328 42073 31331
rect 41472 31300 42073 31328
rect 41472 31288 41478 31300
rect 42061 31297 42073 31300
rect 42107 31328 42119 31331
rect 42886 31328 42892 31340
rect 42107 31300 42892 31328
rect 42107 31297 42119 31300
rect 42061 31291 42119 31297
rect 42886 31288 42892 31300
rect 42944 31328 42950 31340
rect 43073 31331 43131 31337
rect 43073 31328 43085 31331
rect 42944 31300 43085 31328
rect 42944 31288 42950 31300
rect 43073 31297 43085 31300
rect 43119 31297 43131 31331
rect 43073 31291 43131 31297
rect 39574 31260 39580 31272
rect 39224 31232 39580 31260
rect 39574 31220 39580 31232
rect 39632 31220 39638 31272
rect 40589 31263 40647 31269
rect 40589 31229 40601 31263
rect 40635 31260 40647 31263
rect 41690 31260 41696 31272
rect 40635 31232 41696 31260
rect 40635 31229 40647 31232
rect 40589 31223 40647 31229
rect 41690 31220 41696 31232
rect 41748 31220 41754 31272
rect 42702 31220 42708 31272
rect 42760 31260 42766 31272
rect 43990 31260 43996 31272
rect 42760 31232 43996 31260
rect 42760 31220 42766 31232
rect 43990 31220 43996 31232
rect 44048 31220 44054 31272
rect 37829 31195 37887 31201
rect 37829 31192 37841 31195
rect 37332 31164 37841 31192
rect 37332 31152 37338 31164
rect 37829 31161 37841 31164
rect 37875 31161 37887 31195
rect 37829 31155 37887 31161
rect 38102 31152 38108 31204
rect 38160 31192 38166 31204
rect 40034 31192 40040 31204
rect 38160 31164 40040 31192
rect 38160 31152 38166 31164
rect 40034 31152 40040 31164
rect 40092 31152 40098 31204
rect 40126 31152 40132 31204
rect 40184 31192 40190 31204
rect 41049 31195 41107 31201
rect 41049 31192 41061 31195
rect 40184 31164 41061 31192
rect 40184 31152 40190 31164
rect 41049 31161 41061 31164
rect 41095 31161 41107 31195
rect 41049 31155 41107 31161
rect 19536 31096 20760 31124
rect 21269 31127 21327 31133
rect 19429 31087 19487 31093
rect 21269 31093 21281 31127
rect 21315 31124 21327 31127
rect 21634 31124 21640 31136
rect 21315 31096 21640 31124
rect 21315 31093 21327 31096
rect 21269 31087 21327 31093
rect 21634 31084 21640 31096
rect 21692 31084 21698 31136
rect 24026 31084 24032 31136
rect 24084 31124 24090 31136
rect 24121 31127 24179 31133
rect 24121 31124 24133 31127
rect 24084 31096 24133 31124
rect 24084 31084 24090 31096
rect 24121 31093 24133 31096
rect 24167 31093 24179 31127
rect 24121 31087 24179 31093
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 29730 31124 29736 31136
rect 25004 31096 29736 31124
rect 25004 31084 25010 31096
rect 29730 31084 29736 31096
rect 29788 31084 29794 31136
rect 29914 31084 29920 31136
rect 29972 31084 29978 31136
rect 30006 31084 30012 31136
rect 30064 31124 30070 31136
rect 31205 31127 31263 31133
rect 31205 31124 31217 31127
rect 30064 31096 31217 31124
rect 30064 31084 30070 31096
rect 31205 31093 31217 31096
rect 31251 31093 31263 31127
rect 31205 31087 31263 31093
rect 32306 31084 32312 31136
rect 32364 31084 32370 31136
rect 32766 31084 32772 31136
rect 32824 31084 32830 31136
rect 33318 31084 33324 31136
rect 33376 31084 33382 31136
rect 35710 31084 35716 31136
rect 35768 31084 35774 31136
rect 36173 31127 36231 31133
rect 36173 31093 36185 31127
rect 36219 31124 36231 31127
rect 36262 31124 36268 31136
rect 36219 31096 36268 31124
rect 36219 31093 36231 31096
rect 36173 31087 36231 31093
rect 36262 31084 36268 31096
rect 36320 31084 36326 31136
rect 36722 31084 36728 31136
rect 36780 31084 36786 31136
rect 37642 31084 37648 31136
rect 37700 31124 37706 31136
rect 37921 31127 37979 31133
rect 37921 31124 37933 31127
rect 37700 31096 37933 31124
rect 37700 31084 37706 31096
rect 37921 31093 37933 31096
rect 37967 31093 37979 31127
rect 37921 31087 37979 31093
rect 38378 31084 38384 31136
rect 38436 31084 38442 31136
rect 39206 31084 39212 31136
rect 39264 31124 39270 31136
rect 39301 31127 39359 31133
rect 39301 31124 39313 31127
rect 39264 31096 39313 31124
rect 39264 31084 39270 31096
rect 39301 31093 39313 31096
rect 39347 31093 39359 31127
rect 39301 31087 39359 31093
rect 40218 31084 40224 31136
rect 40276 31124 40282 31136
rect 40862 31124 40868 31136
rect 40276 31096 40868 31124
rect 40276 31084 40282 31096
rect 40862 31084 40868 31096
rect 40920 31084 40926 31136
rect 41966 31084 41972 31136
rect 42024 31124 42030 31136
rect 42613 31127 42671 31133
rect 42613 31124 42625 31127
rect 42024 31096 42625 31124
rect 42024 31084 42030 31096
rect 42613 31093 42625 31096
rect 42659 31093 42671 31127
rect 42613 31087 42671 31093
rect 42794 31084 42800 31136
rect 42852 31124 42858 31136
rect 42981 31127 43039 31133
rect 42981 31124 42993 31127
rect 42852 31096 42993 31124
rect 42852 31084 42858 31096
rect 42981 31093 42993 31096
rect 43027 31124 43039 31127
rect 43254 31124 43260 31136
rect 43027 31096 43260 31124
rect 43027 31093 43039 31096
rect 42981 31087 43039 31093
rect 43254 31084 43260 31096
rect 43312 31084 43318 31136
rect 1104 31034 43884 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 43884 31034
rect 1104 30960 43884 30982
rect 12618 30880 12624 30932
rect 12676 30920 12682 30932
rect 12713 30923 12771 30929
rect 12713 30920 12725 30923
rect 12676 30892 12725 30920
rect 12676 30880 12682 30892
rect 12713 30889 12725 30892
rect 12759 30889 12771 30923
rect 12713 30883 12771 30889
rect 13173 30923 13231 30929
rect 13173 30889 13185 30923
rect 13219 30920 13231 30923
rect 13262 30920 13268 30932
rect 13219 30892 13268 30920
rect 13219 30889 13231 30892
rect 13173 30883 13231 30889
rect 13262 30880 13268 30892
rect 13320 30880 13326 30932
rect 14369 30923 14427 30929
rect 14369 30889 14381 30923
rect 14415 30920 14427 30923
rect 15010 30920 15016 30932
rect 14415 30892 15016 30920
rect 14415 30889 14427 30892
rect 14369 30883 14427 30889
rect 11882 30812 11888 30864
rect 11940 30852 11946 30864
rect 14384 30852 14412 30883
rect 15010 30880 15016 30892
rect 15068 30880 15074 30932
rect 18138 30880 18144 30932
rect 18196 30880 18202 30932
rect 18601 30923 18659 30929
rect 18601 30889 18613 30923
rect 18647 30920 18659 30923
rect 18690 30920 18696 30932
rect 18647 30892 18696 30920
rect 18647 30889 18659 30892
rect 18601 30883 18659 30889
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 18782 30880 18788 30932
rect 18840 30920 18846 30932
rect 20622 30920 20628 30932
rect 18840 30892 20628 30920
rect 18840 30880 18846 30892
rect 20622 30880 20628 30892
rect 20680 30880 20686 30932
rect 20714 30880 20720 30932
rect 20772 30920 20778 30932
rect 22094 30920 22100 30932
rect 20772 30892 22100 30920
rect 20772 30880 20778 30892
rect 22094 30880 22100 30892
rect 22152 30880 22158 30932
rect 23382 30880 23388 30932
rect 23440 30920 23446 30932
rect 23661 30923 23719 30929
rect 23661 30920 23673 30923
rect 23440 30892 23673 30920
rect 23440 30880 23446 30892
rect 23661 30889 23673 30892
rect 23707 30889 23719 30923
rect 23661 30883 23719 30889
rect 28902 30880 28908 30932
rect 28960 30920 28966 30932
rect 29730 30920 29736 30932
rect 28960 30892 29736 30920
rect 28960 30880 28966 30892
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 30926 30880 30932 30932
rect 30984 30920 30990 30932
rect 31297 30923 31355 30929
rect 31297 30920 31309 30923
rect 30984 30892 31309 30920
rect 30984 30880 30990 30892
rect 31297 30889 31309 30892
rect 31343 30889 31355 30923
rect 31297 30883 31355 30889
rect 33045 30923 33103 30929
rect 33045 30889 33057 30923
rect 33091 30920 33103 30923
rect 33778 30920 33784 30932
rect 33091 30892 33784 30920
rect 33091 30889 33103 30892
rect 33045 30883 33103 30889
rect 33778 30880 33784 30892
rect 33836 30880 33842 30932
rect 35802 30880 35808 30932
rect 35860 30920 35866 30932
rect 36630 30920 36636 30932
rect 35860 30892 36636 30920
rect 35860 30880 35866 30892
rect 36630 30880 36636 30892
rect 36688 30880 36694 30932
rect 36814 30880 36820 30932
rect 36872 30920 36878 30932
rect 37001 30923 37059 30929
rect 37001 30920 37013 30923
rect 36872 30892 37013 30920
rect 36872 30880 36878 30892
rect 37001 30889 37013 30892
rect 37047 30889 37059 30923
rect 37001 30883 37059 30889
rect 37550 30880 37556 30932
rect 37608 30880 37614 30932
rect 37734 30880 37740 30932
rect 37792 30920 37798 30932
rect 38013 30923 38071 30929
rect 38013 30920 38025 30923
rect 37792 30892 38025 30920
rect 37792 30880 37798 30892
rect 38013 30889 38025 30892
rect 38059 30889 38071 30923
rect 38013 30883 38071 30889
rect 38197 30923 38255 30929
rect 38197 30889 38209 30923
rect 38243 30889 38255 30923
rect 38197 30883 38255 30889
rect 20990 30852 20996 30864
rect 11940 30824 14412 30852
rect 16132 30824 20996 30852
rect 11940 30812 11946 30824
rect 16132 30793 16160 30824
rect 20990 30812 20996 30824
rect 21048 30812 21054 30864
rect 21358 30812 21364 30864
rect 21416 30812 21422 30864
rect 21910 30812 21916 30864
rect 21968 30812 21974 30864
rect 22281 30855 22339 30861
rect 22281 30821 22293 30855
rect 22327 30852 22339 30855
rect 23109 30855 23167 30861
rect 23109 30852 23121 30855
rect 22327 30824 23121 30852
rect 22327 30821 22339 30824
rect 22281 30815 22339 30821
rect 23109 30821 23121 30824
rect 23155 30821 23167 30855
rect 23109 30815 23167 30821
rect 26050 30812 26056 30864
rect 26108 30852 26114 30864
rect 27614 30852 27620 30864
rect 26108 30824 27620 30852
rect 26108 30812 26114 30824
rect 27614 30812 27620 30824
rect 27672 30812 27678 30864
rect 28994 30852 29000 30864
rect 27724 30824 29000 30852
rect 16117 30787 16175 30793
rect 16117 30753 16129 30787
rect 16163 30753 16175 30787
rect 16117 30747 16175 30753
rect 18414 30744 18420 30796
rect 18472 30784 18478 30796
rect 19426 30784 19432 30796
rect 18472 30756 19432 30784
rect 18472 30744 18478 30756
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 20438 30784 20444 30796
rect 19628 30756 20444 30784
rect 12894 30676 12900 30728
rect 12952 30676 12958 30728
rect 12986 30676 12992 30728
rect 13044 30676 13050 30728
rect 13265 30719 13323 30725
rect 13265 30685 13277 30719
rect 13311 30716 13323 30719
rect 13446 30716 13452 30728
rect 13311 30688 13452 30716
rect 13311 30685 13323 30688
rect 13265 30679 13323 30685
rect 13446 30676 13452 30688
rect 13504 30676 13510 30728
rect 15838 30676 15844 30728
rect 15896 30716 15902 30728
rect 15896 30688 18828 30716
rect 15896 30676 15902 30688
rect 17770 30608 17776 30660
rect 17828 30648 17834 30660
rect 18601 30651 18659 30657
rect 18601 30648 18613 30651
rect 17828 30620 18613 30648
rect 17828 30608 17834 30620
rect 18601 30617 18613 30620
rect 18647 30617 18659 30651
rect 18800 30648 18828 30688
rect 18874 30676 18880 30728
rect 18932 30676 18938 30728
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19628 30725 19656 30756
rect 20438 30744 20444 30756
rect 20496 30784 20502 30796
rect 24765 30787 24823 30793
rect 24765 30784 24777 30787
rect 20496 30756 24777 30784
rect 20496 30744 20502 30756
rect 24765 30753 24777 30756
rect 24811 30753 24823 30787
rect 24765 30747 24823 30753
rect 19613 30719 19671 30725
rect 19613 30716 19625 30719
rect 19392 30688 19625 30716
rect 19392 30676 19398 30688
rect 19613 30685 19625 30688
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19702 30676 19708 30728
rect 19760 30676 19766 30728
rect 19886 30676 19892 30728
rect 19944 30676 19950 30728
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30716 20039 30719
rect 21082 30716 21088 30728
rect 20027 30688 21088 30716
rect 20027 30685 20039 30688
rect 19981 30679 20039 30685
rect 21082 30676 21088 30688
rect 21140 30676 21146 30728
rect 21174 30676 21180 30728
rect 21232 30716 21238 30728
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 21232 30688 21281 30716
rect 21232 30676 21238 30688
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 21453 30719 21511 30725
rect 21453 30685 21465 30719
rect 21499 30685 21511 30719
rect 21453 30679 21511 30685
rect 21468 30648 21496 30679
rect 21634 30676 21640 30728
rect 21692 30716 21698 30728
rect 22097 30719 22155 30725
rect 22097 30716 22109 30719
rect 21692 30688 22109 30716
rect 21692 30676 21698 30688
rect 22097 30685 22109 30688
rect 22143 30685 22155 30719
rect 22097 30679 22155 30685
rect 22370 30676 22376 30728
rect 22428 30676 22434 30728
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30716 23075 30719
rect 23106 30716 23112 30728
rect 23063 30688 23112 30716
rect 23063 30685 23075 30688
rect 23017 30679 23075 30685
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30716 23259 30719
rect 23750 30716 23756 30728
rect 23247 30688 23756 30716
rect 23247 30685 23259 30688
rect 23201 30679 23259 30685
rect 23216 30648 23244 30679
rect 23750 30676 23756 30688
rect 23808 30676 23814 30728
rect 24946 30676 24952 30728
rect 25004 30676 25010 30728
rect 25222 30676 25228 30728
rect 25280 30716 25286 30728
rect 25409 30719 25467 30725
rect 25409 30716 25421 30719
rect 25280 30688 25421 30716
rect 25280 30676 25286 30688
rect 25409 30685 25421 30688
rect 25455 30716 25467 30719
rect 25590 30716 25596 30728
rect 25455 30688 25596 30716
rect 25455 30685 25467 30688
rect 25409 30679 25467 30685
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 25685 30719 25743 30725
rect 25685 30685 25697 30719
rect 25731 30716 25743 30719
rect 25774 30716 25780 30728
rect 25731 30688 25780 30716
rect 25731 30685 25743 30688
rect 25685 30679 25743 30685
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 25866 30676 25872 30728
rect 25924 30676 25930 30728
rect 27617 30719 27675 30725
rect 27617 30685 27629 30719
rect 27663 30716 27675 30719
rect 27724 30716 27752 30824
rect 28994 30812 29000 30824
rect 29052 30812 29058 30864
rect 30190 30812 30196 30864
rect 30248 30852 30254 30864
rect 32493 30855 32551 30861
rect 32493 30852 32505 30855
rect 30248 30824 32505 30852
rect 30248 30812 30254 30824
rect 32493 30821 32505 30824
rect 32539 30821 32551 30855
rect 38212 30852 38240 30883
rect 38470 30880 38476 30932
rect 38528 30920 38534 30932
rect 39485 30923 39543 30929
rect 39485 30920 39497 30923
rect 38528 30892 39497 30920
rect 38528 30880 38534 30892
rect 39485 30889 39497 30892
rect 39531 30889 39543 30923
rect 39485 30883 39543 30889
rect 40126 30880 40132 30932
rect 40184 30880 40190 30932
rect 40954 30852 40960 30864
rect 32493 30815 32551 30821
rect 34164 30824 40960 30852
rect 34164 30796 34192 30824
rect 40954 30812 40960 30824
rect 41012 30812 41018 30864
rect 28810 30784 28816 30796
rect 28000 30756 28816 30784
rect 27663 30688 27752 30716
rect 27663 30685 27675 30688
rect 27617 30679 27675 30685
rect 27890 30676 27896 30728
rect 27948 30676 27954 30728
rect 28000 30725 28028 30756
rect 28810 30744 28816 30756
rect 28868 30744 28874 30796
rect 30742 30744 30748 30796
rect 30800 30784 30806 30796
rect 31846 30784 31852 30796
rect 30800 30756 31852 30784
rect 30800 30744 30806 30756
rect 31846 30744 31852 30756
rect 31904 30744 31910 30796
rect 33689 30787 33747 30793
rect 33689 30784 33701 30787
rect 32692 30756 33701 30784
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 28261 30719 28319 30725
rect 28261 30685 28273 30719
rect 28307 30685 28319 30719
rect 28261 30679 28319 30685
rect 18800 30620 23244 30648
rect 24964 30648 24992 30676
rect 26697 30651 26755 30657
rect 26697 30648 26709 30651
rect 24964 30620 26709 30648
rect 18601 30611 18659 30617
rect 26697 30617 26709 30620
rect 26743 30648 26755 30651
rect 27338 30648 27344 30660
rect 26743 30620 27344 30648
rect 26743 30617 26755 30620
rect 26697 30611 26755 30617
rect 27338 30608 27344 30620
rect 27396 30608 27402 30660
rect 28276 30648 28304 30679
rect 28442 30676 28448 30728
rect 28500 30676 28506 30728
rect 29914 30676 29920 30728
rect 29972 30676 29978 30728
rect 30193 30719 30251 30725
rect 30193 30685 30205 30719
rect 30239 30716 30251 30719
rect 30926 30716 30932 30728
rect 30239 30688 30932 30716
rect 30239 30685 30251 30688
rect 30193 30679 30251 30685
rect 30926 30676 30932 30688
rect 30984 30676 30990 30728
rect 31389 30719 31447 30725
rect 31389 30685 31401 30719
rect 31435 30716 31447 30719
rect 32306 30716 32312 30728
rect 31435 30688 32312 30716
rect 31435 30685 31447 30688
rect 31389 30679 31447 30685
rect 32306 30676 32312 30688
rect 32364 30676 32370 30728
rect 32582 30676 32588 30728
rect 32640 30716 32646 30728
rect 32692 30725 32720 30756
rect 33689 30753 33701 30756
rect 33735 30753 33747 30787
rect 33689 30747 33747 30753
rect 34146 30744 34152 30796
rect 34204 30744 34210 30796
rect 36538 30744 36544 30796
rect 36596 30784 36602 30796
rect 41230 30784 41236 30796
rect 36596 30756 38516 30784
rect 36596 30744 36602 30756
rect 32677 30719 32735 30725
rect 32677 30716 32689 30719
rect 32640 30688 32689 30716
rect 32640 30676 32646 30688
rect 32677 30685 32689 30688
rect 32723 30685 32735 30719
rect 32677 30679 32735 30685
rect 32766 30676 32772 30728
rect 32824 30676 32830 30728
rect 33594 30676 33600 30728
rect 33652 30676 33658 30728
rect 33965 30719 34023 30725
rect 33965 30685 33977 30719
rect 34011 30716 34023 30719
rect 34422 30716 34428 30728
rect 34011 30688 34428 30716
rect 34011 30685 34023 30688
rect 33965 30679 34023 30685
rect 34422 30676 34428 30688
rect 34480 30676 34486 30728
rect 34698 30676 34704 30728
rect 34756 30716 34762 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34756 30688 34897 30716
rect 34756 30676 34762 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35434 30676 35440 30728
rect 35492 30676 35498 30728
rect 35618 30676 35624 30728
rect 35676 30676 35682 30728
rect 36262 30676 36268 30728
rect 36320 30676 36326 30728
rect 36449 30719 36507 30725
rect 36449 30685 36461 30719
rect 36495 30685 36507 30719
rect 36449 30679 36507 30685
rect 37185 30719 37243 30725
rect 37185 30685 37197 30719
rect 37231 30716 37243 30719
rect 37274 30716 37280 30728
rect 37231 30688 37280 30716
rect 37231 30685 37243 30688
rect 37185 30679 37243 30685
rect 30282 30648 30288 30660
rect 28276 30620 30288 30648
rect 30282 30608 30288 30620
rect 30340 30608 30346 30660
rect 32858 30608 32864 30660
rect 32916 30648 32922 30660
rect 33137 30651 33195 30657
rect 33137 30648 33149 30651
rect 32916 30620 33149 30648
rect 32916 30608 32922 30620
rect 33137 30617 33149 30620
rect 33183 30648 33195 30651
rect 36081 30651 36139 30657
rect 36081 30648 36093 30651
rect 33183 30620 36093 30648
rect 33183 30617 33195 30620
rect 33137 30611 33195 30617
rect 36081 30617 36093 30620
rect 36127 30617 36139 30651
rect 36464 30648 36492 30679
rect 37274 30676 37280 30688
rect 37332 30676 37338 30728
rect 37369 30719 37427 30725
rect 37369 30685 37381 30719
rect 37415 30716 37427 30719
rect 38102 30716 38108 30728
rect 37415 30688 38108 30716
rect 37415 30685 37427 30688
rect 37369 30679 37427 30685
rect 38102 30676 38108 30688
rect 38160 30676 38166 30728
rect 36630 30648 36636 30660
rect 36464 30620 36636 30648
rect 36081 30611 36139 30617
rect 36630 30608 36636 30620
rect 36688 30648 36694 30660
rect 36909 30651 36967 30657
rect 36909 30648 36921 30651
rect 36688 30620 36921 30648
rect 36688 30608 36694 30620
rect 36909 30617 36921 30620
rect 36955 30617 36967 30651
rect 38381 30651 38439 30657
rect 38381 30648 38393 30651
rect 36909 30611 36967 30617
rect 37384 30620 38393 30648
rect 37384 30592 37412 30620
rect 38381 30617 38393 30620
rect 38427 30617 38439 30651
rect 38488 30648 38516 30756
rect 39500 30756 41236 30784
rect 39301 30719 39359 30725
rect 39301 30685 39313 30719
rect 39347 30716 39359 30719
rect 39390 30716 39396 30728
rect 39347 30688 39396 30716
rect 39347 30685 39359 30688
rect 39301 30679 39359 30685
rect 39390 30676 39396 30688
rect 39448 30676 39454 30728
rect 39500 30725 39528 30756
rect 41230 30744 41236 30756
rect 41288 30744 41294 30796
rect 42521 30787 42579 30793
rect 42521 30753 42533 30787
rect 42567 30784 42579 30787
rect 42702 30784 42708 30796
rect 42567 30756 42708 30784
rect 42567 30753 42579 30756
rect 42521 30747 42579 30753
rect 42702 30744 42708 30756
rect 42760 30744 42766 30796
rect 42794 30744 42800 30796
rect 42852 30744 42858 30796
rect 39485 30719 39543 30725
rect 39485 30685 39497 30719
rect 39531 30685 39543 30719
rect 39485 30679 39543 30685
rect 39850 30676 39856 30728
rect 39908 30716 39914 30728
rect 40037 30719 40095 30725
rect 40037 30716 40049 30719
rect 39908 30688 40049 30716
rect 39908 30676 39914 30688
rect 40037 30685 40049 30688
rect 40083 30685 40095 30719
rect 40037 30679 40095 30685
rect 40218 30676 40224 30728
rect 40276 30676 40282 30728
rect 40678 30676 40684 30728
rect 40736 30676 40742 30728
rect 40862 30676 40868 30728
rect 40920 30676 40926 30728
rect 41966 30676 41972 30728
rect 42024 30676 42030 30728
rect 40773 30651 40831 30657
rect 40773 30648 40785 30651
rect 38488 30620 40785 30648
rect 38381 30611 38439 30617
rect 40773 30617 40785 30620
rect 40819 30617 40831 30651
rect 40773 30611 40831 30617
rect 11974 30540 11980 30592
rect 12032 30580 12038 30592
rect 13906 30580 13912 30592
rect 12032 30552 13912 30580
rect 12032 30540 12038 30552
rect 13906 30540 13912 30552
rect 13964 30580 13970 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 13964 30552 15485 30580
rect 13964 30540 13970 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 15473 30543 15531 30549
rect 15654 30540 15660 30592
rect 15712 30580 15718 30592
rect 15841 30583 15899 30589
rect 15841 30580 15853 30583
rect 15712 30552 15853 30580
rect 15712 30540 15718 30552
rect 15841 30549 15853 30552
rect 15887 30549 15899 30583
rect 15841 30543 15899 30549
rect 15930 30540 15936 30592
rect 15988 30540 15994 30592
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 17313 30583 17371 30589
rect 17313 30580 17325 30583
rect 17000 30552 17325 30580
rect 17000 30540 17006 30552
rect 17313 30549 17325 30552
rect 17359 30549 17371 30583
rect 17313 30543 17371 30549
rect 18785 30583 18843 30589
rect 18785 30549 18797 30583
rect 18831 30580 18843 30583
rect 19150 30580 19156 30592
rect 18831 30552 19156 30580
rect 18831 30549 18843 30552
rect 18785 30543 18843 30549
rect 19150 30540 19156 30552
rect 19208 30540 19214 30592
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 19702 30540 19708 30592
rect 19760 30580 19766 30592
rect 20070 30580 20076 30592
rect 19760 30552 20076 30580
rect 19760 30540 19766 30552
rect 20070 30540 20076 30552
rect 20128 30580 20134 30592
rect 20530 30580 20536 30592
rect 20128 30552 20536 30580
rect 20128 30540 20134 30552
rect 20530 30540 20536 30552
rect 20588 30580 20594 30592
rect 23106 30580 23112 30592
rect 20588 30552 23112 30580
rect 20588 30540 20594 30552
rect 23106 30540 23112 30552
rect 23164 30580 23170 30592
rect 25130 30580 25136 30592
rect 23164 30552 25136 30580
rect 23164 30540 23170 30552
rect 25130 30540 25136 30552
rect 25188 30540 25194 30592
rect 27246 30540 27252 30592
rect 27304 30540 27310 30592
rect 28902 30540 28908 30592
rect 28960 30580 28966 30592
rect 29089 30583 29147 30589
rect 29089 30580 29101 30583
rect 28960 30552 29101 30580
rect 28960 30540 28966 30552
rect 29089 30549 29101 30552
rect 29135 30549 29147 30583
rect 29089 30543 29147 30549
rect 29178 30540 29184 30592
rect 29236 30580 29242 30592
rect 29733 30583 29791 30589
rect 29733 30580 29745 30583
rect 29236 30552 29745 30580
rect 29236 30540 29242 30552
rect 29733 30549 29745 30552
rect 29779 30549 29791 30583
rect 29733 30543 29791 30549
rect 29914 30540 29920 30592
rect 29972 30580 29978 30592
rect 30101 30583 30159 30589
rect 30101 30580 30113 30583
rect 29972 30552 30113 30580
rect 29972 30540 29978 30552
rect 30101 30549 30113 30552
rect 30147 30580 30159 30583
rect 30650 30580 30656 30592
rect 30147 30552 30656 30580
rect 30147 30549 30159 30552
rect 30101 30543 30159 30549
rect 30650 30540 30656 30552
rect 30708 30540 30714 30592
rect 31938 30540 31944 30592
rect 31996 30540 32002 30592
rect 37366 30540 37372 30592
rect 37424 30540 37430 30592
rect 38181 30583 38239 30589
rect 38181 30549 38193 30583
rect 38227 30580 38239 30583
rect 38562 30580 38568 30592
rect 38227 30552 38568 30580
rect 38227 30549 38239 30552
rect 38181 30543 38239 30549
rect 38562 30540 38568 30552
rect 38620 30540 38626 30592
rect 38838 30540 38844 30592
rect 38896 30580 38902 30592
rect 41322 30580 41328 30592
rect 38896 30552 41328 30580
rect 38896 30540 38902 30552
rect 41322 30540 41328 30552
rect 41380 30540 41386 30592
rect 41690 30540 41696 30592
rect 41748 30540 41754 30592
rect 1104 30490 43884 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 43884 30490
rect 1104 30416 43884 30438
rect 17954 30336 17960 30388
rect 18012 30376 18018 30388
rect 18325 30379 18383 30385
rect 18325 30376 18337 30379
rect 18012 30348 18337 30376
rect 18012 30336 18018 30348
rect 18325 30345 18337 30348
rect 18371 30345 18383 30379
rect 19978 30376 19984 30388
rect 18325 30339 18383 30345
rect 19260 30348 19984 30376
rect 12894 30308 12900 30320
rect 12084 30280 12900 30308
rect 12084 30249 12112 30280
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 16482 30308 16488 30320
rect 15120 30280 16488 30308
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30209 12127 30243
rect 12069 30203 12127 30209
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30240 12311 30243
rect 12986 30240 12992 30252
rect 12299 30212 12992 30240
rect 12299 30209 12311 30212
rect 12253 30203 12311 30209
rect 12986 30200 12992 30212
rect 13044 30200 13050 30252
rect 15120 30240 15148 30280
rect 16482 30268 16488 30280
rect 16540 30268 16546 30320
rect 18046 30268 18052 30320
rect 18104 30308 18110 30320
rect 18233 30311 18291 30317
rect 18233 30308 18245 30311
rect 18104 30280 18245 30308
rect 18104 30268 18110 30280
rect 18233 30277 18245 30280
rect 18279 30308 18291 30311
rect 18782 30308 18788 30320
rect 18279 30280 18788 30308
rect 18279 30277 18291 30280
rect 18233 30271 18291 30277
rect 18782 30268 18788 30280
rect 18840 30268 18846 30320
rect 19260 30308 19288 30348
rect 19978 30336 19984 30348
rect 20036 30336 20042 30388
rect 20622 30336 20628 30388
rect 20680 30376 20686 30388
rect 27246 30376 27252 30388
rect 20680 30348 27252 30376
rect 20680 30336 20686 30348
rect 27246 30336 27252 30348
rect 27304 30336 27310 30388
rect 27338 30336 27344 30388
rect 27396 30376 27402 30388
rect 31846 30376 31852 30388
rect 27396 30348 31852 30376
rect 27396 30336 27402 30348
rect 31846 30336 31852 30348
rect 31904 30376 31910 30388
rect 32398 30376 32404 30388
rect 31904 30348 32404 30376
rect 31904 30336 31910 30348
rect 32398 30336 32404 30348
rect 32456 30336 32462 30388
rect 35618 30336 35624 30388
rect 35676 30376 35682 30388
rect 38194 30376 38200 30388
rect 35676 30348 38200 30376
rect 35676 30336 35682 30348
rect 19168 30280 19288 30308
rect 13832 30212 15148 30240
rect 13832 30184 13860 30212
rect 16114 30200 16120 30252
rect 16172 30200 16178 30252
rect 16301 30243 16359 30249
rect 16301 30209 16313 30243
rect 16347 30240 16359 30243
rect 16758 30240 16764 30252
rect 16347 30212 16764 30240
rect 16347 30209 16359 30212
rect 16301 30203 16359 30209
rect 16758 30200 16764 30212
rect 16816 30200 16822 30252
rect 19168 30238 19196 30280
rect 19334 30268 19340 30320
rect 19392 30268 19398 30320
rect 19429 30311 19487 30317
rect 19429 30277 19441 30311
rect 19475 30308 19487 30311
rect 20165 30311 20223 30317
rect 20165 30308 20177 30311
rect 19475 30280 20177 30308
rect 19475 30277 19487 30280
rect 19429 30271 19487 30277
rect 20165 30277 20177 30280
rect 20211 30277 20223 30311
rect 20165 30271 20223 30277
rect 21082 30268 21088 30320
rect 21140 30268 21146 30320
rect 22462 30308 22468 30320
rect 21284 30280 22468 30308
rect 19240 30243 19298 30249
rect 19240 30238 19252 30243
rect 19168 30210 19252 30238
rect 19240 30209 19252 30210
rect 19286 30209 19298 30243
rect 19240 30203 19298 30209
rect 12161 30175 12219 30181
rect 12161 30141 12173 30175
rect 12207 30172 12219 30175
rect 12713 30175 12771 30181
rect 12713 30172 12725 30175
rect 12207 30144 12725 30172
rect 12207 30141 12219 30144
rect 12161 30135 12219 30141
rect 12713 30141 12725 30144
rect 12759 30141 12771 30175
rect 12713 30135 12771 30141
rect 13814 30132 13820 30184
rect 13872 30132 13878 30184
rect 14090 30132 14096 30184
rect 14148 30132 14154 30184
rect 15473 30175 15531 30181
rect 15473 30141 15485 30175
rect 15519 30172 15531 30175
rect 18414 30172 18420 30184
rect 15519 30144 18420 30172
rect 15519 30141 15531 30144
rect 15473 30135 15531 30141
rect 18414 30132 18420 30144
rect 18472 30132 18478 30184
rect 18509 30175 18567 30181
rect 18509 30141 18521 30175
rect 18555 30172 18567 30175
rect 19352 30172 19380 30268
rect 19518 30200 19524 30252
rect 19576 30249 19582 30252
rect 19576 30243 19615 30249
rect 19603 30209 19615 30243
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19576 30203 19615 30209
rect 19704 30209 19717 30240
rect 19751 30209 19763 30243
rect 19704 30203 19763 30209
rect 19576 30200 19582 30203
rect 18555 30144 19380 30172
rect 18555 30141 18567 30144
rect 18509 30135 18567 30141
rect 13078 30064 13084 30116
rect 13136 30064 13142 30116
rect 16298 30064 16304 30116
rect 16356 30064 16362 30116
rect 17494 30064 17500 30116
rect 17552 30104 17558 30116
rect 19242 30104 19248 30116
rect 17552 30076 19248 30104
rect 17552 30064 17558 30076
rect 19242 30064 19248 30076
rect 19300 30104 19306 30116
rect 19704 30104 19732 30203
rect 19978 30200 19984 30252
rect 20036 30240 20042 30252
rect 20349 30243 20407 30249
rect 20349 30240 20361 30243
rect 20036 30212 20361 30240
rect 20036 30200 20042 30212
rect 20349 30209 20361 30212
rect 20395 30209 20407 30243
rect 20349 30203 20407 30209
rect 20438 30200 20444 30252
rect 20496 30200 20502 30252
rect 21284 30249 21312 30280
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30209 21327 30243
rect 21269 30203 21327 30209
rect 22002 30200 22008 30252
rect 22060 30200 22066 30252
rect 22204 30249 22232 30280
rect 22462 30268 22468 30280
rect 22520 30308 22526 30320
rect 23017 30311 23075 30317
rect 23017 30308 23029 30311
rect 22520 30280 23029 30308
rect 22520 30268 22526 30280
rect 23017 30277 23029 30280
rect 23063 30308 23075 30311
rect 24949 30311 25007 30317
rect 24949 30308 24961 30311
rect 23063 30280 24961 30308
rect 23063 30277 23075 30280
rect 23017 30271 23075 30277
rect 24949 30277 24961 30280
rect 24995 30277 25007 30311
rect 25774 30308 25780 30320
rect 24949 30271 25007 30277
rect 25056 30280 25780 30308
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 22833 30243 22891 30249
rect 22833 30209 22845 30243
rect 22879 30209 22891 30243
rect 22833 30203 22891 30209
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30240 23995 30243
rect 25056 30240 25084 30280
rect 25774 30268 25780 30280
rect 25832 30308 25838 30320
rect 26694 30308 26700 30320
rect 25832 30280 26700 30308
rect 25832 30268 25838 30280
rect 26694 30268 26700 30280
rect 26752 30268 26758 30320
rect 27798 30308 27804 30320
rect 27356 30280 27804 30308
rect 23983 30212 25084 30240
rect 25133 30243 25191 30249
rect 23983 30209 23995 30212
rect 23937 30203 23995 30209
rect 25133 30209 25145 30243
rect 25179 30209 25191 30243
rect 25133 30203 25191 30209
rect 20165 30175 20223 30181
rect 20165 30141 20177 30175
rect 20211 30172 20223 30175
rect 20254 30172 20260 30184
rect 20211 30144 20260 30172
rect 20211 30141 20223 30144
rect 20165 30135 20223 30141
rect 20254 30132 20260 30144
rect 20312 30172 20318 30184
rect 21174 30172 21180 30184
rect 20312 30144 21180 30172
rect 20312 30132 20318 30144
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 21453 30175 21511 30181
rect 21453 30141 21465 30175
rect 21499 30172 21511 30175
rect 22848 30172 22876 30203
rect 23382 30172 23388 30184
rect 21499 30144 23388 30172
rect 21499 30141 21511 30144
rect 21453 30135 21511 30141
rect 23382 30132 23388 30144
rect 23440 30132 23446 30184
rect 19300 30076 19732 30104
rect 19300 30064 19306 30076
rect 21266 30064 21272 30116
rect 21324 30104 21330 30116
rect 21324 30076 22692 30104
rect 21324 30064 21330 30076
rect 22664 30048 22692 30076
rect 25038 30064 25044 30116
rect 25096 30104 25102 30116
rect 25148 30104 25176 30203
rect 25314 30200 25320 30252
rect 25372 30200 25378 30252
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30240 25467 30243
rect 25590 30240 25596 30252
rect 25455 30212 25596 30240
rect 25455 30209 25467 30212
rect 25409 30203 25467 30209
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 25866 30200 25872 30252
rect 25924 30200 25930 30252
rect 27356 30184 27384 30280
rect 27798 30268 27804 30280
rect 27856 30268 27862 30320
rect 28721 30311 28779 30317
rect 28721 30277 28733 30311
rect 28767 30308 28779 30311
rect 29086 30308 29092 30320
rect 28767 30280 29092 30308
rect 28767 30277 28779 30280
rect 28721 30271 28779 30277
rect 29086 30268 29092 30280
rect 29144 30268 29150 30320
rect 29362 30268 29368 30320
rect 29420 30308 29426 30320
rect 29914 30308 29920 30320
rect 29420 30280 29920 30308
rect 29420 30268 29426 30280
rect 29914 30268 29920 30280
rect 29972 30268 29978 30320
rect 30285 30311 30343 30317
rect 30285 30277 30297 30311
rect 30331 30308 30343 30311
rect 30742 30308 30748 30320
rect 30331 30280 30748 30308
rect 30331 30277 30343 30280
rect 30285 30271 30343 30277
rect 30742 30268 30748 30280
rect 30800 30268 30806 30320
rect 31202 30268 31208 30320
rect 31260 30268 31266 30320
rect 32030 30268 32036 30320
rect 32088 30308 32094 30320
rect 32585 30311 32643 30317
rect 32585 30308 32597 30311
rect 32088 30280 32597 30308
rect 32088 30268 32094 30280
rect 32585 30277 32597 30280
rect 32631 30277 32643 30311
rect 36817 30311 36875 30317
rect 36817 30308 36829 30311
rect 32585 30271 32643 30277
rect 32784 30280 36829 30308
rect 27433 30243 27491 30249
rect 27433 30209 27445 30243
rect 27479 30240 27491 30243
rect 27614 30240 27620 30252
rect 27479 30212 27620 30240
rect 27479 30209 27491 30212
rect 27433 30203 27491 30209
rect 27614 30200 27620 30212
rect 27672 30240 27678 30252
rect 28442 30240 28448 30252
rect 27672 30212 28448 30240
rect 27672 30200 27678 30212
rect 28442 30200 28448 30212
rect 28500 30200 28506 30252
rect 28629 30243 28687 30249
rect 28629 30209 28641 30243
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 27338 30132 27344 30184
rect 27396 30132 27402 30184
rect 28644 30172 28672 30203
rect 28810 30200 28816 30252
rect 28868 30200 28874 30252
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30240 29607 30243
rect 30006 30240 30012 30252
rect 29595 30212 30012 30240
rect 29595 30209 29607 30212
rect 29549 30203 29607 30209
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 30650 30200 30656 30252
rect 30708 30240 30714 30252
rect 31220 30240 31248 30268
rect 30708 30212 31248 30240
rect 31389 30243 31447 30249
rect 30708 30200 30714 30212
rect 31389 30209 31401 30243
rect 31435 30209 31447 30243
rect 31389 30203 31447 30209
rect 31665 30243 31723 30249
rect 31665 30209 31677 30243
rect 31711 30240 31723 30243
rect 32784 30240 32812 30280
rect 36817 30277 36829 30280
rect 36863 30308 36875 30311
rect 36998 30308 37004 30320
rect 36863 30280 37004 30308
rect 36863 30277 36875 30280
rect 36817 30271 36875 30277
rect 36998 30268 37004 30280
rect 37056 30268 37062 30320
rect 31711 30212 32812 30240
rect 32861 30243 32919 30249
rect 31711 30209 31723 30212
rect 31665 30203 31723 30209
rect 32861 30209 32873 30243
rect 32907 30240 32919 30243
rect 32950 30240 32956 30252
rect 32907 30212 32956 30240
rect 32907 30209 32919 30212
rect 32861 30203 32919 30209
rect 29638 30172 29644 30184
rect 28644 30144 29644 30172
rect 29638 30132 29644 30144
rect 29696 30132 29702 30184
rect 31021 30175 31079 30181
rect 31021 30141 31033 30175
rect 31067 30141 31079 30175
rect 31021 30135 31079 30141
rect 31036 30104 31064 30135
rect 31202 30132 31208 30184
rect 31260 30132 31266 30184
rect 31404 30172 31432 30203
rect 32950 30200 32956 30212
rect 33008 30200 33014 30252
rect 33962 30200 33968 30252
rect 34020 30240 34026 30252
rect 34057 30243 34115 30249
rect 34057 30240 34069 30243
rect 34020 30212 34069 30240
rect 34020 30200 34026 30212
rect 34057 30209 34069 30212
rect 34103 30240 34115 30243
rect 34146 30240 34152 30252
rect 34103 30212 34152 30240
rect 34103 30209 34115 30212
rect 34057 30203 34115 30209
rect 34146 30200 34152 30212
rect 34204 30200 34210 30252
rect 34514 30200 34520 30252
rect 34572 30200 34578 30252
rect 35342 30200 35348 30252
rect 35400 30240 35406 30252
rect 35437 30243 35495 30249
rect 35437 30240 35449 30243
rect 35400 30212 35449 30240
rect 35400 30200 35406 30212
rect 35437 30209 35449 30212
rect 35483 30209 35495 30243
rect 35437 30203 35495 30209
rect 31938 30172 31944 30184
rect 31404 30144 31944 30172
rect 31938 30132 31944 30144
rect 31996 30132 32002 30184
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30141 32643 30175
rect 32585 30135 32643 30141
rect 32769 30175 32827 30181
rect 32769 30141 32781 30175
rect 32815 30172 32827 30175
rect 33686 30172 33692 30184
rect 32815 30144 33692 30172
rect 32815 30141 32827 30144
rect 32769 30135 32827 30141
rect 25096 30076 31064 30104
rect 25096 30064 25102 30076
rect 13173 30039 13231 30045
rect 13173 30005 13185 30039
rect 13219 30036 13231 30039
rect 13538 30036 13544 30048
rect 13219 30008 13544 30036
rect 13219 30005 13231 30008
rect 13173 29999 13231 30005
rect 13538 29996 13544 30008
rect 13596 29996 13602 30048
rect 17862 29996 17868 30048
rect 17920 29996 17926 30048
rect 18138 29996 18144 30048
rect 18196 30036 18202 30048
rect 19061 30039 19119 30045
rect 19061 30036 19073 30039
rect 18196 30008 19073 30036
rect 18196 29996 18202 30008
rect 19061 30005 19073 30008
rect 19107 30005 19119 30039
rect 19061 29999 19119 30005
rect 20162 29996 20168 30048
rect 20220 30036 20226 30048
rect 20438 30036 20444 30048
rect 20220 30008 20444 30036
rect 20220 29996 20226 30008
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 21174 29996 21180 30048
rect 21232 30036 21238 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21232 30008 22017 30036
rect 21232 29996 21238 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22005 29999 22063 30005
rect 22646 29996 22652 30048
rect 22704 29996 22710 30048
rect 24302 29996 24308 30048
rect 24360 30036 24366 30048
rect 24397 30039 24455 30045
rect 24397 30036 24409 30039
rect 24360 30008 24409 30036
rect 24360 29996 24366 30008
rect 24397 30005 24409 30008
rect 24443 30036 24455 30039
rect 24670 30036 24676 30048
rect 24443 30008 24676 30036
rect 24443 30005 24455 30008
rect 24397 29999 24455 30005
rect 24670 29996 24676 30008
rect 24728 29996 24734 30048
rect 26142 29996 26148 30048
rect 26200 30036 26206 30048
rect 26513 30039 26571 30045
rect 26513 30036 26525 30039
rect 26200 30008 26525 30036
rect 26200 29996 26206 30008
rect 26513 30005 26525 30008
rect 26559 30036 26571 30039
rect 26786 30036 26792 30048
rect 26559 30008 26792 30036
rect 26559 30005 26571 30008
rect 26513 29999 26571 30005
rect 26786 29996 26792 30008
rect 26844 29996 26850 30048
rect 27706 29996 27712 30048
rect 27764 29996 27770 30048
rect 29733 30039 29791 30045
rect 29733 30005 29745 30039
rect 29779 30036 29791 30039
rect 29822 30036 29828 30048
rect 29779 30008 29828 30036
rect 29779 30005 29791 30008
rect 29733 29999 29791 30005
rect 29822 29996 29828 30008
rect 29880 29996 29886 30048
rect 32600 30036 32628 30135
rect 33686 30132 33692 30144
rect 33744 30132 33750 30184
rect 33873 30175 33931 30181
rect 33873 30141 33885 30175
rect 33919 30172 33931 30175
rect 35452 30172 35480 30203
rect 35710 30200 35716 30252
rect 35768 30200 35774 30252
rect 35802 30200 35808 30252
rect 35860 30200 35866 30252
rect 36725 30243 36783 30249
rect 36725 30209 36737 30243
rect 36771 30209 36783 30243
rect 36725 30203 36783 30209
rect 36909 30243 36967 30249
rect 36909 30209 36921 30243
rect 36955 30209 36967 30243
rect 36909 30203 36967 30209
rect 36446 30172 36452 30184
rect 33919 30144 34008 30172
rect 35452 30144 36452 30172
rect 33919 30141 33931 30144
rect 33873 30135 33931 30141
rect 33980 30116 34008 30144
rect 36446 30132 36452 30144
rect 36504 30172 36510 30184
rect 36740 30172 36768 30203
rect 36504 30144 36768 30172
rect 36504 30132 36510 30144
rect 33962 30064 33968 30116
rect 34020 30064 34026 30116
rect 36924 30104 36952 30203
rect 37274 30200 37280 30252
rect 37332 30240 37338 30252
rect 37568 30249 37596 30348
rect 38194 30336 38200 30348
rect 38252 30336 38258 30388
rect 40034 30336 40040 30388
rect 40092 30376 40098 30388
rect 40862 30376 40868 30388
rect 40092 30348 40868 30376
rect 40092 30336 40098 30348
rect 40862 30336 40868 30348
rect 40920 30376 40926 30388
rect 41138 30376 41144 30388
rect 40920 30348 41144 30376
rect 40920 30336 40926 30348
rect 41138 30336 41144 30348
rect 41196 30336 41202 30388
rect 41322 30336 41328 30388
rect 41380 30376 41386 30388
rect 41690 30376 41696 30388
rect 41380 30348 41696 30376
rect 41380 30336 41386 30348
rect 41690 30336 41696 30348
rect 41748 30336 41754 30388
rect 37918 30268 37924 30320
rect 37976 30308 37982 30320
rect 38013 30311 38071 30317
rect 38013 30308 38025 30311
rect 37976 30280 38025 30308
rect 37976 30268 37982 30280
rect 38013 30277 38025 30280
rect 38059 30277 38071 30311
rect 38013 30271 38071 30277
rect 38102 30268 38108 30320
rect 38160 30308 38166 30320
rect 39853 30311 39911 30317
rect 39853 30308 39865 30311
rect 38160 30280 39865 30308
rect 38160 30268 38166 30280
rect 39853 30277 39865 30280
rect 39899 30277 39911 30311
rect 39853 30271 39911 30277
rect 40586 30268 40592 30320
rect 40644 30308 40650 30320
rect 40773 30311 40831 30317
rect 40773 30308 40785 30311
rect 40644 30280 40785 30308
rect 40644 30268 40650 30280
rect 40773 30277 40785 30280
rect 40819 30277 40831 30311
rect 40773 30271 40831 30277
rect 40957 30311 41015 30317
rect 40957 30277 40969 30311
rect 41003 30308 41015 30311
rect 41414 30308 41420 30320
rect 41003 30280 41420 30308
rect 41003 30277 41015 30280
rect 40957 30271 41015 30277
rect 41414 30268 41420 30280
rect 41472 30268 41478 30320
rect 37461 30243 37519 30249
rect 37461 30240 37473 30243
rect 37332 30212 37473 30240
rect 37332 30200 37338 30212
rect 37461 30209 37473 30212
rect 37507 30209 37519 30243
rect 37461 30203 37519 30209
rect 37553 30243 37611 30249
rect 37553 30209 37565 30243
rect 37599 30209 37611 30243
rect 37553 30203 37611 30209
rect 37734 30200 37740 30252
rect 37792 30200 37798 30252
rect 37826 30200 37832 30252
rect 37884 30249 37890 30252
rect 37884 30240 37896 30249
rect 37884 30212 37929 30240
rect 37884 30203 37896 30212
rect 37884 30200 37890 30203
rect 38194 30200 38200 30252
rect 38252 30240 38258 30252
rect 38933 30243 38991 30249
rect 38933 30240 38945 30243
rect 38252 30212 38945 30240
rect 38252 30200 38258 30212
rect 38933 30209 38945 30212
rect 38979 30240 38991 30243
rect 38979 30212 39160 30240
rect 38979 30209 38991 30212
rect 38933 30203 38991 30209
rect 38746 30132 38752 30184
rect 38804 30172 38810 30184
rect 39025 30175 39083 30181
rect 39025 30172 39037 30175
rect 38804 30144 39037 30172
rect 38804 30132 38810 30144
rect 39025 30141 39037 30144
rect 39071 30141 39083 30175
rect 39132 30172 39160 30212
rect 39574 30200 39580 30252
rect 39632 30240 39638 30252
rect 39761 30243 39819 30249
rect 39761 30240 39773 30243
rect 39632 30212 39773 30240
rect 39632 30200 39638 30212
rect 39761 30209 39773 30212
rect 39807 30209 39819 30243
rect 39761 30203 39819 30209
rect 39945 30243 40003 30249
rect 39945 30209 39957 30243
rect 39991 30240 40003 30243
rect 40126 30240 40132 30252
rect 39991 30212 40132 30240
rect 39991 30209 40003 30212
rect 39945 30203 40003 30209
rect 40126 30200 40132 30212
rect 40184 30200 40190 30252
rect 41141 30243 41199 30249
rect 41141 30209 41153 30243
rect 41187 30209 41199 30243
rect 41141 30203 41199 30209
rect 42061 30243 42119 30249
rect 42061 30209 42073 30243
rect 42107 30240 42119 30243
rect 43073 30243 43131 30249
rect 42107 30212 42656 30240
rect 42107 30209 42119 30212
rect 42061 30203 42119 30209
rect 41156 30172 41184 30203
rect 42628 30181 42656 30212
rect 43073 30209 43085 30243
rect 43119 30240 43131 30243
rect 43254 30240 43260 30252
rect 43119 30212 43260 30240
rect 43119 30209 43131 30212
rect 43073 30203 43131 30209
rect 43254 30200 43260 30212
rect 43312 30200 43318 30252
rect 42613 30175 42671 30181
rect 39132 30144 42104 30172
rect 39025 30135 39083 30141
rect 42076 30116 42104 30144
rect 42613 30141 42625 30175
rect 42659 30141 42671 30175
rect 42613 30135 42671 30141
rect 39574 30104 39580 30116
rect 36924 30076 39580 30104
rect 39574 30064 39580 30076
rect 39632 30064 39638 30116
rect 40494 30064 40500 30116
rect 40552 30104 40558 30116
rect 41877 30107 41935 30113
rect 41877 30104 41889 30107
rect 40552 30076 41889 30104
rect 40552 30064 40558 30076
rect 41877 30073 41889 30076
rect 41923 30073 41935 30107
rect 41877 30067 41935 30073
rect 42058 30064 42064 30116
rect 42116 30064 42122 30116
rect 32766 30036 32772 30048
rect 32600 30008 32772 30036
rect 32766 29996 32772 30008
rect 32824 30036 32830 30048
rect 38378 30036 38384 30048
rect 32824 30008 38384 30036
rect 32824 29996 32830 30008
rect 38378 29996 38384 30008
rect 38436 29996 38442 30048
rect 39022 29996 39028 30048
rect 39080 29996 39086 30048
rect 39301 30039 39359 30045
rect 39301 30005 39313 30039
rect 39347 30036 39359 30039
rect 39666 30036 39672 30048
rect 39347 30008 39672 30036
rect 39347 30005 39359 30008
rect 39301 29999 39359 30005
rect 39666 29996 39672 30008
rect 39724 29996 39730 30048
rect 42794 29996 42800 30048
rect 42852 29996 42858 30048
rect 1104 29946 43884 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 43884 29946
rect 1104 29872 43884 29894
rect 11974 29792 11980 29844
rect 12032 29792 12038 29844
rect 12621 29835 12679 29841
rect 12621 29801 12633 29835
rect 12667 29832 12679 29835
rect 12986 29832 12992 29844
rect 12667 29804 12992 29832
rect 12667 29801 12679 29804
rect 12621 29795 12679 29801
rect 12986 29792 12992 29804
rect 13044 29792 13050 29844
rect 13725 29835 13783 29841
rect 13725 29801 13737 29835
rect 13771 29832 13783 29835
rect 14090 29832 14096 29844
rect 13771 29804 14096 29832
rect 13771 29801 13783 29804
rect 13725 29795 13783 29801
rect 14090 29792 14096 29804
rect 14148 29792 14154 29844
rect 18598 29832 18604 29844
rect 16684 29804 18604 29832
rect 13630 29764 13636 29776
rect 12176 29736 13636 29764
rect 12176 29705 12204 29736
rect 13630 29724 13636 29736
rect 13688 29724 13694 29776
rect 12161 29699 12219 29705
rect 12161 29665 12173 29699
rect 12207 29665 12219 29699
rect 12161 29659 12219 29665
rect 15473 29699 15531 29705
rect 15473 29665 15485 29699
rect 15519 29696 15531 29699
rect 16114 29696 16120 29708
rect 15519 29668 16120 29696
rect 15519 29665 15531 29668
rect 15473 29659 15531 29665
rect 16114 29656 16120 29668
rect 16172 29696 16178 29708
rect 16684 29705 16712 29804
rect 18598 29792 18604 29804
rect 18656 29792 18662 29844
rect 18690 29792 18696 29844
rect 18748 29832 18754 29844
rect 20346 29832 20352 29844
rect 18748 29804 20352 29832
rect 18748 29792 18754 29804
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 20990 29792 20996 29844
rect 21048 29832 21054 29844
rect 21048 29804 21864 29832
rect 21048 29792 21054 29804
rect 16850 29724 16856 29776
rect 16908 29764 16914 29776
rect 18877 29767 18935 29773
rect 18877 29764 18889 29767
rect 16908 29736 18889 29764
rect 16908 29724 16914 29736
rect 18877 29733 18889 29736
rect 18923 29733 18935 29767
rect 18877 29727 18935 29733
rect 21453 29767 21511 29773
rect 21453 29733 21465 29767
rect 21499 29733 21511 29767
rect 21836 29764 21864 29804
rect 21910 29792 21916 29844
rect 21968 29792 21974 29844
rect 22370 29792 22376 29844
rect 22428 29792 22434 29844
rect 25685 29835 25743 29841
rect 25685 29801 25697 29835
rect 25731 29832 25743 29835
rect 26050 29832 26056 29844
rect 25731 29804 26056 29832
rect 25731 29801 25743 29804
rect 25685 29795 25743 29801
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 27525 29835 27583 29841
rect 27525 29801 27537 29835
rect 27571 29832 27583 29835
rect 27614 29832 27620 29844
rect 27571 29804 27620 29832
rect 27571 29801 27583 29804
rect 27525 29795 27583 29801
rect 27614 29792 27620 29804
rect 27672 29792 27678 29844
rect 27706 29792 27712 29844
rect 27764 29832 27770 29844
rect 35986 29832 35992 29844
rect 27764 29804 35992 29832
rect 27764 29792 27770 29804
rect 35986 29792 35992 29804
rect 36044 29792 36050 29844
rect 36081 29835 36139 29841
rect 36081 29801 36093 29835
rect 36127 29832 36139 29835
rect 36906 29832 36912 29844
rect 36127 29804 36912 29832
rect 36127 29801 36139 29804
rect 36081 29795 36139 29801
rect 36906 29792 36912 29804
rect 36964 29792 36970 29844
rect 36998 29792 37004 29844
rect 37056 29792 37062 29844
rect 39206 29792 39212 29844
rect 39264 29792 39270 29844
rect 39574 29792 39580 29844
rect 39632 29832 39638 29844
rect 41233 29835 41291 29841
rect 41233 29832 41245 29835
rect 39632 29804 41245 29832
rect 39632 29792 39638 29804
rect 41233 29801 41245 29804
rect 41279 29801 41291 29835
rect 41233 29795 41291 29801
rect 41322 29792 41328 29844
rect 41380 29832 41386 29844
rect 41417 29835 41475 29841
rect 41417 29832 41429 29835
rect 41380 29804 41429 29832
rect 41380 29792 41386 29804
rect 41417 29801 41429 29804
rect 41463 29801 41475 29835
rect 41417 29795 41475 29801
rect 24026 29764 24032 29776
rect 21836 29736 24032 29764
rect 21453 29727 21511 29733
rect 16485 29699 16543 29705
rect 16485 29696 16497 29699
rect 16172 29668 16497 29696
rect 16172 29656 16178 29668
rect 16485 29665 16497 29668
rect 16531 29665 16543 29699
rect 16485 29659 16543 29665
rect 16669 29699 16727 29705
rect 16669 29665 16681 29699
rect 16715 29665 16727 29699
rect 19705 29699 19763 29705
rect 19705 29696 19717 29699
rect 16669 29659 16727 29665
rect 17328 29668 19717 29696
rect 11425 29631 11483 29637
rect 11425 29597 11437 29631
rect 11471 29628 11483 29631
rect 11882 29628 11888 29640
rect 11471 29600 11888 29628
rect 11471 29597 11483 29600
rect 11425 29591 11483 29597
rect 11882 29588 11888 29600
rect 11940 29588 11946 29640
rect 12802 29588 12808 29640
rect 12860 29588 12866 29640
rect 12986 29588 12992 29640
rect 13044 29588 13050 29640
rect 13081 29631 13139 29637
rect 13081 29597 13093 29631
rect 13127 29628 13139 29631
rect 13170 29628 13176 29640
rect 13127 29600 13176 29628
rect 13127 29597 13139 29600
rect 13081 29591 13139 29597
rect 13170 29588 13176 29600
rect 13228 29588 13234 29640
rect 13538 29588 13544 29640
rect 13596 29588 13602 29640
rect 14274 29588 14280 29640
rect 14332 29588 14338 29640
rect 14461 29631 14519 29637
rect 14461 29597 14473 29631
rect 14507 29597 14519 29631
rect 14461 29591 14519 29597
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29628 15439 29631
rect 15930 29628 15936 29640
rect 15427 29600 15936 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 12161 29563 12219 29569
rect 12161 29529 12173 29563
rect 12207 29560 12219 29563
rect 14476 29560 14504 29591
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16298 29588 16304 29640
rect 16356 29628 16362 29640
rect 17221 29631 17279 29637
rect 17221 29628 17233 29631
rect 16356 29600 17233 29628
rect 16356 29588 16362 29600
rect 17221 29597 17233 29600
rect 17267 29597 17279 29631
rect 17221 29591 17279 29597
rect 12207 29532 14504 29560
rect 12207 29529 12219 29532
rect 12161 29523 12219 29529
rect 16114 29520 16120 29572
rect 16172 29560 16178 29572
rect 17328 29560 17356 29668
rect 19705 29665 19717 29668
rect 19751 29665 19763 29699
rect 19705 29659 19763 29665
rect 17405 29631 17463 29637
rect 17405 29597 17417 29631
rect 17451 29628 17463 29631
rect 17494 29628 17500 29640
rect 17451 29600 17500 29628
rect 17451 29597 17463 29600
rect 17405 29591 17463 29597
rect 17494 29588 17500 29600
rect 17552 29588 17558 29640
rect 17862 29588 17868 29640
rect 17920 29588 17926 29640
rect 18138 29588 18144 29640
rect 18196 29588 18202 29640
rect 18690 29588 18696 29640
rect 18748 29588 18754 29640
rect 18874 29588 18880 29640
rect 18932 29588 18938 29640
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19981 29631 20039 29637
rect 19981 29628 19993 29631
rect 19024 29600 19993 29628
rect 19024 29588 19030 29600
rect 19981 29597 19993 29600
rect 20027 29597 20039 29631
rect 19981 29591 20039 29597
rect 20070 29588 20076 29640
rect 20128 29588 20134 29640
rect 20162 29588 20168 29640
rect 20220 29588 20226 29640
rect 20346 29588 20352 29640
rect 20404 29588 20410 29640
rect 21174 29588 21180 29640
rect 21232 29588 21238 29640
rect 21468 29628 21496 29727
rect 24026 29724 24032 29736
rect 24084 29724 24090 29776
rect 27798 29724 27804 29776
rect 27856 29764 27862 29776
rect 27985 29767 28043 29773
rect 27985 29764 27997 29767
rect 27856 29736 27997 29764
rect 27856 29724 27862 29736
rect 27985 29733 27997 29736
rect 28031 29733 28043 29767
rect 27985 29727 28043 29733
rect 31018 29724 31024 29776
rect 31076 29764 31082 29776
rect 31113 29767 31171 29773
rect 31113 29764 31125 29767
rect 31076 29736 31125 29764
rect 31076 29724 31082 29736
rect 31113 29733 31125 29736
rect 31159 29733 31171 29767
rect 31113 29727 31171 29733
rect 33226 29724 33232 29776
rect 33284 29764 33290 29776
rect 34054 29764 34060 29776
rect 33284 29736 34060 29764
rect 33284 29724 33290 29736
rect 34054 29724 34060 29736
rect 34112 29764 34118 29776
rect 35069 29767 35127 29773
rect 35069 29764 35081 29767
rect 34112 29736 35081 29764
rect 34112 29724 34118 29736
rect 35069 29733 35081 29736
rect 35115 29764 35127 29767
rect 35342 29764 35348 29776
rect 35115 29736 35348 29764
rect 35115 29733 35127 29736
rect 35069 29727 35127 29733
rect 35342 29724 35348 29736
rect 35400 29724 35406 29776
rect 36449 29767 36507 29773
rect 36449 29733 36461 29767
rect 36495 29764 36507 29767
rect 37826 29764 37832 29776
rect 36495 29736 37832 29764
rect 36495 29733 36507 29736
rect 36449 29727 36507 29733
rect 37826 29724 37832 29736
rect 37884 29764 37890 29776
rect 38013 29767 38071 29773
rect 38013 29764 38025 29767
rect 37884 29736 38025 29764
rect 37884 29724 37890 29736
rect 38013 29733 38025 29736
rect 38059 29733 38071 29767
rect 38013 29727 38071 29733
rect 38562 29724 38568 29776
rect 38620 29764 38626 29776
rect 38620 29736 40540 29764
rect 38620 29724 38626 29736
rect 23290 29656 23296 29708
rect 23348 29696 23354 29708
rect 23937 29699 23995 29705
rect 23937 29696 23949 29699
rect 23348 29668 23949 29696
rect 23348 29656 23354 29668
rect 23937 29665 23949 29668
rect 23983 29665 23995 29699
rect 23937 29659 23995 29665
rect 22097 29631 22155 29637
rect 22097 29628 22109 29631
rect 21468 29600 22109 29628
rect 22097 29597 22109 29600
rect 22143 29597 22155 29631
rect 22097 29591 22155 29597
rect 22186 29588 22192 29640
rect 22244 29588 22250 29640
rect 22465 29631 22523 29637
rect 22465 29597 22477 29631
rect 22511 29628 22523 29631
rect 22554 29628 22560 29640
rect 22511 29600 22560 29628
rect 22511 29597 22523 29600
rect 22465 29591 22523 29597
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22704 29600 23121 29628
rect 22704 29588 22710 29600
rect 23109 29597 23121 29600
rect 23155 29597 23167 29631
rect 23109 29591 23167 29597
rect 23385 29631 23443 29637
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 19334 29560 19340 29572
rect 16172 29532 17356 29560
rect 18064 29532 19340 29560
rect 16172 29520 16178 29532
rect 12986 29452 12992 29504
rect 13044 29492 13050 29504
rect 14277 29495 14335 29501
rect 14277 29492 14289 29495
rect 13044 29464 14289 29492
rect 13044 29452 13050 29464
rect 14277 29461 14289 29464
rect 14323 29461 14335 29495
rect 14277 29455 14335 29461
rect 15838 29452 15844 29504
rect 15896 29492 15902 29504
rect 16025 29495 16083 29501
rect 16025 29492 16037 29495
rect 15896 29464 16037 29492
rect 15896 29452 15902 29464
rect 16025 29461 16037 29464
rect 16071 29461 16083 29495
rect 16025 29455 16083 29461
rect 16390 29452 16396 29504
rect 16448 29452 16454 29504
rect 17310 29452 17316 29504
rect 17368 29452 17374 29504
rect 17954 29452 17960 29504
rect 18012 29501 18018 29504
rect 18064 29501 18092 29532
rect 19334 29520 19340 29532
rect 19392 29520 19398 29572
rect 20990 29520 20996 29572
rect 21048 29560 21054 29572
rect 21269 29563 21327 29569
rect 21269 29560 21281 29563
rect 21048 29532 21281 29560
rect 21048 29520 21054 29532
rect 21269 29529 21281 29532
rect 21315 29529 21327 29563
rect 21269 29523 21327 29529
rect 21453 29563 21511 29569
rect 21453 29529 21465 29563
rect 21499 29560 21511 29563
rect 22925 29563 22983 29569
rect 22925 29560 22937 29563
rect 21499 29532 22937 29560
rect 21499 29529 21511 29532
rect 21453 29523 21511 29529
rect 22925 29529 22937 29532
rect 22971 29529 22983 29563
rect 23400 29560 23428 29591
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 24044 29637 24072 29724
rect 24946 29656 24952 29708
rect 25004 29696 25010 29708
rect 36998 29696 37004 29708
rect 25004 29668 25176 29696
rect 25004 29656 25010 29668
rect 23845 29631 23903 29637
rect 23845 29628 23857 29631
rect 23532 29600 23857 29628
rect 23532 29588 23538 29600
rect 23845 29597 23857 29600
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29597 24087 29631
rect 24029 29591 24087 29597
rect 24578 29588 24584 29640
rect 24636 29628 24642 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24636 29600 24777 29628
rect 24636 29588 24642 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 24854 29588 24860 29640
rect 24912 29588 24918 29640
rect 25148 29637 25176 29668
rect 32692 29668 37004 29696
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29628 25191 29631
rect 25866 29628 25872 29640
rect 25179 29600 25872 29628
rect 25179 29597 25191 29600
rect 25133 29591 25191 29597
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 26145 29631 26203 29637
rect 26145 29597 26157 29631
rect 26191 29628 26203 29631
rect 26786 29628 26792 29640
rect 26191 29600 26792 29628
rect 26191 29597 26203 29600
rect 26145 29591 26203 29597
rect 26786 29588 26792 29600
rect 26844 29628 26850 29640
rect 29089 29631 29147 29637
rect 29089 29628 29101 29631
rect 26844 29600 29101 29628
rect 26844 29588 26850 29600
rect 29089 29597 29101 29600
rect 29135 29597 29147 29631
rect 29089 29591 29147 29597
rect 29730 29588 29736 29640
rect 29788 29588 29794 29640
rect 29822 29588 29828 29640
rect 29880 29628 29886 29640
rect 32692 29637 32720 29668
rect 29989 29631 30047 29637
rect 29989 29628 30001 29631
rect 29880 29600 30001 29628
rect 29880 29588 29886 29600
rect 29989 29597 30001 29600
rect 30035 29597 30047 29631
rect 29989 29591 30047 29597
rect 32677 29631 32735 29637
rect 32677 29597 32689 29631
rect 32723 29597 32735 29631
rect 32677 29591 32735 29597
rect 32861 29631 32919 29637
rect 32861 29597 32873 29631
rect 32907 29628 32919 29631
rect 33226 29628 33232 29640
rect 32907 29600 33232 29628
rect 32907 29597 32919 29600
rect 32861 29591 32919 29597
rect 33226 29588 33232 29600
rect 33284 29588 33290 29640
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29628 33379 29631
rect 33410 29628 33416 29640
rect 33367 29600 33416 29628
rect 33367 29597 33379 29600
rect 33321 29591 33379 29597
rect 33410 29588 33416 29600
rect 33468 29588 33474 29640
rect 33505 29631 33563 29637
rect 33505 29597 33517 29631
rect 33551 29628 33563 29631
rect 33870 29628 33876 29640
rect 33551 29600 33876 29628
rect 33551 29597 33563 29600
rect 33505 29591 33563 29597
rect 33870 29588 33876 29600
rect 33928 29588 33934 29640
rect 33980 29637 34008 29668
rect 36998 29656 37004 29668
rect 37056 29656 37062 29708
rect 37185 29699 37243 29705
rect 37185 29665 37197 29699
rect 37231 29696 37243 29699
rect 38102 29696 38108 29708
rect 37231 29668 38108 29696
rect 37231 29665 37243 29668
rect 37185 29659 37243 29665
rect 38102 29656 38108 29668
rect 38160 29656 38166 29708
rect 40236 29705 40264 29736
rect 38841 29699 38899 29705
rect 38841 29665 38853 29699
rect 38887 29696 38899 29699
rect 40037 29699 40095 29705
rect 40037 29696 40049 29699
rect 38887 29668 40049 29696
rect 38887 29665 38899 29668
rect 38841 29659 38899 29665
rect 40037 29665 40049 29668
rect 40083 29665 40095 29699
rect 40037 29659 40095 29665
rect 40221 29699 40279 29705
rect 40221 29665 40233 29699
rect 40267 29665 40279 29699
rect 40221 29659 40279 29665
rect 40310 29656 40316 29708
rect 40368 29656 40374 29708
rect 40402 29656 40408 29708
rect 40460 29656 40466 29708
rect 40512 29696 40540 29736
rect 40586 29724 40592 29776
rect 40644 29764 40650 29776
rect 42242 29764 42248 29776
rect 40644 29736 42248 29764
rect 40644 29724 40650 29736
rect 42242 29724 42248 29736
rect 42300 29724 42306 29776
rect 42886 29724 42892 29776
rect 42944 29724 42950 29776
rect 41138 29696 41144 29708
rect 40512 29668 41144 29696
rect 41138 29656 41144 29668
rect 41196 29656 41202 29708
rect 41414 29656 41420 29708
rect 41472 29696 41478 29708
rect 41472 29668 41644 29696
rect 41472 29656 41478 29668
rect 33965 29631 34023 29637
rect 33965 29597 33977 29631
rect 34011 29597 34023 29631
rect 33965 29591 34023 29597
rect 34054 29588 34060 29640
rect 34112 29628 34118 29640
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 34112 29600 34161 29628
rect 34112 29588 34118 29600
rect 34149 29597 34161 29600
rect 34195 29628 34207 29631
rect 34238 29628 34244 29640
rect 34195 29600 34244 29628
rect 34195 29597 34207 29600
rect 34149 29591 34207 29597
rect 34238 29588 34244 29600
rect 34296 29588 34302 29640
rect 34514 29588 34520 29640
rect 34572 29628 34578 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34572 29600 34897 29628
rect 34572 29588 34578 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 36170 29588 36176 29640
rect 36228 29628 36234 29640
rect 36265 29631 36323 29637
rect 36265 29628 36277 29631
rect 36228 29600 36277 29628
rect 36228 29588 36234 29600
rect 36265 29597 36277 29600
rect 36311 29597 36323 29631
rect 36265 29591 36323 29597
rect 36541 29631 36599 29637
rect 36541 29597 36553 29631
rect 36587 29628 36599 29631
rect 37090 29628 37096 29640
rect 36587 29600 37096 29628
rect 36587 29597 36599 29600
rect 36541 29591 36599 29597
rect 37090 29588 37096 29600
rect 37148 29588 37154 29640
rect 37274 29588 37280 29640
rect 37332 29588 37338 29640
rect 37918 29588 37924 29640
rect 37976 29628 37982 29640
rect 38013 29631 38071 29637
rect 38013 29628 38025 29631
rect 37976 29600 38025 29628
rect 37976 29588 37982 29600
rect 38013 29597 38025 29600
rect 38059 29597 38071 29631
rect 38013 29591 38071 29597
rect 38197 29631 38255 29637
rect 38197 29597 38209 29631
rect 38243 29628 38255 29631
rect 38562 29628 38568 29640
rect 38243 29600 38568 29628
rect 38243 29597 38255 29600
rect 38197 29591 38255 29597
rect 38562 29588 38568 29600
rect 38620 29588 38626 29640
rect 38933 29631 38991 29637
rect 38933 29597 38945 29631
rect 38979 29597 38991 29631
rect 38933 29591 38991 29597
rect 39301 29631 39359 29637
rect 39301 29597 39313 29631
rect 39347 29628 39359 29631
rect 39942 29628 39948 29640
rect 39347 29600 39948 29628
rect 39347 29597 39359 29600
rect 39301 29591 39359 29597
rect 24210 29560 24216 29572
rect 23400 29532 24216 29560
rect 22925 29523 22983 29529
rect 23492 29504 23520 29532
rect 24210 29520 24216 29532
rect 24268 29520 24274 29572
rect 24949 29563 25007 29569
rect 24949 29529 24961 29563
rect 24995 29560 25007 29563
rect 25222 29560 25228 29572
rect 24995 29532 25228 29560
rect 24995 29529 25007 29532
rect 24949 29523 25007 29529
rect 25222 29520 25228 29532
rect 25280 29520 25286 29572
rect 26412 29563 26470 29569
rect 26412 29529 26424 29563
rect 26458 29560 26470 29563
rect 28626 29560 28632 29572
rect 26458 29532 28632 29560
rect 26458 29529 26470 29532
rect 26412 29523 26470 29529
rect 28626 29520 28632 29532
rect 28684 29520 28690 29572
rect 31202 29520 31208 29572
rect 31260 29560 31266 29572
rect 31665 29563 31723 29569
rect 31665 29560 31677 29563
rect 31260 29532 31677 29560
rect 31260 29520 31266 29532
rect 31665 29529 31677 29532
rect 31711 29529 31723 29563
rect 32493 29563 32551 29569
rect 32493 29560 32505 29563
rect 31665 29523 31723 29529
rect 31864 29532 32505 29560
rect 18012 29455 18021 29501
rect 18049 29495 18107 29501
rect 18049 29461 18061 29495
rect 18095 29461 18107 29495
rect 18049 29455 18107 29461
rect 18012 29452 18018 29455
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 22002 29492 22008 29504
rect 19208 29464 22008 29492
rect 19208 29452 19214 29464
rect 22002 29452 22008 29464
rect 22060 29492 22066 29504
rect 23474 29492 23480 29504
rect 22060 29464 23480 29492
rect 22060 29452 22066 29464
rect 23474 29452 23480 29464
rect 23532 29452 23538 29504
rect 24578 29452 24584 29504
rect 24636 29452 24642 29504
rect 28534 29452 28540 29504
rect 28592 29452 28598 29504
rect 31110 29452 31116 29504
rect 31168 29492 31174 29504
rect 31864 29492 31892 29532
rect 32493 29529 32505 29532
rect 32539 29529 32551 29563
rect 32493 29523 32551 29529
rect 34422 29520 34428 29572
rect 34480 29560 34486 29572
rect 36722 29560 36728 29572
rect 34480 29532 36728 29560
rect 34480 29520 34486 29532
rect 36722 29520 36728 29532
rect 36780 29520 36786 29572
rect 36998 29520 37004 29572
rect 37056 29520 37062 29572
rect 38948 29560 38976 29591
rect 39942 29588 39948 29600
rect 40000 29588 40006 29640
rect 40497 29631 40555 29637
rect 40497 29628 40509 29631
rect 40052 29600 40509 29628
rect 37108 29532 38976 29560
rect 31168 29464 31892 29492
rect 31168 29452 31174 29464
rect 31938 29452 31944 29504
rect 31996 29452 32002 29504
rect 33413 29495 33471 29501
rect 33413 29461 33425 29495
rect 33459 29492 33471 29495
rect 34054 29492 34060 29504
rect 33459 29464 34060 29492
rect 33459 29461 33471 29464
rect 33413 29455 33471 29461
rect 34054 29452 34060 29464
rect 34112 29452 34118 29504
rect 34333 29495 34391 29501
rect 34333 29461 34345 29495
rect 34379 29492 34391 29495
rect 34514 29492 34520 29504
rect 34379 29464 34520 29492
rect 34379 29461 34391 29464
rect 34333 29455 34391 29461
rect 34514 29452 34520 29464
rect 34572 29452 34578 29504
rect 35158 29452 35164 29504
rect 35216 29492 35222 29504
rect 37108 29492 37136 29532
rect 39022 29520 39028 29572
rect 39080 29560 39086 29572
rect 40052 29560 40080 29600
rect 40497 29597 40509 29600
rect 40543 29597 40555 29631
rect 40497 29591 40555 29597
rect 41506 29588 41512 29640
rect 41564 29588 41570 29640
rect 41616 29637 41644 29668
rect 41601 29631 41659 29637
rect 41601 29597 41613 29631
rect 41647 29628 41659 29631
rect 41647 29600 42472 29628
rect 41647 29597 41659 29600
rect 41601 29591 41659 29597
rect 39080 29532 40080 29560
rect 39080 29520 39086 29532
rect 41322 29520 41328 29572
rect 41380 29560 41386 29572
rect 42242 29560 42248 29572
rect 41380 29532 42248 29560
rect 41380 29520 41386 29532
rect 42242 29520 42248 29532
rect 42300 29520 42306 29572
rect 42444 29569 42472 29600
rect 42429 29563 42487 29569
rect 42429 29529 42441 29563
rect 42475 29560 42487 29563
rect 42610 29560 42616 29572
rect 42475 29532 42616 29560
rect 42475 29529 42487 29532
rect 42429 29523 42487 29529
rect 42610 29520 42616 29532
rect 42668 29520 42674 29572
rect 42886 29520 42892 29572
rect 42944 29560 42950 29572
rect 43073 29563 43131 29569
rect 43073 29560 43085 29563
rect 42944 29532 43085 29560
rect 42944 29520 42950 29532
rect 43073 29529 43085 29532
rect 43119 29529 43131 29563
rect 43073 29523 43131 29529
rect 43254 29520 43260 29572
rect 43312 29520 43318 29572
rect 35216 29464 37136 29492
rect 35216 29452 35222 29464
rect 37182 29452 37188 29504
rect 37240 29492 37246 29504
rect 37461 29495 37519 29501
rect 37461 29492 37473 29495
rect 37240 29464 37473 29492
rect 37240 29452 37246 29464
rect 37461 29461 37473 29464
rect 37507 29461 37519 29495
rect 37461 29455 37519 29461
rect 39298 29452 39304 29504
rect 39356 29492 39362 29504
rect 39485 29495 39543 29501
rect 39485 29492 39497 29495
rect 39356 29464 39497 29492
rect 39356 29452 39362 29464
rect 39485 29461 39497 29464
rect 39531 29461 39543 29495
rect 39485 29455 39543 29461
rect 39574 29452 39580 29504
rect 39632 29492 39638 29504
rect 42061 29495 42119 29501
rect 42061 29492 42073 29495
rect 39632 29464 42073 29492
rect 39632 29452 39638 29464
rect 42061 29461 42073 29464
rect 42107 29461 42119 29495
rect 42061 29455 42119 29461
rect 1104 29402 43884 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 43884 29402
rect 1104 29328 43884 29350
rect 12802 29248 12808 29300
rect 12860 29288 12866 29300
rect 13541 29291 13599 29297
rect 13541 29288 13553 29291
rect 12860 29260 13553 29288
rect 12860 29248 12866 29260
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 12636 29084 12664 29115
rect 12894 29112 12900 29164
rect 12952 29112 12958 29164
rect 13004 29161 13032 29260
rect 13541 29257 13553 29260
rect 13587 29288 13599 29291
rect 14274 29288 14280 29300
rect 13587 29260 14280 29288
rect 13587 29257 13599 29260
rect 13541 29251 13599 29257
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 16390 29248 16396 29300
rect 16448 29288 16454 29300
rect 16945 29291 17003 29297
rect 16945 29288 16957 29291
rect 16448 29260 16957 29288
rect 16448 29248 16454 29260
rect 16945 29257 16957 29260
rect 16991 29257 17003 29291
rect 18046 29288 18052 29300
rect 16945 29251 17003 29257
rect 17236 29260 18052 29288
rect 13906 29180 13912 29232
rect 13964 29180 13970 29232
rect 15013 29223 15071 29229
rect 15013 29189 15025 29223
rect 15059 29220 15071 29223
rect 15194 29220 15200 29232
rect 15059 29192 15200 29220
rect 15059 29189 15071 29192
rect 15013 29183 15071 29189
rect 15194 29180 15200 29192
rect 15252 29180 15258 29232
rect 12989 29155 13047 29161
rect 12989 29121 13001 29155
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 13630 29112 13636 29164
rect 13688 29152 13694 29164
rect 13725 29155 13783 29161
rect 13725 29152 13737 29155
rect 13688 29124 13737 29152
rect 13688 29112 13694 29124
rect 13725 29121 13737 29124
rect 13771 29121 13783 29155
rect 13725 29115 13783 29121
rect 13740 29084 13768 29115
rect 14826 29112 14832 29164
rect 14884 29112 14890 29164
rect 15105 29155 15163 29161
rect 15105 29121 15117 29155
rect 15151 29152 15163 29155
rect 15286 29152 15292 29164
rect 15151 29124 15292 29152
rect 15151 29121 15163 29124
rect 15105 29115 15163 29121
rect 15286 29112 15292 29124
rect 15344 29152 15350 29164
rect 15657 29155 15715 29161
rect 15657 29152 15669 29155
rect 15344 29124 15669 29152
rect 15344 29112 15350 29124
rect 15657 29121 15669 29124
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 15838 29112 15844 29164
rect 15896 29112 15902 29164
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29121 15991 29155
rect 15933 29115 15991 29121
rect 15948 29084 15976 29115
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 16206 29112 16212 29164
rect 16264 29152 16270 29164
rect 16850 29152 16856 29164
rect 16264 29124 16856 29152
rect 16264 29112 16270 29124
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 17129 29155 17187 29161
rect 17129 29121 17141 29155
rect 17175 29152 17187 29155
rect 17236 29152 17264 29260
rect 18046 29248 18052 29260
rect 18104 29248 18110 29300
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18196 29260 18397 29288
rect 18196 29248 18202 29260
rect 17862 29180 17868 29232
rect 17920 29220 17926 29232
rect 17920 29192 18092 29220
rect 17920 29180 17926 29192
rect 18064 29161 18092 29192
rect 18369 29174 18397 29260
rect 18966 29248 18972 29300
rect 19024 29288 19030 29300
rect 19521 29291 19579 29297
rect 19521 29288 19533 29291
rect 19024 29260 19533 29288
rect 19024 29248 19030 29260
rect 19521 29257 19533 29260
rect 19567 29257 19579 29291
rect 19521 29251 19579 29257
rect 20070 29248 20076 29300
rect 20128 29248 20134 29300
rect 20530 29288 20536 29300
rect 20272 29260 20536 29288
rect 18598 29180 18604 29232
rect 18656 29220 18662 29232
rect 19978 29220 19984 29232
rect 18656 29192 19984 29220
rect 18656 29180 18662 29192
rect 19978 29180 19984 29192
rect 20036 29180 20042 29232
rect 18245 29161 18397 29174
rect 17175 29124 17264 29152
rect 17957 29155 18015 29161
rect 17175 29121 17187 29124
rect 17129 29115 17187 29121
rect 17957 29121 17969 29155
rect 18003 29121 18015 29155
rect 17957 29115 18015 29121
rect 18049 29155 18107 29161
rect 18049 29121 18061 29155
rect 18095 29121 18107 29155
rect 18049 29115 18107 29121
rect 18233 29155 18397 29161
rect 18233 29121 18245 29155
rect 18279 29146 18397 29155
rect 18279 29121 18291 29146
rect 18233 29115 18291 29121
rect 16758 29084 16764 29096
rect 12636 29056 13216 29084
rect 13740 29056 14964 29084
rect 15948 29056 16764 29084
rect 13188 29028 13216 29056
rect 12713 29019 12771 29025
rect 12713 28985 12725 29019
rect 12759 29016 12771 29019
rect 12986 29016 12992 29028
rect 12759 28988 12992 29016
rect 12759 28985 12771 28988
rect 12713 28979 12771 28985
rect 12986 28976 12992 28988
rect 13044 28976 13050 29028
rect 13170 28976 13176 29028
rect 13228 29016 13234 29028
rect 14829 29019 14887 29025
rect 14829 29016 14841 29019
rect 13228 28988 14841 29016
rect 13228 28976 13234 28988
rect 14829 28985 14841 28988
rect 14875 28985 14887 29019
rect 14936 29016 14964 29056
rect 16758 29044 16764 29056
rect 16816 29044 16822 29096
rect 16942 29044 16948 29096
rect 17000 29084 17006 29096
rect 17972 29084 18000 29115
rect 18966 29112 18972 29164
rect 19024 29112 19030 29164
rect 19426 29112 19432 29164
rect 19484 29112 19490 29164
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29152 19671 29155
rect 20272 29152 20300 29260
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 21450 29248 21456 29300
rect 21508 29248 21514 29300
rect 22186 29248 22192 29300
rect 22244 29288 22250 29300
rect 22833 29291 22891 29297
rect 22833 29288 22845 29291
rect 22244 29260 22845 29288
rect 22244 29248 22250 29260
rect 22833 29257 22845 29260
rect 22879 29257 22891 29291
rect 22833 29251 22891 29257
rect 23201 29291 23259 29297
rect 23201 29257 23213 29291
rect 23247 29288 23259 29291
rect 23474 29288 23480 29300
rect 23247 29260 23480 29288
rect 23247 29257 23259 29260
rect 23201 29251 23259 29257
rect 23474 29248 23480 29260
rect 23532 29248 23538 29300
rect 25130 29248 25136 29300
rect 25188 29248 25194 29300
rect 26605 29291 26663 29297
rect 26605 29257 26617 29291
rect 26651 29257 26663 29291
rect 26605 29251 26663 29257
rect 20346 29180 20352 29232
rect 20404 29220 20410 29232
rect 20404 29192 22094 29220
rect 20404 29180 20410 29192
rect 19659 29124 20300 29152
rect 20441 29155 20499 29161
rect 19659 29121 19671 29124
rect 19613 29115 19671 29121
rect 20441 29121 20453 29155
rect 20487 29152 20499 29155
rect 20530 29152 20536 29164
rect 20487 29124 20536 29152
rect 20487 29121 20499 29124
rect 20441 29115 20499 29121
rect 18138 29084 18144 29096
rect 17000 29056 18144 29084
rect 17000 29044 17006 29056
rect 18138 29044 18144 29056
rect 18196 29044 18202 29096
rect 18354 29087 18412 29093
rect 18354 29053 18366 29087
rect 18400 29084 18412 29087
rect 19334 29084 19340 29096
rect 18400 29056 19340 29084
rect 18400 29053 18412 29056
rect 18354 29047 18412 29053
rect 19334 29044 19340 29056
rect 19392 29044 19398 29096
rect 19444 29084 19472 29112
rect 20254 29084 20260 29096
rect 19444 29056 20260 29084
rect 20254 29044 20260 29056
rect 20312 29084 20318 29096
rect 20456 29084 20484 29115
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 22066 29152 22094 29192
rect 22738 29180 22744 29232
rect 22796 29220 22802 29232
rect 23845 29223 23903 29229
rect 23845 29220 23857 29223
rect 22796 29192 23857 29220
rect 22796 29180 22802 29192
rect 23845 29189 23857 29192
rect 23891 29220 23903 29223
rect 24854 29220 24860 29232
rect 23891 29192 24860 29220
rect 23891 29189 23903 29192
rect 23845 29183 23903 29189
rect 24854 29180 24860 29192
rect 24912 29180 24918 29232
rect 26620 29220 26648 29251
rect 28350 29248 28356 29300
rect 28408 29288 28414 29300
rect 28537 29291 28595 29297
rect 28537 29288 28549 29291
rect 28408 29260 28549 29288
rect 28408 29248 28414 29260
rect 28537 29257 28549 29260
rect 28583 29257 28595 29291
rect 28537 29251 28595 29257
rect 29365 29291 29423 29297
rect 29365 29257 29377 29291
rect 29411 29288 29423 29291
rect 29638 29288 29644 29300
rect 29411 29260 29644 29288
rect 29411 29257 29423 29260
rect 29365 29251 29423 29257
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 30006 29248 30012 29300
rect 30064 29248 30070 29300
rect 31110 29288 31116 29300
rect 30116 29260 31116 29288
rect 27402 29223 27460 29229
rect 27402 29220 27414 29223
rect 26620 29192 27414 29220
rect 27402 29189 27414 29192
rect 27448 29189 27460 29223
rect 27402 29183 27460 29189
rect 29454 29180 29460 29232
rect 29512 29220 29518 29232
rect 30116 29220 30144 29260
rect 29512 29192 30144 29220
rect 30193 29223 30251 29229
rect 29512 29180 29518 29192
rect 30193 29189 30205 29223
rect 30239 29220 30251 29223
rect 30650 29220 30656 29232
rect 30239 29192 30656 29220
rect 30239 29189 30251 29192
rect 30193 29183 30251 29189
rect 30650 29180 30656 29192
rect 30708 29180 30714 29232
rect 22281 29155 22339 29161
rect 22281 29152 22293 29155
rect 22066 29124 22293 29152
rect 22281 29121 22293 29124
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 20312 29056 20484 29084
rect 20312 29044 20318 29056
rect 20622 29044 20628 29096
rect 20680 29044 20686 29096
rect 22296 29084 22324 29115
rect 23014 29112 23020 29164
rect 23072 29112 23078 29164
rect 23290 29112 23296 29164
rect 23348 29112 23354 29164
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29121 24363 29155
rect 24305 29115 24363 29121
rect 23842 29084 23848 29096
rect 22296 29056 23848 29084
rect 23842 29044 23848 29056
rect 23900 29044 23906 29096
rect 24320 29084 24348 29115
rect 24394 29112 24400 29164
rect 24452 29112 24458 29164
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29152 24639 29155
rect 25038 29152 25044 29164
rect 24627 29124 25044 29152
rect 24627 29121 24639 29124
rect 24581 29115 24639 29121
rect 25038 29112 25044 29124
rect 25096 29112 25102 29164
rect 25314 29112 25320 29164
rect 25372 29152 25378 29164
rect 25409 29155 25467 29161
rect 25409 29152 25421 29155
rect 25372 29124 25421 29152
rect 25372 29112 25378 29124
rect 25409 29121 25421 29124
rect 25455 29121 25467 29155
rect 25409 29115 25467 29121
rect 26418 29112 26424 29164
rect 26476 29112 26482 29164
rect 28994 29152 29000 29164
rect 26712 29124 29000 29152
rect 24762 29084 24768 29096
rect 24320 29056 24768 29084
rect 24762 29044 24768 29056
rect 24820 29084 24826 29096
rect 25590 29084 25596 29096
rect 24820 29056 25596 29084
rect 24820 29044 24826 29056
rect 25590 29044 25596 29056
rect 25648 29084 25654 29096
rect 26712 29084 26740 29124
rect 28966 29112 29000 29124
rect 29052 29112 29058 29164
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 25648 29056 26740 29084
rect 25648 29044 25654 29056
rect 26786 29044 26792 29096
rect 26844 29084 26850 29096
rect 27157 29087 27215 29093
rect 27157 29084 27169 29087
rect 26844 29056 27169 29084
rect 26844 29044 26850 29056
rect 27157 29053 27169 29056
rect 27203 29053 27215 29087
rect 27157 29047 27215 29053
rect 21910 29016 21916 29028
rect 14936 28988 21916 29016
rect 14829 28979 14887 28985
rect 21910 28976 21916 28988
rect 21968 28976 21974 29028
rect 22097 29019 22155 29025
rect 22097 28985 22109 29019
rect 22143 29016 22155 29019
rect 22554 29016 22560 29028
rect 22143 28988 22560 29016
rect 22143 28985 22155 28988
rect 22097 28979 22155 28985
rect 22554 28976 22560 28988
rect 22612 28976 22618 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 24581 29019 24639 29025
rect 24581 29016 24593 29019
rect 23440 28988 24593 29016
rect 23440 28976 23446 28988
rect 24581 28985 24593 28988
rect 24627 28985 24639 29019
rect 28966 29016 28994 29112
rect 29564 29084 29592 29115
rect 30282 29112 30288 29164
rect 30340 29152 30346 29164
rect 30377 29155 30435 29161
rect 30377 29152 30389 29155
rect 30340 29124 30389 29152
rect 30340 29112 30346 29124
rect 30377 29121 30389 29124
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 30837 29155 30895 29161
rect 30837 29121 30849 29155
rect 30883 29152 30895 29155
rect 30926 29152 30932 29164
rect 30883 29124 30932 29152
rect 30883 29121 30895 29124
rect 30837 29115 30895 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31036 29161 31064 29260
rect 31110 29248 31116 29260
rect 31168 29248 31174 29300
rect 31202 29248 31208 29300
rect 31260 29248 31266 29300
rect 32214 29248 32220 29300
rect 32272 29288 32278 29300
rect 32309 29291 32367 29297
rect 32309 29288 32321 29291
rect 32272 29260 32321 29288
rect 32272 29248 32278 29260
rect 32309 29257 32321 29260
rect 32355 29257 32367 29291
rect 32309 29251 32367 29257
rect 34698 29248 34704 29300
rect 34756 29248 34762 29300
rect 34793 29291 34851 29297
rect 34793 29257 34805 29291
rect 34839 29288 34851 29291
rect 35158 29288 35164 29300
rect 34839 29260 35164 29288
rect 34839 29257 34851 29260
rect 34793 29251 34851 29257
rect 35158 29248 35164 29260
rect 35216 29248 35222 29300
rect 36633 29291 36691 29297
rect 36633 29257 36645 29291
rect 36679 29288 36691 29291
rect 36998 29288 37004 29300
rect 36679 29260 37004 29288
rect 36679 29257 36691 29260
rect 36633 29251 36691 29257
rect 36998 29248 37004 29260
rect 37056 29248 37062 29300
rect 37366 29248 37372 29300
rect 37424 29288 37430 29300
rect 37553 29291 37611 29297
rect 37553 29288 37565 29291
rect 37424 29260 37565 29288
rect 37424 29248 37430 29260
rect 37553 29257 37565 29260
rect 37599 29257 37611 29291
rect 37553 29251 37611 29257
rect 37918 29248 37924 29300
rect 37976 29288 37982 29300
rect 40221 29291 40279 29297
rect 37976 29260 39436 29288
rect 37976 29248 37982 29260
rect 34514 29220 34520 29232
rect 34164 29192 34520 29220
rect 31021 29155 31079 29161
rect 31021 29121 31033 29155
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 32490 29112 32496 29164
rect 32548 29112 32554 29164
rect 32674 29112 32680 29164
rect 32732 29112 32738 29164
rect 33321 29155 33379 29161
rect 33321 29121 33333 29155
rect 33367 29152 33379 29155
rect 33410 29152 33416 29164
rect 33367 29124 33416 29152
rect 33367 29121 33379 29124
rect 33321 29115 33379 29121
rect 33410 29112 33416 29124
rect 33468 29152 33474 29164
rect 33594 29152 33600 29164
rect 33468 29124 33600 29152
rect 33468 29112 33474 29124
rect 33594 29112 33600 29124
rect 33652 29112 33658 29164
rect 34164 29161 34192 29192
rect 34514 29180 34520 29192
rect 34572 29180 34578 29232
rect 34716 29220 34744 29248
rect 34882 29220 34888 29232
rect 34624 29192 34888 29220
rect 34149 29155 34207 29161
rect 34149 29121 34161 29155
rect 34195 29121 34207 29155
rect 34149 29115 34207 29121
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29152 34391 29155
rect 34422 29152 34428 29164
rect 34379 29124 34428 29152
rect 34379 29121 34391 29124
rect 34333 29115 34391 29121
rect 34422 29112 34428 29124
rect 34480 29112 34486 29164
rect 34624 29161 34652 29192
rect 34882 29180 34888 29192
rect 34940 29180 34946 29232
rect 35253 29223 35311 29229
rect 35253 29189 35265 29223
rect 35299 29220 35311 29223
rect 35342 29220 35348 29232
rect 35299 29192 35348 29220
rect 35299 29189 35311 29192
rect 35253 29183 35311 29189
rect 35342 29180 35348 29192
rect 35400 29180 35406 29232
rect 38194 29220 38200 29232
rect 36648 29192 38200 29220
rect 34609 29155 34667 29161
rect 34609 29121 34621 29155
rect 34655 29121 34667 29155
rect 34609 29115 34667 29121
rect 34698 29112 34704 29164
rect 34756 29152 34762 29164
rect 36648 29161 36676 29192
rect 38194 29180 38200 29192
rect 38252 29180 38258 29232
rect 38470 29180 38476 29232
rect 38528 29180 38534 29232
rect 39408 29220 39436 29260
rect 40221 29257 40233 29291
rect 40267 29288 40279 29291
rect 41046 29288 41052 29300
rect 40267 29260 41052 29288
rect 40267 29257 40279 29260
rect 40221 29251 40279 29257
rect 41046 29248 41052 29260
rect 41104 29248 41110 29300
rect 41138 29248 41144 29300
rect 41196 29288 41202 29300
rect 42613 29291 42671 29297
rect 42613 29288 42625 29291
rect 41196 29260 42625 29288
rect 41196 29248 41202 29260
rect 42613 29257 42625 29260
rect 42659 29257 42671 29291
rect 42613 29251 42671 29257
rect 39574 29220 39580 29232
rect 39408 29192 39580 29220
rect 35529 29155 35587 29161
rect 35529 29152 35541 29155
rect 34756 29124 35541 29152
rect 34756 29112 34762 29124
rect 35529 29121 35541 29124
rect 35575 29121 35587 29155
rect 35529 29115 35587 29121
rect 36633 29155 36691 29161
rect 36633 29121 36645 29155
rect 36679 29121 36691 29155
rect 36633 29115 36691 29121
rect 36909 29155 36967 29161
rect 36909 29121 36921 29155
rect 36955 29152 36967 29155
rect 37921 29155 37979 29161
rect 37921 29152 37933 29155
rect 36955 29124 37933 29152
rect 36955 29121 36967 29124
rect 36909 29115 36967 29121
rect 37921 29121 37933 29124
rect 37967 29152 37979 29155
rect 38102 29152 38108 29164
rect 37967 29124 38108 29152
rect 37967 29121 37979 29124
rect 37921 29115 37979 29121
rect 38102 29112 38108 29124
rect 38160 29112 38166 29164
rect 38562 29112 38568 29164
rect 38620 29152 38626 29164
rect 39408 29161 39436 29192
rect 39574 29180 39580 29192
rect 39632 29180 39638 29232
rect 40310 29180 40316 29232
rect 40368 29220 40374 29232
rect 40770 29220 40776 29232
rect 40368 29192 40776 29220
rect 40368 29180 40374 29192
rect 40770 29180 40776 29192
rect 40828 29180 40834 29232
rect 39301 29155 39359 29161
rect 39301 29152 39313 29155
rect 38620 29124 39313 29152
rect 38620 29112 38626 29124
rect 39301 29121 39313 29124
rect 39347 29121 39359 29155
rect 39301 29115 39359 29121
rect 39393 29155 39451 29161
rect 39393 29121 39405 29155
rect 39439 29121 39451 29155
rect 39393 29115 39451 29121
rect 31662 29084 31668 29096
rect 29564 29056 31668 29084
rect 31662 29044 31668 29056
rect 31720 29044 31726 29096
rect 31754 29044 31760 29096
rect 31812 29044 31818 29096
rect 31938 29044 31944 29096
rect 31996 29084 32002 29096
rect 35345 29087 35403 29093
rect 35345 29084 35357 29087
rect 31996 29056 35357 29084
rect 31996 29044 32002 29056
rect 35345 29053 35357 29056
rect 35391 29053 35403 29087
rect 35345 29047 35403 29053
rect 37734 29044 37740 29096
rect 37792 29084 37798 29096
rect 37829 29087 37887 29093
rect 37829 29084 37841 29087
rect 37792 29056 37841 29084
rect 37792 29044 37798 29056
rect 37829 29053 37841 29056
rect 37875 29053 37887 29087
rect 38930 29084 38936 29096
rect 37829 29047 37887 29053
rect 37936 29056 38936 29084
rect 29822 29016 29828 29028
rect 28966 28988 29828 29016
rect 24581 28979 24639 28985
rect 29822 28976 29828 28988
rect 29880 29016 29886 29028
rect 31956 29016 31984 29044
rect 29880 28988 31984 29016
rect 29880 28976 29886 28988
rect 33502 28976 33508 29028
rect 33560 28976 33566 29028
rect 33870 28976 33876 29028
rect 33928 29016 33934 29028
rect 34425 29019 34483 29025
rect 34425 29016 34437 29019
rect 33928 28988 34437 29016
rect 33928 28976 33934 28988
rect 34425 28985 34437 28988
rect 34471 28985 34483 29019
rect 34425 28979 34483 28985
rect 34517 29019 34575 29025
rect 34517 28985 34529 29019
rect 34563 29016 34575 29019
rect 34563 28988 34597 29016
rect 34563 28985 34575 28988
rect 34517 28979 34575 28985
rect 13078 28908 13084 28960
rect 13136 28948 13142 28960
rect 13446 28948 13452 28960
rect 13136 28920 13452 28948
rect 13136 28908 13142 28920
rect 13446 28908 13452 28920
rect 13504 28908 13510 28960
rect 18414 28908 18420 28960
rect 18472 28908 18478 28960
rect 25866 28908 25872 28960
rect 25924 28948 25930 28960
rect 29178 28948 29184 28960
rect 25924 28920 29184 28948
rect 25924 28908 25930 28920
rect 29178 28908 29184 28920
rect 29236 28908 29242 28960
rect 29270 28908 29276 28960
rect 29328 28948 29334 28960
rect 31570 28948 31576 28960
rect 29328 28920 31576 28948
rect 29328 28908 29334 28920
rect 31570 28908 31576 28920
rect 31628 28908 31634 28960
rect 34146 28908 34152 28960
rect 34204 28948 34210 28960
rect 34532 28948 34560 28979
rect 34882 28976 34888 29028
rect 34940 29016 34946 29028
rect 35618 29016 35624 29028
rect 34940 28988 35624 29016
rect 34940 28976 34946 28988
rect 35618 28976 35624 28988
rect 35676 28976 35682 29028
rect 35713 29019 35771 29025
rect 35713 28985 35725 29019
rect 35759 29016 35771 29019
rect 35894 29016 35900 29028
rect 35759 28988 35900 29016
rect 35759 28985 35771 28988
rect 35713 28979 35771 28985
rect 35894 28976 35900 28988
rect 35952 28976 35958 29028
rect 36725 29019 36783 29025
rect 36725 28985 36737 29019
rect 36771 29016 36783 29019
rect 37936 29016 37964 29056
rect 38930 29044 38936 29056
rect 38988 29044 38994 29096
rect 39022 29044 39028 29096
rect 39080 29044 39086 29096
rect 39316 29084 39344 29115
rect 39482 29112 39488 29164
rect 39540 29112 39546 29164
rect 39666 29112 39672 29164
rect 39724 29112 39730 29164
rect 40402 29112 40408 29164
rect 40460 29152 40466 29164
rect 41046 29152 41052 29164
rect 40460 29124 41052 29152
rect 40460 29112 40466 29124
rect 41046 29112 41052 29124
rect 41104 29112 41110 29164
rect 41414 29112 41420 29164
rect 41472 29152 41478 29164
rect 41601 29155 41659 29161
rect 41601 29152 41613 29155
rect 41472 29124 41613 29152
rect 41472 29112 41478 29124
rect 41601 29121 41613 29124
rect 41647 29152 41659 29155
rect 41647 29124 42104 29152
rect 41647 29121 41659 29124
rect 41601 29115 41659 29121
rect 39574 29084 39580 29096
rect 39316 29056 39580 29084
rect 39574 29044 39580 29056
rect 39632 29044 39638 29096
rect 40954 29044 40960 29096
rect 41012 29044 41018 29096
rect 41141 29087 41199 29093
rect 41141 29053 41153 29087
rect 41187 29084 41199 29087
rect 41187 29056 41414 29084
rect 41187 29053 41199 29056
rect 41141 29047 41199 29053
rect 36771 28988 37964 29016
rect 36771 28985 36783 28988
rect 36725 28979 36783 28985
rect 38470 28976 38476 29028
rect 38528 29016 38534 29028
rect 40586 29016 40592 29028
rect 38528 28988 40592 29016
rect 38528 28976 38534 28988
rect 40586 28976 40592 28988
rect 40644 28976 40650 29028
rect 34204 28920 34560 28948
rect 34204 28908 34210 28920
rect 35526 28908 35532 28960
rect 35584 28948 35590 28960
rect 37274 28948 37280 28960
rect 35584 28920 37280 28948
rect 35584 28908 35590 28920
rect 37274 28908 37280 28920
rect 37332 28908 37338 28960
rect 37921 28951 37979 28957
rect 37921 28917 37933 28951
rect 37967 28948 37979 28951
rect 40494 28948 40500 28960
rect 37967 28920 40500 28948
rect 37967 28917 37979 28920
rect 37921 28911 37979 28917
rect 40494 28908 40500 28920
rect 40552 28908 40558 28960
rect 41046 28908 41052 28960
rect 41104 28948 41110 28960
rect 41233 28951 41291 28957
rect 41233 28948 41245 28951
rect 41104 28920 41245 28948
rect 41104 28908 41110 28920
rect 41233 28917 41245 28920
rect 41279 28917 41291 28951
rect 41386 28948 41414 29056
rect 41506 29044 41512 29096
rect 41564 29084 41570 29096
rect 41693 29087 41751 29093
rect 41693 29084 41705 29087
rect 41564 29056 41705 29084
rect 41564 29044 41570 29056
rect 41693 29053 41705 29056
rect 41739 29084 41751 29087
rect 42076 29084 42104 29124
rect 42242 29112 42248 29164
rect 42300 29152 42306 29164
rect 42981 29155 43039 29161
rect 42981 29152 42993 29155
rect 42300 29124 42993 29152
rect 42300 29112 42306 29124
rect 42981 29121 42993 29124
rect 43027 29121 43039 29155
rect 42981 29115 43039 29121
rect 42889 29087 42947 29093
rect 42889 29084 42901 29087
rect 41739 29056 42012 29084
rect 42076 29056 42901 29084
rect 41739 29053 41751 29056
rect 41693 29047 41751 29053
rect 41984 28960 42012 29056
rect 42889 29053 42901 29056
rect 42935 29053 42947 29087
rect 42889 29047 42947 29053
rect 41874 28948 41880 28960
rect 41386 28920 41880 28948
rect 41233 28911 41291 28917
rect 41874 28908 41880 28920
rect 41932 28908 41938 28960
rect 41966 28908 41972 28960
rect 42024 28948 42030 28960
rect 42797 28951 42855 28957
rect 42797 28948 42809 28951
rect 42024 28920 42809 28948
rect 42024 28908 42030 28920
rect 42797 28917 42809 28920
rect 42843 28917 42855 28951
rect 42797 28911 42855 28917
rect 1104 28858 43884 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 43884 28858
rect 1104 28784 43884 28806
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 15197 28747 15255 28753
rect 15197 28744 15209 28747
rect 14884 28716 15209 28744
rect 14884 28704 14890 28716
rect 15197 28713 15209 28716
rect 15243 28744 15255 28747
rect 15749 28747 15807 28753
rect 15749 28744 15761 28747
rect 15243 28716 15761 28744
rect 15243 28713 15255 28716
rect 15197 28707 15255 28713
rect 15749 28713 15761 28716
rect 15795 28713 15807 28747
rect 15749 28707 15807 28713
rect 16114 28704 16120 28756
rect 16172 28704 16178 28756
rect 16758 28704 16764 28756
rect 16816 28704 16822 28756
rect 17236 28716 18552 28744
rect 13173 28679 13231 28685
rect 13173 28645 13185 28679
rect 13219 28676 13231 28679
rect 13354 28676 13360 28688
rect 13219 28648 13360 28676
rect 13219 28645 13231 28648
rect 13173 28639 13231 28645
rect 13354 28636 13360 28648
rect 13412 28636 13418 28688
rect 13725 28679 13783 28685
rect 13725 28645 13737 28679
rect 13771 28676 13783 28679
rect 16022 28676 16028 28688
rect 13771 28648 16028 28676
rect 13771 28645 13783 28648
rect 13725 28639 13783 28645
rect 16022 28636 16028 28648
rect 16080 28676 16086 28688
rect 17236 28676 17264 28716
rect 18414 28676 18420 28688
rect 16080 28648 17264 28676
rect 17696 28648 18420 28676
rect 16080 28636 16086 28648
rect 16206 28568 16212 28620
rect 16264 28568 16270 28620
rect 17310 28568 17316 28620
rect 17368 28608 17374 28620
rect 17696 28617 17724 28648
rect 18414 28636 18420 28648
rect 18472 28636 18478 28688
rect 18524 28676 18552 28716
rect 19334 28704 19340 28756
rect 19392 28744 19398 28756
rect 19429 28747 19487 28753
rect 19429 28744 19441 28747
rect 19392 28716 19441 28744
rect 19392 28704 19398 28716
rect 19429 28713 19441 28716
rect 19475 28713 19487 28747
rect 19429 28707 19487 28713
rect 20162 28704 20168 28756
rect 20220 28744 20226 28756
rect 20257 28747 20315 28753
rect 20257 28744 20269 28747
rect 20220 28716 20269 28744
rect 20220 28704 20226 28716
rect 20257 28713 20269 28716
rect 20303 28713 20315 28747
rect 28350 28744 28356 28756
rect 20257 28707 20315 28713
rect 26436 28716 28356 28744
rect 20714 28676 20720 28688
rect 18524 28648 20720 28676
rect 20714 28636 20720 28648
rect 20772 28636 20778 28688
rect 21821 28679 21879 28685
rect 21821 28676 21833 28679
rect 20916 28648 21833 28676
rect 20916 28620 20944 28648
rect 21821 28645 21833 28648
rect 21867 28645 21879 28679
rect 25866 28676 25872 28688
rect 21821 28639 21879 28645
rect 22066 28648 25872 28676
rect 17497 28611 17555 28617
rect 17497 28608 17509 28611
rect 17368 28580 17509 28608
rect 17368 28568 17374 28580
rect 17497 28577 17509 28580
rect 17543 28577 17555 28611
rect 17497 28571 17555 28577
rect 17681 28611 17739 28617
rect 17681 28577 17693 28611
rect 17727 28577 17739 28611
rect 17681 28571 17739 28577
rect 17773 28611 17831 28617
rect 17773 28577 17785 28611
rect 17819 28608 17831 28611
rect 17954 28608 17960 28620
rect 17819 28580 17960 28608
rect 17819 28577 17831 28580
rect 17773 28571 17831 28577
rect 17954 28568 17960 28580
rect 18012 28608 18018 28620
rect 18785 28611 18843 28617
rect 18785 28608 18797 28611
rect 18012 28580 18797 28608
rect 18012 28568 18018 28580
rect 18785 28577 18797 28580
rect 18831 28577 18843 28611
rect 20898 28608 20904 28620
rect 18785 28571 18843 28577
rect 19812 28580 20904 28608
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 12897 28475 12955 28481
rect 12897 28441 12909 28475
rect 12943 28441 12955 28475
rect 13280 28472 13308 28503
rect 13446 28500 13452 28552
rect 13504 28500 13510 28552
rect 15286 28500 15292 28552
rect 15344 28500 15350 28552
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 15933 28543 15991 28549
rect 15933 28540 15945 28543
rect 15896 28512 15945 28540
rect 15896 28500 15902 28512
rect 15933 28509 15945 28512
rect 15979 28509 15991 28543
rect 15933 28503 15991 28509
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 16942 28540 16948 28552
rect 16899 28512 16948 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28540 17647 28543
rect 18046 28540 18052 28552
rect 17635 28512 18052 28540
rect 17635 28509 17647 28512
rect 17589 28503 17647 28509
rect 18046 28500 18052 28512
rect 18104 28540 18110 28552
rect 18506 28540 18512 28552
rect 18104 28512 18512 28540
rect 18104 28500 18110 28512
rect 18506 28500 18512 28512
rect 18564 28500 18570 28552
rect 19812 28549 19840 28580
rect 20898 28568 20904 28580
rect 20956 28568 20962 28620
rect 22066 28608 22094 28648
rect 25866 28636 25872 28648
rect 25924 28636 25930 28688
rect 23382 28608 23388 28620
rect 21836 28580 22094 28608
rect 22848 28580 23388 28608
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 20036 28512 20453 28540
rect 20036 28500 20042 28512
rect 20441 28509 20453 28512
rect 20487 28509 20499 28543
rect 20441 28503 20499 28509
rect 20530 28500 20536 28552
rect 20588 28500 20594 28552
rect 21836 28549 21864 28580
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28509 21879 28543
rect 21821 28503 21879 28509
rect 22097 28543 22155 28549
rect 22097 28509 22109 28543
rect 22143 28540 22155 28543
rect 22186 28540 22192 28552
rect 22143 28512 22192 28540
rect 22143 28509 22155 28512
rect 22097 28503 22155 28509
rect 22186 28500 22192 28512
rect 22244 28500 22250 28552
rect 22848 28549 22876 28580
rect 23382 28568 23388 28580
rect 23440 28568 23446 28620
rect 26053 28611 26111 28617
rect 26053 28577 26065 28611
rect 26099 28608 26111 28611
rect 26326 28608 26332 28620
rect 26099 28580 26332 28608
rect 26099 28577 26111 28580
rect 26053 28571 26111 28577
rect 26326 28568 26332 28580
rect 26384 28568 26390 28620
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28540 23535 28543
rect 23566 28540 23572 28552
rect 23523 28512 23572 28540
rect 23523 28509 23535 28512
rect 23477 28503 23535 28509
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 26237 28543 26295 28549
rect 26237 28509 26249 28543
rect 26283 28540 26295 28543
rect 26436 28540 26464 28716
rect 28350 28704 28356 28716
rect 28408 28704 28414 28756
rect 30101 28747 30159 28753
rect 30101 28713 30113 28747
rect 30147 28744 30159 28747
rect 30282 28744 30288 28756
rect 30147 28716 30288 28744
rect 30147 28713 30159 28716
rect 30101 28707 30159 28713
rect 30282 28704 30288 28716
rect 30340 28704 30346 28756
rect 31386 28704 31392 28756
rect 31444 28744 31450 28756
rect 33778 28744 33784 28756
rect 31444 28716 33784 28744
rect 31444 28704 31450 28716
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 34054 28704 34060 28756
rect 34112 28744 34118 28756
rect 34885 28747 34943 28753
rect 34885 28744 34897 28747
rect 34112 28716 34897 28744
rect 34112 28704 34118 28716
rect 34885 28713 34897 28716
rect 34931 28713 34943 28747
rect 34885 28707 34943 28713
rect 35342 28704 35348 28756
rect 35400 28704 35406 28756
rect 35894 28704 35900 28756
rect 35952 28704 35958 28756
rect 36725 28747 36783 28753
rect 36725 28713 36737 28747
rect 36771 28744 36783 28747
rect 36998 28744 37004 28756
rect 36771 28716 37004 28744
rect 36771 28713 36783 28716
rect 36725 28707 36783 28713
rect 36998 28704 37004 28716
rect 37056 28704 37062 28756
rect 37550 28704 37556 28756
rect 37608 28744 37614 28756
rect 38013 28747 38071 28753
rect 38013 28744 38025 28747
rect 37608 28716 38025 28744
rect 37608 28704 37614 28716
rect 38013 28713 38025 28716
rect 38059 28744 38071 28747
rect 38746 28744 38752 28756
rect 38059 28716 38752 28744
rect 38059 28713 38071 28716
rect 38013 28707 38071 28713
rect 38746 28704 38752 28716
rect 38804 28704 38810 28756
rect 26510 28636 26516 28688
rect 26568 28676 26574 28688
rect 26568 28648 26832 28676
rect 26568 28636 26574 28648
rect 26694 28568 26700 28620
rect 26752 28568 26758 28620
rect 26804 28608 26832 28648
rect 27706 28636 27712 28688
rect 27764 28676 27770 28688
rect 31478 28676 31484 28688
rect 27764 28648 31484 28676
rect 27764 28636 27770 28648
rect 28920 28617 28948 28648
rect 31478 28636 31484 28648
rect 31536 28636 31542 28688
rect 31570 28636 31576 28688
rect 31628 28676 31634 28688
rect 36265 28679 36323 28685
rect 31628 28648 32628 28676
rect 31628 28636 31634 28648
rect 27249 28611 27307 28617
rect 27249 28608 27261 28611
rect 26804 28580 27261 28608
rect 27249 28577 27261 28580
rect 27295 28577 27307 28611
rect 27249 28571 27307 28577
rect 28905 28611 28963 28617
rect 28905 28577 28917 28611
rect 28951 28577 28963 28611
rect 28905 28571 28963 28577
rect 30742 28568 30748 28620
rect 30800 28568 30806 28620
rect 30834 28568 30840 28620
rect 30892 28608 30898 28620
rect 32600 28617 32628 28648
rect 32876 28648 36124 28676
rect 32585 28611 32643 28617
rect 30892 28580 32352 28608
rect 30892 28568 30898 28580
rect 26283 28512 26464 28540
rect 26283 28509 26295 28512
rect 26237 28503 26295 28509
rect 26970 28500 26976 28552
rect 27028 28500 27034 28552
rect 27062 28500 27068 28552
rect 27120 28549 27126 28552
rect 27120 28543 27148 28549
rect 27136 28509 27148 28543
rect 27120 28503 27148 28509
rect 30469 28543 30527 28549
rect 30469 28509 30481 28543
rect 30515 28540 30527 28543
rect 31018 28540 31024 28552
rect 30515 28512 31024 28540
rect 30515 28509 30527 28512
rect 30469 28503 30527 28509
rect 27120 28500 27126 28503
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 14734 28472 14740 28484
rect 13280 28444 14740 28472
rect 12897 28435 12955 28441
rect 12912 28404 12940 28435
rect 14734 28432 14740 28444
rect 14792 28432 14798 28484
rect 19613 28475 19671 28481
rect 19613 28441 19625 28475
rect 19659 28472 19671 28475
rect 20346 28472 20352 28484
rect 19659 28444 20352 28472
rect 19659 28441 19671 28444
rect 19613 28435 19671 28441
rect 20346 28432 20352 28444
rect 20404 28432 20410 28484
rect 13906 28404 13912 28416
rect 12912 28376 13912 28404
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 14829 28407 14887 28413
rect 14829 28373 14841 28407
rect 14875 28404 14887 28407
rect 15102 28404 15108 28416
rect 14875 28376 15108 28404
rect 14875 28373 14887 28376
rect 14829 28367 14887 28373
rect 15102 28364 15108 28376
rect 15160 28364 15166 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 17313 28407 17371 28413
rect 17313 28404 17325 28407
rect 15252 28376 17325 28404
rect 15252 28364 15258 28376
rect 17313 28373 17325 28376
rect 17359 28373 17371 28407
rect 17313 28367 17371 28373
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 18325 28407 18383 28413
rect 18325 28404 18337 28407
rect 18288 28376 18337 28404
rect 18288 28364 18294 28376
rect 18325 28373 18337 28376
rect 18371 28373 18383 28407
rect 20548 28404 20576 28500
rect 22005 28475 22063 28481
rect 22005 28441 22017 28475
rect 22051 28472 22063 28475
rect 23385 28475 23443 28481
rect 23385 28472 23397 28475
rect 22051 28444 23397 28472
rect 22051 28441 22063 28444
rect 22005 28435 22063 28441
rect 23385 28441 23397 28444
rect 23431 28441 23443 28475
rect 23385 28435 23443 28441
rect 25593 28475 25651 28481
rect 25593 28441 25605 28475
rect 25639 28472 25651 28475
rect 25958 28472 25964 28484
rect 25639 28444 25964 28472
rect 25639 28441 25651 28444
rect 25593 28435 25651 28441
rect 25958 28432 25964 28444
rect 26016 28432 26022 28484
rect 28074 28472 28080 28484
rect 27724 28444 28080 28472
rect 22649 28407 22707 28413
rect 22649 28404 22661 28407
rect 20548 28376 22661 28404
rect 18325 28367 18383 28373
rect 22649 28373 22661 28376
rect 22695 28373 22707 28407
rect 22649 28367 22707 28373
rect 24026 28364 24032 28416
rect 24084 28364 24090 28416
rect 25038 28364 25044 28416
rect 25096 28364 25102 28416
rect 25682 28364 25688 28416
rect 25740 28404 25746 28416
rect 26970 28404 26976 28416
rect 25740 28376 26976 28404
rect 25740 28364 25746 28376
rect 26970 28364 26976 28376
rect 27028 28364 27034 28416
rect 27062 28364 27068 28416
rect 27120 28404 27126 28416
rect 27724 28404 27752 28444
rect 28074 28432 28080 28444
rect 28132 28432 28138 28484
rect 30098 28432 30104 28484
rect 30156 28472 30162 28484
rect 31481 28475 31539 28481
rect 30156 28444 31432 28472
rect 30156 28432 30162 28444
rect 27120 28376 27752 28404
rect 27120 28364 27126 28376
rect 27890 28364 27896 28416
rect 27948 28364 27954 28416
rect 28350 28364 28356 28416
rect 28408 28364 28414 28416
rect 28626 28364 28632 28416
rect 28684 28404 28690 28416
rect 28721 28407 28779 28413
rect 28721 28404 28733 28407
rect 28684 28376 28733 28404
rect 28684 28364 28690 28376
rect 28721 28373 28733 28376
rect 28767 28373 28779 28407
rect 28721 28367 28779 28373
rect 28810 28364 28816 28416
rect 28868 28364 28874 28416
rect 30558 28364 30564 28416
rect 30616 28364 30622 28416
rect 31202 28364 31208 28416
rect 31260 28404 31266 28416
rect 31297 28407 31355 28413
rect 31297 28404 31309 28407
rect 31260 28376 31309 28404
rect 31260 28364 31266 28376
rect 31297 28373 31309 28376
rect 31343 28373 31355 28407
rect 31404 28404 31432 28444
rect 31481 28441 31493 28475
rect 31527 28472 31539 28475
rect 31570 28472 31576 28484
rect 31527 28444 31576 28472
rect 31527 28441 31539 28444
rect 31481 28435 31539 28441
rect 31570 28432 31576 28444
rect 31628 28432 31634 28484
rect 31665 28475 31723 28481
rect 31665 28441 31677 28475
rect 31711 28472 31723 28475
rect 32324 28472 32352 28580
rect 32585 28577 32597 28611
rect 32631 28577 32643 28611
rect 32585 28571 32643 28577
rect 32401 28543 32459 28549
rect 32401 28509 32413 28543
rect 32447 28540 32459 28543
rect 32876 28540 32904 28648
rect 34698 28568 34704 28620
rect 34756 28608 34762 28620
rect 34977 28611 35035 28617
rect 34977 28608 34989 28611
rect 34756 28580 34989 28608
rect 34756 28568 34762 28580
rect 34977 28577 34989 28580
rect 35023 28577 35035 28611
rect 34977 28571 35035 28577
rect 32447 28512 32904 28540
rect 32447 28509 32459 28512
rect 32401 28503 32459 28509
rect 32950 28500 32956 28552
rect 33008 28540 33014 28552
rect 33045 28543 33103 28549
rect 33045 28540 33057 28543
rect 33008 28512 33057 28540
rect 33008 28500 33014 28512
rect 33045 28509 33057 28512
rect 33091 28509 33103 28543
rect 33045 28503 33103 28509
rect 33870 28500 33876 28552
rect 33928 28500 33934 28552
rect 33962 28500 33968 28552
rect 34020 28500 34026 28552
rect 34054 28500 34060 28552
rect 34112 28540 34118 28552
rect 34149 28543 34207 28549
rect 34149 28540 34161 28543
rect 34112 28512 34161 28540
rect 34112 28500 34118 28512
rect 34149 28509 34161 28512
rect 34195 28509 34207 28543
rect 34149 28503 34207 28509
rect 34606 28500 34612 28552
rect 34664 28540 34670 28552
rect 35161 28543 35219 28549
rect 35161 28540 35173 28543
rect 34664 28512 35173 28540
rect 34664 28500 34670 28512
rect 35161 28509 35173 28512
rect 35207 28509 35219 28543
rect 35161 28503 35219 28509
rect 35802 28500 35808 28552
rect 35860 28500 35866 28552
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 36096 28549 36124 28648
rect 36265 28645 36277 28679
rect 36311 28645 36323 28679
rect 36265 28639 36323 28645
rect 36280 28608 36308 28639
rect 37826 28636 37832 28688
rect 37884 28676 37890 28688
rect 38286 28676 38292 28688
rect 37884 28648 38292 28676
rect 37884 28636 37890 28648
rect 38010 28608 38016 28620
rect 36280 28580 38016 28608
rect 38010 28568 38016 28580
rect 38068 28568 38074 28620
rect 38212 28617 38240 28648
rect 38286 28636 38292 28648
rect 38344 28636 38350 28688
rect 41046 28636 41052 28688
rect 41104 28676 41110 28688
rect 41322 28676 41328 28688
rect 41104 28648 41328 28676
rect 41104 28636 41110 28648
rect 41322 28636 41328 28648
rect 41380 28676 41386 28688
rect 41509 28679 41567 28685
rect 41509 28676 41521 28679
rect 41380 28648 41521 28676
rect 41380 28636 41386 28648
rect 41509 28645 41521 28648
rect 41555 28645 41567 28679
rect 41509 28639 41567 28645
rect 42521 28679 42579 28685
rect 42521 28645 42533 28679
rect 42567 28676 42579 28679
rect 42978 28676 42984 28688
rect 42567 28648 42984 28676
rect 42567 28645 42579 28648
rect 42521 28639 42579 28645
rect 42978 28636 42984 28648
rect 43036 28636 43042 28688
rect 38197 28611 38255 28617
rect 38197 28577 38209 28611
rect 38243 28577 38255 28611
rect 38197 28571 38255 28577
rect 41414 28568 41420 28620
rect 41472 28568 41478 28620
rect 42794 28568 42800 28620
rect 42852 28608 42858 28620
rect 43254 28608 43260 28620
rect 42852 28580 43260 28608
rect 42852 28568 42858 28580
rect 43254 28568 43260 28580
rect 43312 28568 43318 28620
rect 35989 28543 36047 28549
rect 35989 28540 36001 28543
rect 35952 28512 36001 28540
rect 35952 28500 35958 28512
rect 35989 28509 36001 28512
rect 36035 28509 36047 28543
rect 35989 28503 36047 28509
rect 36081 28543 36139 28549
rect 36081 28509 36093 28543
rect 36127 28540 36139 28543
rect 36170 28540 36176 28552
rect 36127 28512 36176 28540
rect 36127 28509 36139 28512
rect 36081 28503 36139 28509
rect 36170 28500 36176 28512
rect 36228 28500 36234 28552
rect 37001 28543 37059 28549
rect 37001 28509 37013 28543
rect 37047 28509 37059 28543
rect 37001 28503 37059 28509
rect 37185 28543 37243 28549
rect 37185 28509 37197 28543
rect 37231 28540 37243 28543
rect 38289 28543 38347 28549
rect 37231 28512 37320 28540
rect 37231 28509 37243 28512
rect 37185 28503 37243 28509
rect 33888 28472 33916 28500
rect 31711 28444 31745 28472
rect 32324 28444 33916 28472
rect 31711 28441 31723 28444
rect 31665 28435 31723 28441
rect 31680 28404 31708 28435
rect 33980 28404 34008 28500
rect 34333 28475 34391 28481
rect 34333 28441 34345 28475
rect 34379 28472 34391 28475
rect 34422 28472 34428 28484
rect 34379 28444 34428 28472
rect 34379 28441 34391 28444
rect 34333 28435 34391 28441
rect 34422 28432 34428 28444
rect 34480 28432 34486 28484
rect 34885 28475 34943 28481
rect 34885 28441 34897 28475
rect 34931 28441 34943 28475
rect 34885 28435 34943 28441
rect 31404 28376 34008 28404
rect 34900 28404 34928 28435
rect 35342 28432 35348 28484
rect 35400 28472 35406 28484
rect 37016 28472 37044 28503
rect 35400 28444 37044 28472
rect 35400 28432 35406 28444
rect 36538 28404 36544 28416
rect 34900 28376 36544 28404
rect 31297 28367 31355 28373
rect 36538 28364 36544 28376
rect 36596 28364 36602 28416
rect 36906 28364 36912 28416
rect 36964 28364 36970 28416
rect 37292 28404 37320 28512
rect 38289 28509 38301 28543
rect 38335 28540 38347 28543
rect 38470 28540 38476 28552
rect 38335 28512 38476 28540
rect 38335 28509 38347 28512
rect 38289 28503 38347 28509
rect 38470 28500 38476 28512
rect 38528 28500 38534 28552
rect 40034 28500 40040 28552
rect 40092 28540 40098 28552
rect 40218 28540 40224 28552
rect 40092 28512 40224 28540
rect 40092 28500 40098 28512
rect 40218 28500 40224 28512
rect 40276 28540 40282 28552
rect 40405 28543 40463 28549
rect 40405 28540 40417 28543
rect 40276 28512 40417 28540
rect 40276 28500 40282 28512
rect 40405 28509 40417 28512
rect 40451 28509 40463 28543
rect 40405 28503 40463 28509
rect 40589 28543 40647 28549
rect 40589 28509 40601 28543
rect 40635 28540 40647 28543
rect 40635 28512 41828 28540
rect 40635 28509 40647 28512
rect 40589 28503 40647 28509
rect 38010 28432 38016 28484
rect 38068 28472 38074 28484
rect 38194 28472 38200 28484
rect 38068 28444 38200 28472
rect 38068 28432 38074 28444
rect 38194 28432 38200 28444
rect 38252 28432 38258 28484
rect 38562 28472 38568 28484
rect 38304 28444 38568 28472
rect 38304 28404 38332 28444
rect 38562 28432 38568 28444
rect 38620 28432 38626 28484
rect 39025 28475 39083 28481
rect 39025 28441 39037 28475
rect 39071 28441 39083 28475
rect 39025 28435 39083 28441
rect 37292 28376 38332 28404
rect 38473 28407 38531 28413
rect 38473 28373 38485 28407
rect 38519 28404 38531 28407
rect 39040 28404 39068 28435
rect 39114 28432 39120 28484
rect 39172 28472 39178 28484
rect 39393 28475 39451 28481
rect 39393 28472 39405 28475
rect 39172 28444 39405 28472
rect 39172 28432 39178 28444
rect 39393 28441 39405 28444
rect 39439 28472 39451 28475
rect 39666 28472 39672 28484
rect 39439 28444 39672 28472
rect 39439 28441 39451 28444
rect 39393 28435 39451 28441
rect 39666 28432 39672 28444
rect 39724 28432 39730 28484
rect 40497 28475 40555 28481
rect 40497 28441 40509 28475
rect 40543 28472 40555 28475
rect 41690 28472 41696 28484
rect 40543 28444 41696 28472
rect 40543 28441 40555 28444
rect 40497 28435 40555 28441
rect 41690 28432 41696 28444
rect 41748 28432 41754 28484
rect 41800 28472 41828 28512
rect 41874 28500 41880 28552
rect 41932 28500 41938 28552
rect 41966 28500 41972 28552
rect 42024 28500 42030 28552
rect 42886 28500 42892 28552
rect 42944 28500 42950 28552
rect 42904 28472 42932 28500
rect 41800 28444 42932 28472
rect 38519 28376 39068 28404
rect 38519 28373 38531 28376
rect 38473 28367 38531 28373
rect 40678 28364 40684 28416
rect 40736 28404 40742 28416
rect 41141 28407 41199 28413
rect 41141 28404 41153 28407
rect 40736 28376 41153 28404
rect 40736 28364 40742 28376
rect 41141 28373 41153 28376
rect 41187 28373 41199 28407
rect 41141 28367 41199 28373
rect 1104 28314 43884 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 43884 28314
rect 1104 28240 43884 28262
rect 14734 28160 14740 28212
rect 14792 28200 14798 28212
rect 14829 28203 14887 28209
rect 14829 28200 14841 28203
rect 14792 28172 14841 28200
rect 14792 28160 14798 28172
rect 14829 28169 14841 28172
rect 14875 28169 14887 28203
rect 14829 28163 14887 28169
rect 16942 28160 16948 28212
rect 17000 28160 17006 28212
rect 18601 28203 18659 28209
rect 18601 28169 18613 28203
rect 18647 28200 18659 28203
rect 21450 28200 21456 28212
rect 18647 28172 21456 28200
rect 18647 28169 18659 28172
rect 18601 28163 18659 28169
rect 21450 28160 21456 28172
rect 21508 28160 21514 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22281 28203 22339 28209
rect 22281 28200 22293 28203
rect 22152 28172 22293 28200
rect 22152 28160 22158 28172
rect 22281 28169 22293 28172
rect 22327 28169 22339 28203
rect 22281 28163 22339 28169
rect 23014 28160 23020 28212
rect 23072 28200 23078 28212
rect 23385 28203 23443 28209
rect 23385 28200 23397 28203
rect 23072 28172 23397 28200
rect 23072 28160 23078 28172
rect 23385 28169 23397 28172
rect 23431 28169 23443 28203
rect 23385 28163 23443 28169
rect 25593 28203 25651 28209
rect 25593 28169 25605 28203
rect 25639 28200 25651 28203
rect 25682 28200 25688 28212
rect 25639 28172 25688 28200
rect 25639 28169 25651 28172
rect 25593 28163 25651 28169
rect 25682 28160 25688 28172
rect 25740 28160 25746 28212
rect 26418 28160 26424 28212
rect 26476 28200 26482 28212
rect 27157 28203 27215 28209
rect 27157 28200 27169 28203
rect 26476 28172 27169 28200
rect 26476 28160 26482 28172
rect 27157 28169 27169 28172
rect 27203 28169 27215 28203
rect 27157 28163 27215 28169
rect 27617 28203 27675 28209
rect 27617 28169 27629 28203
rect 27663 28200 27675 28203
rect 28350 28200 28356 28212
rect 27663 28172 28356 28200
rect 27663 28169 27675 28172
rect 27617 28163 27675 28169
rect 28350 28160 28356 28172
rect 28408 28160 28414 28212
rect 28905 28203 28963 28209
rect 28905 28169 28917 28203
rect 28951 28200 28963 28203
rect 30834 28200 30840 28212
rect 28951 28172 30840 28200
rect 28951 28169 28963 28172
rect 28905 28163 28963 28169
rect 30834 28160 30840 28172
rect 30892 28160 30898 28212
rect 32677 28203 32735 28209
rect 32677 28169 32689 28203
rect 32723 28200 32735 28203
rect 32766 28200 32772 28212
rect 32723 28172 32772 28200
rect 32723 28169 32735 28172
rect 32677 28163 32735 28169
rect 32766 28160 32772 28172
rect 32824 28160 32830 28212
rect 32950 28160 32956 28212
rect 33008 28160 33014 28212
rect 33226 28160 33232 28212
rect 33284 28200 33290 28212
rect 33413 28203 33471 28209
rect 33413 28200 33425 28203
rect 33284 28172 33425 28200
rect 33284 28160 33290 28172
rect 33413 28169 33425 28172
rect 33459 28169 33471 28203
rect 33413 28163 33471 28169
rect 34422 28160 34428 28212
rect 34480 28200 34486 28212
rect 35434 28200 35440 28212
rect 34480 28172 35440 28200
rect 34480 28160 34486 28172
rect 35434 28160 35440 28172
rect 35492 28160 35498 28212
rect 35894 28160 35900 28212
rect 35952 28160 35958 28212
rect 36354 28160 36360 28212
rect 36412 28160 36418 28212
rect 40862 28160 40868 28212
rect 40920 28200 40926 28212
rect 41325 28203 41383 28209
rect 41325 28200 41337 28203
rect 40920 28172 41337 28200
rect 40920 28160 40926 28172
rect 41325 28169 41337 28172
rect 41371 28169 41383 28203
rect 41325 28163 41383 28169
rect 41782 28160 41788 28212
rect 41840 28200 41846 28212
rect 41969 28203 42027 28209
rect 41969 28200 41981 28203
rect 41840 28172 41981 28200
rect 41840 28160 41846 28172
rect 41969 28169 41981 28172
rect 42015 28169 42027 28203
rect 41969 28163 42027 28169
rect 18046 28132 18052 28144
rect 17604 28104 18052 28132
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28064 12863 28067
rect 13170 28064 13176 28076
rect 12851 28036 13176 28064
rect 12851 28033 12863 28036
rect 12805 28027 12863 28033
rect 13170 28024 13176 28036
rect 13228 28024 13234 28076
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 17310 28024 17316 28076
rect 17368 28064 17374 28076
rect 17604 28073 17632 28104
rect 18046 28092 18052 28104
rect 18104 28132 18110 28144
rect 18104 28104 18368 28132
rect 18104 28092 18110 28104
rect 17405 28067 17463 28073
rect 17405 28064 17417 28067
rect 17368 28036 17417 28064
rect 17368 28024 17374 28036
rect 17405 28033 17417 28036
rect 17451 28033 17463 28067
rect 17405 28027 17463 28033
rect 17589 28067 17647 28073
rect 17589 28033 17601 28067
rect 17635 28033 17647 28067
rect 17589 28027 17647 28033
rect 18230 28024 18236 28076
rect 18288 28024 18294 28076
rect 18340 28064 18368 28104
rect 20898 28092 20904 28144
rect 20956 28092 20962 28144
rect 21358 28092 21364 28144
rect 21416 28092 21422 28144
rect 24026 28092 24032 28144
rect 24084 28132 24090 28144
rect 26786 28132 26792 28144
rect 24084 28104 26792 28132
rect 24084 28092 24090 28104
rect 23569 28067 23627 28073
rect 18340 28036 23520 28064
rect 12897 27999 12955 28005
rect 12897 27965 12909 27999
rect 12943 27996 12955 27999
rect 12986 27996 12992 28008
rect 12943 27968 12992 27996
rect 12943 27965 12955 27968
rect 12897 27959 12955 27965
rect 12986 27956 12992 27968
rect 13044 27956 13050 28008
rect 15102 27956 15108 28008
rect 15160 27956 15166 28008
rect 17497 27999 17555 28005
rect 17497 27965 17509 27999
rect 17543 27996 17555 27999
rect 18141 27999 18199 28005
rect 18141 27996 18153 27999
rect 17543 27968 18153 27996
rect 17543 27965 17555 27968
rect 17497 27959 17555 27965
rect 18141 27965 18153 27968
rect 18187 27965 18199 27999
rect 18141 27959 18199 27965
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27996 20499 27999
rect 20622 27996 20628 28008
rect 20487 27968 20628 27996
rect 20487 27965 20499 27968
rect 20441 27959 20499 27965
rect 20622 27956 20628 27968
rect 20680 27956 20686 28008
rect 19978 27888 19984 27940
rect 20036 27928 20042 27940
rect 20533 27931 20591 27937
rect 20533 27928 20545 27931
rect 20036 27900 20545 27928
rect 20036 27888 20042 27900
rect 20533 27897 20545 27900
rect 20579 27897 20591 27931
rect 20533 27891 20591 27897
rect 13173 27863 13231 27869
rect 13173 27829 13185 27863
rect 13219 27860 13231 27863
rect 13906 27860 13912 27872
rect 13219 27832 13912 27860
rect 13219 27829 13231 27832
rect 13173 27823 13231 27829
rect 13906 27820 13912 27832
rect 13964 27860 13970 27872
rect 14550 27860 14556 27872
rect 13964 27832 14556 27860
rect 13964 27820 13970 27832
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 22922 27820 22928 27872
rect 22980 27820 22986 27872
rect 23492 27860 23520 28036
rect 23569 28033 23581 28067
rect 23615 28064 23627 28067
rect 23934 28064 23940 28076
rect 23615 28036 23940 28064
rect 23615 28033 23627 28036
rect 23569 28027 23627 28033
rect 23934 28024 23940 28036
rect 23992 28024 23998 28076
rect 24228 28073 24256 28104
rect 26786 28092 26792 28104
rect 26844 28092 26850 28144
rect 27525 28135 27583 28141
rect 27525 28101 27537 28135
rect 27571 28132 27583 28135
rect 28258 28132 28264 28144
rect 27571 28104 28264 28132
rect 27571 28101 27583 28104
rect 27525 28095 27583 28101
rect 28258 28092 28264 28104
rect 28316 28092 28322 28144
rect 32490 28132 32496 28144
rect 30576 28104 32496 28132
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 24480 28067 24538 28073
rect 24480 28033 24492 28067
rect 24526 28064 24538 28067
rect 25498 28064 25504 28076
rect 24526 28036 25504 28064
rect 24526 28033 24538 28036
rect 24480 28027 24538 28033
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 28537 28067 28595 28073
rect 28537 28033 28549 28067
rect 28583 28064 28595 28067
rect 28718 28064 28724 28076
rect 28583 28036 28724 28064
rect 28583 28033 28595 28036
rect 28537 28027 28595 28033
rect 28718 28024 28724 28036
rect 28776 28024 28782 28076
rect 29362 28024 29368 28076
rect 29420 28024 29426 28076
rect 29546 28024 29552 28076
rect 29604 28024 29610 28076
rect 30576 28073 30604 28104
rect 32490 28092 32496 28104
rect 32548 28092 32554 28144
rect 32585 28135 32643 28141
rect 32585 28101 32597 28135
rect 32631 28132 32643 28135
rect 37090 28132 37096 28144
rect 32631 28104 37096 28132
rect 32631 28101 32643 28104
rect 32585 28095 32643 28101
rect 37090 28092 37096 28104
rect 37148 28092 37154 28144
rect 38102 28092 38108 28144
rect 38160 28092 38166 28144
rect 42794 28132 42800 28144
rect 40052 28104 42800 28132
rect 30561 28067 30619 28073
rect 30561 28033 30573 28067
rect 30607 28033 30619 28067
rect 30561 28027 30619 28033
rect 30745 28067 30803 28073
rect 30745 28033 30757 28067
rect 30791 28033 30803 28067
rect 30745 28027 30803 28033
rect 23750 27956 23756 28008
rect 23808 27956 23814 28008
rect 27338 27956 27344 28008
rect 27396 27996 27402 28008
rect 27709 27999 27767 28005
rect 27709 27996 27721 27999
rect 27396 27968 27721 27996
rect 27396 27956 27402 27968
rect 27709 27965 27721 27968
rect 27755 27965 27767 27999
rect 27709 27959 27767 27965
rect 27890 27956 27896 28008
rect 27948 27996 27954 28008
rect 28445 27999 28503 28005
rect 28445 27996 28457 27999
rect 27948 27968 28457 27996
rect 27948 27956 27954 27968
rect 28445 27965 28457 27968
rect 28491 27965 28503 27999
rect 30760 27996 30788 28027
rect 31202 28024 31208 28076
rect 31260 28024 31266 28076
rect 31386 28024 31392 28076
rect 31444 28064 31450 28076
rect 32309 28067 32367 28073
rect 32309 28064 32321 28067
rect 31444 28036 32321 28064
rect 31444 28024 31450 28036
rect 32309 28033 32321 28036
rect 32355 28033 32367 28067
rect 32309 28027 32367 28033
rect 34149 28067 34207 28073
rect 34149 28033 34161 28067
rect 34195 28064 34207 28067
rect 34195 28036 34284 28064
rect 34195 28033 34207 28036
rect 34149 28027 34207 28033
rect 34256 28008 34284 28036
rect 34514 28024 34520 28076
rect 34572 28024 34578 28076
rect 34701 28067 34759 28073
rect 34701 28033 34713 28067
rect 34747 28064 34759 28067
rect 34747 28036 35112 28064
rect 34747 28033 34759 28036
rect 34701 28027 34759 28033
rect 32582 27996 32588 28008
rect 30760 27968 32588 27996
rect 28445 27959 28503 27965
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 32766 27956 32772 28008
rect 32824 28005 32830 28008
rect 32824 27999 32852 28005
rect 32840 27965 32852 27999
rect 32824 27959 32852 27965
rect 32824 27956 32830 27959
rect 34238 27956 34244 28008
rect 34296 27956 34302 28008
rect 34330 27956 34336 28008
rect 34388 27956 34394 28008
rect 34422 27956 34428 28008
rect 34480 27956 34486 28008
rect 35084 27996 35112 28036
rect 35158 28024 35164 28076
rect 35216 28064 35222 28076
rect 35529 28067 35587 28073
rect 35529 28064 35541 28067
rect 35216 28036 35541 28064
rect 35216 28024 35222 28036
rect 35529 28033 35541 28036
rect 35575 28033 35587 28067
rect 35529 28027 35587 28033
rect 35713 28067 35771 28073
rect 35713 28033 35725 28067
rect 35759 28064 35771 28067
rect 36446 28064 36452 28076
rect 35759 28036 36452 28064
rect 35759 28033 35771 28036
rect 35713 28027 35771 28033
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 38010 28064 38016 28076
rect 38068 28073 38074 28076
rect 37976 28036 38016 28064
rect 38010 28024 38016 28036
rect 38068 28027 38076 28073
rect 38120 28064 38148 28092
rect 40052 28076 40080 28104
rect 42794 28092 42800 28104
rect 42852 28092 42858 28144
rect 38197 28067 38255 28073
rect 38197 28064 38209 28067
rect 38120 28036 38209 28064
rect 38197 28033 38209 28036
rect 38243 28033 38255 28067
rect 38197 28027 38255 28033
rect 39025 28067 39083 28073
rect 39025 28033 39037 28067
rect 39071 28064 39083 28067
rect 40034 28064 40040 28076
rect 39071 28036 40040 28064
rect 39071 28033 39083 28036
rect 39025 28027 39083 28033
rect 38068 28024 38074 28027
rect 40034 28024 40040 28036
rect 40092 28024 40098 28076
rect 40129 28067 40187 28073
rect 40129 28033 40141 28067
rect 40175 28064 40187 28067
rect 40586 28064 40592 28076
rect 40175 28036 40592 28064
rect 40175 28033 40187 28036
rect 40129 28027 40187 28033
rect 40586 28024 40592 28036
rect 40644 28064 40650 28076
rect 41230 28064 41236 28076
rect 40644 28036 41236 28064
rect 40644 28024 40650 28036
rect 41230 28024 41236 28036
rect 41288 28024 41294 28076
rect 43257 28067 43315 28073
rect 43257 28033 43269 28067
rect 43303 28064 43315 28067
rect 43438 28064 43444 28076
rect 43303 28036 43444 28064
rect 43303 28033 43315 28036
rect 43257 28027 43315 28033
rect 43438 28024 43444 28036
rect 43496 28064 43502 28076
rect 43990 28064 43996 28076
rect 43496 28036 43996 28064
rect 43496 28024 43502 28036
rect 43990 28024 43996 28036
rect 44048 28024 44054 28076
rect 35986 27996 35992 28008
rect 35084 27968 35992 27996
rect 35986 27956 35992 27968
rect 36044 27956 36050 28008
rect 36998 27956 37004 28008
rect 37056 27996 37062 28008
rect 39209 27999 39267 28005
rect 39209 27996 39221 27999
rect 37056 27968 39221 27996
rect 37056 27956 37062 27968
rect 39209 27965 39221 27968
rect 39255 27996 39267 27999
rect 39850 27996 39856 28008
rect 39255 27968 39856 27996
rect 39255 27965 39267 27968
rect 39209 27959 39267 27965
rect 39850 27956 39856 27968
rect 39908 27956 39914 28008
rect 40402 27956 40408 28008
rect 40460 27996 40466 28008
rect 40957 27999 41015 28005
rect 40957 27996 40969 27999
rect 40460 27968 40969 27996
rect 40460 27956 40466 27968
rect 40957 27965 40969 27968
rect 41003 27965 41015 27999
rect 40957 27959 41015 27965
rect 41046 27956 41052 28008
rect 41104 27956 41110 28008
rect 41509 27999 41567 28005
rect 41509 27965 41521 27999
rect 41555 27996 41567 27999
rect 41966 27996 41972 28008
rect 41555 27968 41972 27996
rect 41555 27965 41567 27968
rect 41509 27959 41567 27965
rect 29457 27931 29515 27937
rect 29457 27928 29469 27931
rect 25148 27900 29469 27928
rect 25148 27860 25176 27900
rect 29457 27897 29469 27900
rect 29503 27897 29515 27931
rect 29457 27891 29515 27897
rect 29914 27888 29920 27940
rect 29972 27928 29978 27940
rect 30745 27931 30803 27937
rect 29972 27900 30696 27928
rect 29972 27888 29978 27900
rect 23492 27832 25176 27860
rect 25866 27820 25872 27872
rect 25924 27860 25930 27872
rect 26053 27863 26111 27869
rect 26053 27860 26065 27863
rect 25924 27832 26065 27860
rect 25924 27820 25930 27832
rect 26053 27829 26065 27832
rect 26099 27829 26111 27863
rect 26053 27823 26111 27829
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 29638 27860 29644 27872
rect 29052 27832 29644 27860
rect 29052 27820 29058 27832
rect 29638 27820 29644 27832
rect 29696 27860 29702 27872
rect 30009 27863 30067 27869
rect 30009 27860 30021 27863
rect 29696 27832 30021 27860
rect 29696 27820 29702 27832
rect 30009 27829 30021 27832
rect 30055 27860 30067 27863
rect 30282 27860 30288 27872
rect 30055 27832 30288 27860
rect 30055 27829 30067 27832
rect 30009 27823 30067 27829
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 30668 27860 30696 27900
rect 30745 27897 30757 27931
rect 30791 27928 30803 27931
rect 32122 27928 32128 27940
rect 30791 27900 32128 27928
rect 30791 27897 30803 27900
rect 30745 27891 30803 27897
rect 32122 27888 32128 27900
rect 32180 27888 32186 27940
rect 32306 27888 32312 27940
rect 32364 27928 32370 27940
rect 33965 27931 34023 27937
rect 33965 27928 33977 27931
rect 32364 27900 33977 27928
rect 32364 27888 32370 27900
rect 33965 27897 33977 27900
rect 34011 27897 34023 27931
rect 33965 27891 34023 27897
rect 37458 27888 37464 27940
rect 37516 27888 37522 27940
rect 38562 27888 38568 27940
rect 38620 27928 38626 27940
rect 38620 27900 38976 27928
rect 38620 27888 38626 27900
rect 31386 27860 31392 27872
rect 30668 27832 31392 27860
rect 31386 27820 31392 27832
rect 31444 27820 31450 27872
rect 33778 27820 33784 27872
rect 33836 27860 33842 27872
rect 35529 27863 35587 27869
rect 35529 27860 35541 27863
rect 33836 27832 35541 27860
rect 33836 27820 33842 27832
rect 35529 27829 35541 27832
rect 35575 27860 35587 27863
rect 36906 27860 36912 27872
rect 35575 27832 36912 27860
rect 35575 27829 35587 27832
rect 35529 27823 35587 27829
rect 36906 27820 36912 27832
rect 36964 27820 36970 27872
rect 37826 27820 37832 27872
rect 37884 27860 37890 27872
rect 38013 27863 38071 27869
rect 38013 27860 38025 27863
rect 37884 27832 38025 27860
rect 37884 27820 37890 27832
rect 38013 27829 38025 27832
rect 38059 27829 38071 27863
rect 38013 27823 38071 27829
rect 38194 27820 38200 27872
rect 38252 27860 38258 27872
rect 38381 27863 38439 27869
rect 38381 27860 38393 27863
rect 38252 27832 38393 27860
rect 38252 27820 38258 27832
rect 38381 27829 38393 27832
rect 38427 27829 38439 27863
rect 38381 27823 38439 27829
rect 38654 27820 38660 27872
rect 38712 27860 38718 27872
rect 38841 27863 38899 27869
rect 38841 27860 38853 27863
rect 38712 27832 38853 27860
rect 38712 27820 38718 27832
rect 38841 27829 38853 27832
rect 38887 27829 38899 27863
rect 38948 27860 38976 27900
rect 39942 27888 39948 27940
rect 40000 27928 40006 27940
rect 41524 27928 41552 27959
rect 41966 27956 41972 27968
rect 42024 27956 42030 28008
rect 40000 27900 41552 27928
rect 40000 27888 40006 27900
rect 39206 27860 39212 27872
rect 38948 27832 39212 27860
rect 38841 27823 38899 27829
rect 39206 27820 39212 27832
rect 39264 27820 39270 27872
rect 39390 27820 39396 27872
rect 39448 27860 39454 27872
rect 40037 27863 40095 27869
rect 40037 27860 40049 27863
rect 39448 27832 40049 27860
rect 39448 27820 39454 27832
rect 40037 27829 40049 27832
rect 40083 27829 40095 27863
rect 40037 27823 40095 27829
rect 43070 27820 43076 27872
rect 43128 27860 43134 27872
rect 43165 27863 43223 27869
rect 43165 27860 43177 27863
rect 43128 27832 43177 27860
rect 43128 27820 43134 27832
rect 43165 27829 43177 27832
rect 43211 27860 43223 27863
rect 43530 27860 43536 27872
rect 43211 27832 43536 27860
rect 43211 27829 43223 27832
rect 43165 27823 43223 27829
rect 43530 27820 43536 27832
rect 43588 27820 43594 27872
rect 1104 27770 43884 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 43884 27770
rect 1104 27696 43884 27718
rect 26050 27656 26056 27668
rect 23768 27628 26056 27656
rect 20254 27548 20260 27600
rect 20312 27588 20318 27600
rect 20438 27588 20444 27600
rect 20312 27560 20444 27588
rect 20312 27548 20318 27560
rect 20438 27548 20444 27560
rect 20496 27548 20502 27600
rect 23658 27548 23664 27600
rect 23716 27588 23722 27600
rect 23768 27588 23796 27628
rect 26050 27616 26056 27628
rect 26108 27656 26114 27668
rect 26237 27659 26295 27665
rect 26237 27656 26249 27659
rect 26108 27628 26249 27656
rect 26108 27616 26114 27628
rect 26237 27625 26249 27628
rect 26283 27625 26295 27659
rect 26237 27619 26295 27625
rect 27338 27616 27344 27668
rect 27396 27616 27402 27668
rect 27982 27656 27988 27668
rect 27448 27628 27988 27656
rect 23716 27560 23796 27588
rect 23716 27548 23722 27560
rect 23842 27548 23848 27600
rect 23900 27548 23906 27600
rect 25498 27548 25504 27600
rect 25556 27548 25562 27600
rect 26694 27588 26700 27600
rect 26436 27560 26700 27588
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14277 27523 14335 27529
rect 14277 27520 14289 27523
rect 13872 27492 14289 27520
rect 13872 27480 13878 27492
rect 14277 27489 14289 27492
rect 14323 27520 14335 27523
rect 21361 27523 21419 27529
rect 21361 27520 21373 27523
rect 14323 27492 21373 27520
rect 14323 27489 14335 27492
rect 14277 27483 14335 27489
rect 21361 27489 21373 27492
rect 21407 27489 21419 27523
rect 24394 27520 24400 27532
rect 21361 27483 21419 27489
rect 23860 27492 24400 27520
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 18966 27412 18972 27464
rect 19024 27452 19030 27464
rect 19024 27424 19564 27452
rect 19024 27412 19030 27424
rect 15933 27387 15991 27393
rect 15933 27353 15945 27387
rect 15979 27384 15991 27387
rect 19426 27384 19432 27396
rect 15979 27356 19432 27384
rect 15979 27353 15991 27356
rect 15933 27347 15991 27353
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 19536 27384 19564 27424
rect 21450 27412 21456 27464
rect 21508 27452 21514 27464
rect 21617 27455 21675 27461
rect 21617 27452 21629 27455
rect 21508 27424 21629 27452
rect 21508 27412 21514 27424
rect 21617 27421 21629 27424
rect 21663 27421 21675 27455
rect 21617 27415 21675 27421
rect 23750 27412 23756 27464
rect 23808 27452 23814 27464
rect 23860 27452 23888 27492
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 25038 27480 25044 27532
rect 25096 27520 25102 27532
rect 26436 27529 26464 27560
rect 26694 27548 26700 27560
rect 26752 27588 26758 27600
rect 27448 27588 27476 27628
rect 27982 27616 27988 27628
rect 28040 27616 28046 27668
rect 29089 27659 29147 27665
rect 29089 27625 29101 27659
rect 29135 27656 29147 27659
rect 29362 27656 29368 27668
rect 29135 27628 29368 27656
rect 29135 27625 29147 27628
rect 29089 27619 29147 27625
rect 29362 27616 29368 27628
rect 29420 27616 29426 27668
rect 29546 27616 29552 27668
rect 29604 27656 29610 27668
rect 29733 27659 29791 27665
rect 29733 27656 29745 27659
rect 29604 27628 29745 27656
rect 29604 27616 29610 27628
rect 29733 27625 29745 27628
rect 29779 27625 29791 27659
rect 32766 27656 32772 27668
rect 29733 27619 29791 27625
rect 31588 27628 32772 27656
rect 26752 27560 27476 27588
rect 27709 27591 27767 27597
rect 26752 27548 26758 27560
rect 27709 27557 27721 27591
rect 27755 27588 27767 27591
rect 27798 27588 27804 27600
rect 27755 27560 27804 27588
rect 27755 27557 27767 27560
rect 27709 27551 27767 27557
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 31588 27597 31616 27628
rect 32766 27616 32772 27628
rect 32824 27616 32830 27668
rect 34422 27616 34428 27668
rect 34480 27656 34486 27668
rect 34974 27656 34980 27668
rect 34480 27628 34980 27656
rect 34480 27616 34486 27628
rect 34974 27616 34980 27628
rect 35032 27656 35038 27668
rect 35342 27656 35348 27668
rect 35032 27628 35348 27656
rect 35032 27616 35038 27628
rect 35342 27616 35348 27628
rect 35400 27616 35406 27668
rect 35526 27616 35532 27668
rect 35584 27656 35590 27668
rect 35805 27659 35863 27665
rect 35805 27656 35817 27659
rect 35584 27628 35817 27656
rect 35584 27616 35590 27628
rect 35805 27625 35817 27628
rect 35851 27625 35863 27659
rect 35805 27619 35863 27625
rect 36354 27616 36360 27668
rect 36412 27656 36418 27668
rect 36630 27656 36636 27668
rect 36412 27628 36636 27656
rect 36412 27616 36418 27628
rect 36630 27616 36636 27628
rect 36688 27616 36694 27668
rect 38102 27616 38108 27668
rect 38160 27656 38166 27668
rect 38838 27656 38844 27668
rect 38160 27628 38844 27656
rect 38160 27616 38166 27628
rect 38838 27616 38844 27628
rect 38896 27656 38902 27668
rect 39393 27659 39451 27665
rect 39393 27656 39405 27659
rect 38896 27628 39405 27656
rect 38896 27616 38902 27628
rect 39393 27625 39405 27628
rect 39439 27656 39451 27659
rect 40402 27656 40408 27668
rect 39439 27628 40408 27656
rect 39439 27625 39451 27628
rect 39393 27619 39451 27625
rect 40402 27616 40408 27628
rect 40460 27616 40466 27668
rect 40494 27616 40500 27668
rect 40552 27656 40558 27668
rect 40552 27628 41184 27656
rect 40552 27616 40558 27628
rect 41156 27600 41184 27628
rect 41414 27616 41420 27668
rect 41472 27616 41478 27668
rect 42337 27659 42395 27665
rect 42337 27656 42349 27659
rect 41524 27628 42349 27656
rect 31297 27591 31355 27597
rect 31297 27557 31309 27591
rect 31343 27588 31355 27591
rect 31573 27591 31631 27597
rect 31343 27560 31524 27588
rect 31343 27557 31355 27560
rect 31297 27551 31355 27557
rect 26421 27523 26479 27529
rect 26421 27520 26433 27523
rect 25096 27492 26433 27520
rect 25096 27480 25102 27492
rect 26421 27489 26433 27492
rect 26467 27489 26479 27523
rect 30469 27523 30527 27529
rect 30469 27520 30481 27523
rect 26421 27483 26479 27489
rect 26528 27492 30481 27520
rect 23808 27424 23888 27452
rect 23808 27412 23814 27424
rect 23934 27412 23940 27464
rect 23992 27452 23998 27464
rect 24762 27452 24768 27464
rect 23992 27424 24768 27452
rect 23992 27412 23998 27424
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 25682 27412 25688 27464
rect 25740 27412 25746 27464
rect 26528 27461 26556 27492
rect 30469 27489 30481 27492
rect 30515 27489 30527 27523
rect 30469 27483 30527 27489
rect 31386 27480 31392 27532
rect 31444 27480 31450 27532
rect 31496 27520 31524 27560
rect 31573 27557 31585 27591
rect 31619 27557 31631 27591
rect 31573 27551 31631 27557
rect 31662 27548 31668 27600
rect 31720 27588 31726 27600
rect 32033 27591 32091 27597
rect 32033 27588 32045 27591
rect 31720 27560 32045 27588
rect 31720 27548 31726 27560
rect 32033 27557 32045 27560
rect 32079 27557 32091 27591
rect 32033 27551 32091 27557
rect 32674 27548 32680 27600
rect 32732 27588 32738 27600
rect 34333 27591 34391 27597
rect 34333 27588 34345 27591
rect 32732 27560 34345 27588
rect 32732 27548 32738 27560
rect 34333 27557 34345 27560
rect 34379 27588 34391 27591
rect 34606 27588 34612 27600
rect 34379 27560 34612 27588
rect 34379 27557 34391 27560
rect 34333 27551 34391 27557
rect 34606 27548 34612 27560
rect 34664 27548 34670 27600
rect 35084 27560 36768 27588
rect 31938 27520 31944 27532
rect 31496 27492 31944 27520
rect 31938 27480 31944 27492
rect 31996 27480 32002 27532
rect 33134 27520 33140 27532
rect 32232 27492 33140 27520
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 25792 27424 26525 27452
rect 24581 27387 24639 27393
rect 24581 27384 24593 27387
rect 19536 27356 24593 27384
rect 24581 27353 24593 27356
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 24946 27344 24952 27396
rect 25004 27344 25010 27396
rect 20622 27276 20628 27328
rect 20680 27316 20686 27328
rect 20717 27319 20775 27325
rect 20717 27316 20729 27319
rect 20680 27288 20729 27316
rect 20680 27276 20686 27288
rect 20717 27285 20729 27288
rect 20763 27285 20775 27319
rect 20717 27279 20775 27285
rect 22646 27276 22652 27328
rect 22704 27316 22710 27328
rect 22741 27319 22799 27325
rect 22741 27316 22753 27319
rect 22704 27288 22753 27316
rect 22704 27276 22710 27288
rect 22741 27285 22753 27288
rect 22787 27285 22799 27319
rect 22741 27279 22799 27285
rect 22830 27276 22836 27328
rect 22888 27316 22894 27328
rect 24486 27316 24492 27328
rect 22888 27288 24492 27316
rect 22888 27276 22894 27288
rect 24486 27276 24492 27288
rect 24544 27316 24550 27328
rect 25792 27316 25820 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 27522 27412 27528 27464
rect 27580 27412 27586 27464
rect 27614 27412 27620 27464
rect 27672 27452 27678 27464
rect 27801 27455 27859 27461
rect 27801 27452 27813 27455
rect 27672 27424 27813 27452
rect 27672 27412 27678 27424
rect 27801 27421 27813 27424
rect 27847 27452 27859 27455
rect 27890 27452 27896 27464
rect 27847 27424 27896 27452
rect 27847 27421 27859 27424
rect 27801 27415 27859 27421
rect 27890 27412 27896 27424
rect 27948 27412 27954 27464
rect 28074 27412 28080 27464
rect 28132 27452 28138 27464
rect 28997 27455 29055 27461
rect 28997 27452 29009 27455
rect 28132 27424 29009 27452
rect 28132 27412 28138 27424
rect 28997 27421 29009 27424
rect 29043 27421 29055 27455
rect 28997 27415 29055 27421
rect 29178 27412 29184 27464
rect 29236 27412 29242 27464
rect 30009 27455 30067 27461
rect 30009 27421 30021 27455
rect 30055 27452 30067 27455
rect 30282 27452 30288 27464
rect 30055 27424 30288 27452
rect 30055 27421 30067 27424
rect 30009 27415 30067 27421
rect 30282 27412 30288 27424
rect 30340 27412 30346 27464
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27452 31263 27455
rect 32232 27452 32260 27492
rect 33134 27480 33140 27492
rect 33192 27520 33198 27532
rect 33597 27523 33655 27529
rect 33597 27520 33609 27523
rect 33192 27492 33609 27520
rect 33192 27480 33198 27492
rect 33597 27489 33609 27492
rect 33643 27489 33655 27523
rect 33597 27483 33655 27489
rect 34238 27480 34244 27532
rect 34296 27520 34302 27532
rect 35084 27520 35112 27560
rect 34296 27492 35112 27520
rect 34296 27480 34302 27492
rect 31251 27424 32260 27452
rect 31251 27421 31263 27424
rect 31205 27415 31263 27421
rect 32306 27412 32312 27464
rect 32364 27412 32370 27464
rect 32401 27455 32459 27461
rect 32401 27421 32413 27455
rect 32447 27452 32459 27455
rect 32766 27452 32772 27464
rect 32447 27424 32772 27452
rect 32447 27421 32459 27424
rect 32401 27415 32459 27421
rect 32766 27412 32772 27424
rect 32824 27412 32830 27464
rect 33410 27412 33416 27464
rect 33468 27412 33474 27464
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27452 33563 27455
rect 33551 27424 33640 27452
rect 33551 27421 33563 27424
rect 33505 27415 33563 27421
rect 33612 27396 33640 27424
rect 34054 27412 34060 27464
rect 34112 27452 34118 27464
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 34112 27424 34161 27452
rect 34112 27412 34118 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34330 27412 34336 27464
rect 34388 27412 34394 27464
rect 34992 27461 35020 27492
rect 35710 27480 35716 27532
rect 35768 27520 35774 27532
rect 35768 27492 35940 27520
rect 35768 27480 35774 27492
rect 34977 27455 35035 27461
rect 34977 27421 34989 27455
rect 35023 27421 35035 27455
rect 34977 27415 35035 27421
rect 35066 27412 35072 27464
rect 35124 27452 35130 27464
rect 35161 27455 35219 27461
rect 35161 27452 35173 27455
rect 35124 27424 35173 27452
rect 35124 27412 35130 27424
rect 35161 27421 35173 27424
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 35618 27412 35624 27464
rect 35676 27461 35682 27464
rect 35676 27452 35685 27461
rect 35805 27455 35863 27461
rect 35676 27424 35721 27452
rect 35676 27415 35685 27424
rect 35805 27421 35817 27455
rect 35851 27421 35863 27455
rect 35912 27452 35940 27492
rect 36354 27480 36360 27532
rect 36412 27480 36418 27532
rect 36538 27452 36544 27464
rect 35912 27424 36544 27452
rect 35805 27415 35863 27421
rect 35676 27412 35682 27415
rect 26050 27344 26056 27396
rect 26108 27384 26114 27396
rect 26237 27387 26295 27393
rect 26237 27384 26249 27387
rect 26108 27356 26249 27384
rect 26108 27344 26114 27356
rect 26237 27353 26249 27356
rect 26283 27384 26295 27387
rect 28810 27384 28816 27396
rect 26283 27356 28816 27384
rect 26283 27353 26295 27356
rect 26237 27347 26295 27353
rect 28810 27344 28816 27356
rect 28868 27344 28874 27396
rect 29733 27387 29791 27393
rect 29733 27353 29745 27387
rect 29779 27384 29791 27387
rect 30190 27384 30196 27396
rect 29779 27356 30196 27384
rect 29779 27353 29791 27356
rect 29733 27347 29791 27353
rect 30190 27344 30196 27356
rect 30248 27344 30254 27396
rect 31573 27387 31631 27393
rect 31573 27353 31585 27387
rect 31619 27384 31631 27387
rect 32030 27384 32036 27396
rect 31619 27356 32036 27384
rect 31619 27353 31631 27356
rect 31573 27347 31631 27353
rect 32030 27344 32036 27356
rect 32088 27344 32094 27396
rect 32122 27344 32128 27396
rect 32180 27384 32186 27396
rect 32585 27387 32643 27393
rect 32585 27384 32597 27387
rect 32180 27356 32597 27384
rect 32180 27344 32186 27356
rect 32585 27353 32597 27356
rect 32631 27353 32643 27387
rect 32585 27347 32643 27353
rect 33594 27344 33600 27396
rect 33652 27384 33658 27396
rect 33652 27356 34284 27384
rect 33652 27344 33658 27356
rect 24544 27288 25820 27316
rect 26697 27319 26755 27325
rect 24544 27276 24550 27288
rect 26697 27285 26709 27319
rect 26743 27316 26755 27319
rect 27246 27316 27252 27328
rect 26743 27288 27252 27316
rect 26743 27285 26755 27288
rect 26697 27279 26755 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 27338 27276 27344 27328
rect 27396 27316 27402 27328
rect 28261 27319 28319 27325
rect 28261 27316 28273 27319
rect 27396 27288 28273 27316
rect 27396 27276 27402 27288
rect 28261 27285 28273 27288
rect 28307 27316 28319 27319
rect 28626 27316 28632 27328
rect 28307 27288 28632 27316
rect 28307 27285 28319 27288
rect 28261 27279 28319 27285
rect 28626 27276 28632 27288
rect 28684 27276 28690 27328
rect 29917 27319 29975 27325
rect 29917 27285 29929 27319
rect 29963 27316 29975 27319
rect 30374 27316 30380 27328
rect 29963 27288 30380 27316
rect 29963 27285 29975 27288
rect 29917 27279 29975 27285
rect 30374 27276 30380 27288
rect 30432 27276 30438 27328
rect 32214 27276 32220 27328
rect 32272 27276 32278 27328
rect 34256 27316 34284 27356
rect 35526 27344 35532 27396
rect 35584 27384 35590 27396
rect 35820 27384 35848 27415
rect 36538 27412 36544 27424
rect 36596 27412 36602 27464
rect 36633 27455 36691 27461
rect 36633 27421 36645 27455
rect 36679 27452 36691 27455
rect 36740 27452 36768 27560
rect 37090 27548 37096 27600
rect 37148 27588 37154 27600
rect 37553 27591 37611 27597
rect 37553 27588 37565 27591
rect 37148 27560 37565 27588
rect 37148 27548 37154 27560
rect 37553 27557 37565 27560
rect 37599 27557 37611 27591
rect 37553 27551 37611 27557
rect 37734 27548 37740 27600
rect 37792 27588 37798 27600
rect 39942 27588 39948 27600
rect 37792 27560 39948 27588
rect 37792 27548 37798 27560
rect 39942 27548 39948 27560
rect 40000 27588 40006 27600
rect 40221 27591 40279 27597
rect 40221 27588 40233 27591
rect 40000 27560 40233 27588
rect 40000 27548 40006 27560
rect 40221 27557 40233 27560
rect 40267 27557 40279 27591
rect 40221 27551 40279 27557
rect 41138 27548 41144 27600
rect 41196 27588 41202 27600
rect 41524 27588 41552 27628
rect 42337 27625 42349 27628
rect 42383 27625 42395 27659
rect 42337 27619 42395 27625
rect 41196 27560 41552 27588
rect 41196 27548 41202 27560
rect 42058 27548 42064 27600
rect 42116 27588 42122 27600
rect 43073 27591 43131 27597
rect 43073 27588 43085 27591
rect 42116 27560 43085 27588
rect 42116 27548 42122 27560
rect 43073 27557 43085 27560
rect 43119 27557 43131 27591
rect 43073 27551 43131 27557
rect 38378 27480 38384 27532
rect 38436 27480 38442 27532
rect 41230 27520 41236 27532
rect 38488 27492 38700 27520
rect 36998 27452 37004 27464
rect 36679 27424 37004 27452
rect 36679 27421 36691 27424
rect 36633 27415 36691 27421
rect 36998 27412 37004 27424
rect 37056 27412 37062 27464
rect 37921 27455 37979 27461
rect 37921 27421 37933 27455
rect 37967 27452 37979 27455
rect 38010 27452 38016 27464
rect 37967 27424 38016 27452
rect 37967 27421 37979 27424
rect 37921 27415 37979 27421
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 38102 27412 38108 27464
rect 38160 27452 38166 27464
rect 38488 27452 38516 27492
rect 38160 27424 38516 27452
rect 38160 27412 38166 27424
rect 38562 27412 38568 27464
rect 38620 27412 38626 27464
rect 38672 27461 38700 27492
rect 40420 27492 41236 27520
rect 38657 27455 38715 27461
rect 38657 27421 38669 27455
rect 38703 27421 38715 27455
rect 38657 27415 38715 27421
rect 39301 27455 39359 27461
rect 39301 27421 39313 27455
rect 39347 27421 39359 27455
rect 39301 27415 39359 27421
rect 35584 27356 35848 27384
rect 37737 27387 37795 27393
rect 35584 27344 35590 27356
rect 37737 27353 37749 27387
rect 37783 27384 37795 27387
rect 39022 27384 39028 27396
rect 37783 27356 39028 27384
rect 37783 27353 37795 27356
rect 37737 27347 37795 27353
rect 39022 27344 39028 27356
rect 39080 27344 39086 27396
rect 39316 27384 39344 27415
rect 39482 27412 39488 27464
rect 39540 27412 39546 27464
rect 40420 27461 40448 27492
rect 41230 27480 41236 27492
rect 41288 27520 41294 27532
rect 42429 27523 42487 27529
rect 42429 27520 42441 27523
rect 41288 27492 42441 27520
rect 41288 27480 41294 27492
rect 40405 27455 40463 27461
rect 40405 27421 40417 27455
rect 40451 27421 40463 27455
rect 40405 27415 40463 27421
rect 40862 27412 40868 27464
rect 40920 27452 40926 27464
rect 40957 27455 41015 27461
rect 40957 27452 40969 27455
rect 40920 27424 40969 27452
rect 40920 27412 40926 27424
rect 40957 27421 40969 27424
rect 41003 27452 41015 27455
rect 41046 27452 41052 27464
rect 41003 27424 41052 27452
rect 41003 27421 41015 27424
rect 40957 27415 41015 27421
rect 41046 27412 41052 27424
rect 41104 27412 41110 27464
rect 41325 27455 41383 27461
rect 41325 27421 41337 27455
rect 41371 27452 41383 27455
rect 41506 27452 41512 27464
rect 41371 27424 41512 27452
rect 41371 27421 41383 27424
rect 41325 27415 41383 27421
rect 41506 27412 41512 27424
rect 41564 27412 41570 27464
rect 41616 27461 41644 27492
rect 42429 27489 42441 27492
rect 42475 27520 42487 27523
rect 42475 27492 43208 27520
rect 42475 27489 42487 27492
rect 42429 27483 42487 27489
rect 41601 27455 41659 27461
rect 41601 27421 41613 27455
rect 41647 27421 41659 27455
rect 41601 27415 41659 27421
rect 42521 27455 42579 27461
rect 42521 27421 42533 27455
rect 42567 27452 42579 27455
rect 42610 27452 42616 27464
rect 42567 27424 42616 27452
rect 42567 27421 42579 27424
rect 42521 27415 42579 27421
rect 42610 27412 42616 27424
rect 42668 27412 42674 27464
rect 43180 27461 43208 27492
rect 42981 27455 43039 27461
rect 42981 27421 42993 27455
rect 43027 27421 43039 27455
rect 42981 27415 43039 27421
rect 43165 27455 43223 27461
rect 43165 27421 43177 27455
rect 43211 27421 43223 27455
rect 43165 27415 43223 27421
rect 40218 27384 40224 27396
rect 39316 27356 40224 27384
rect 34974 27316 34980 27328
rect 34256 27288 34980 27316
rect 34974 27276 34980 27288
rect 35032 27276 35038 27328
rect 35069 27319 35127 27325
rect 35069 27285 35081 27319
rect 35115 27316 35127 27319
rect 35158 27316 35164 27328
rect 35115 27288 35164 27316
rect 35115 27285 35127 27288
rect 35069 27279 35127 27285
rect 35158 27276 35164 27288
rect 35216 27276 35222 27328
rect 36354 27276 36360 27328
rect 36412 27276 36418 27328
rect 36446 27276 36452 27328
rect 36504 27316 36510 27328
rect 38381 27319 38439 27325
rect 38381 27316 38393 27319
rect 36504 27288 38393 27316
rect 36504 27276 36510 27288
rect 38381 27285 38393 27288
rect 38427 27285 38439 27319
rect 38381 27279 38439 27285
rect 38470 27276 38476 27328
rect 38528 27316 38534 27328
rect 39316 27316 39344 27356
rect 40218 27344 40224 27356
rect 40276 27344 40282 27396
rect 41064 27384 41092 27412
rect 41782 27384 41788 27396
rect 41064 27356 41788 27384
rect 41782 27344 41788 27356
rect 41840 27384 41846 27396
rect 42996 27384 43024 27415
rect 41840 27356 43024 27384
rect 41840 27344 41846 27356
rect 38528 27288 39344 27316
rect 38528 27276 38534 27288
rect 40494 27276 40500 27328
rect 40552 27316 40558 27328
rect 41141 27319 41199 27325
rect 41141 27316 41153 27319
rect 40552 27288 41153 27316
rect 40552 27276 40558 27288
rect 41141 27285 41153 27288
rect 41187 27285 41199 27319
rect 41141 27279 41199 27285
rect 41322 27276 41328 27328
rect 41380 27316 41386 27328
rect 42153 27319 42211 27325
rect 42153 27316 42165 27319
rect 41380 27288 42165 27316
rect 41380 27276 41386 27288
rect 42153 27285 42165 27288
rect 42199 27285 42211 27319
rect 42153 27279 42211 27285
rect 1104 27226 43884 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 43884 27226
rect 1104 27152 43884 27174
rect 16209 27115 16267 27121
rect 16209 27081 16221 27115
rect 16255 27112 16267 27115
rect 18138 27112 18144 27124
rect 16255 27084 18144 27112
rect 16255 27081 16267 27084
rect 16209 27075 16267 27081
rect 18138 27072 18144 27084
rect 18196 27072 18202 27124
rect 20714 27072 20720 27124
rect 20772 27112 20778 27124
rect 22005 27115 22063 27121
rect 22005 27112 22017 27115
rect 20772 27084 22017 27112
rect 20772 27072 20778 27084
rect 22005 27081 22017 27084
rect 22051 27081 22063 27115
rect 22005 27075 22063 27081
rect 24673 27115 24731 27121
rect 24673 27081 24685 27115
rect 24719 27112 24731 27115
rect 24946 27112 24952 27124
rect 24719 27084 24952 27112
rect 24719 27081 24731 27084
rect 24673 27075 24731 27081
rect 24946 27072 24952 27084
rect 25004 27072 25010 27124
rect 25682 27072 25688 27124
rect 25740 27072 25746 27124
rect 25774 27072 25780 27124
rect 25832 27112 25838 27124
rect 26053 27115 26111 27121
rect 26053 27112 26065 27115
rect 25832 27084 26065 27112
rect 25832 27072 25838 27084
rect 26053 27081 26065 27084
rect 26099 27081 26111 27115
rect 26053 27075 26111 27081
rect 29178 27072 29184 27124
rect 29236 27072 29242 27124
rect 30374 27072 30380 27124
rect 30432 27072 30438 27124
rect 30834 27072 30840 27124
rect 30892 27112 30898 27124
rect 31757 27115 31815 27121
rect 31757 27112 31769 27115
rect 30892 27084 31769 27112
rect 30892 27072 30898 27084
rect 31757 27081 31769 27084
rect 31803 27081 31815 27115
rect 31757 27075 31815 27081
rect 32214 27072 32220 27124
rect 32272 27112 32278 27124
rect 32401 27115 32459 27121
rect 32401 27112 32413 27115
rect 32272 27084 32413 27112
rect 32272 27072 32278 27084
rect 32401 27081 32413 27084
rect 32447 27081 32459 27115
rect 32401 27075 32459 27081
rect 35437 27115 35495 27121
rect 35437 27081 35449 27115
rect 35483 27112 35495 27115
rect 35802 27112 35808 27124
rect 35483 27084 35808 27112
rect 35483 27081 35495 27084
rect 35437 27075 35495 27081
rect 35802 27072 35808 27084
rect 35860 27072 35866 27124
rect 36170 27072 36176 27124
rect 36228 27072 36234 27124
rect 36538 27072 36544 27124
rect 36596 27112 36602 27124
rect 40678 27112 40684 27124
rect 36596 27084 40684 27112
rect 36596 27072 36602 27084
rect 40678 27072 40684 27084
rect 40736 27072 40742 27124
rect 42610 27072 42616 27124
rect 42668 27072 42674 27124
rect 17120 27047 17178 27053
rect 17120 27013 17132 27047
rect 17166 27044 17178 27047
rect 17218 27044 17224 27056
rect 17166 27016 17224 27044
rect 17166 27013 17178 27016
rect 17120 27007 17178 27013
rect 17218 27004 17224 27016
rect 17276 27004 17282 27056
rect 20438 27004 20444 27056
rect 20496 27044 20502 27056
rect 22830 27044 22836 27056
rect 20496 27016 22836 27044
rect 20496 27004 20502 27016
rect 22830 27004 22836 27016
rect 22888 27004 22894 27056
rect 22922 27004 22928 27056
rect 22980 27044 22986 27056
rect 23017 27047 23075 27053
rect 23017 27044 23029 27047
rect 22980 27016 23029 27044
rect 22980 27004 22986 27016
rect 23017 27013 23029 27016
rect 23063 27044 23075 27047
rect 28534 27044 28540 27056
rect 23063 27016 23704 27044
rect 23063 27013 23075 27016
rect 23017 27007 23075 27013
rect 23676 26988 23704 27016
rect 28368 27016 28540 27044
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 14660 26948 16865 26976
rect 14274 26868 14280 26920
rect 14332 26908 14338 26920
rect 14660 26917 14688 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 20622 26976 20628 26988
rect 19567 26948 20628 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 20622 26936 20628 26948
rect 20680 26936 20686 26988
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 14645 26911 14703 26917
rect 14645 26908 14657 26911
rect 14332 26880 14657 26908
rect 14332 26868 14338 26880
rect 14645 26877 14657 26880
rect 14691 26877 14703 26911
rect 14645 26871 14703 26877
rect 14826 26868 14832 26920
rect 14884 26908 14890 26920
rect 14921 26911 14979 26917
rect 14921 26908 14933 26911
rect 14884 26880 14933 26908
rect 14884 26868 14890 26880
rect 14921 26877 14933 26880
rect 14967 26877 14979 26911
rect 14921 26871 14979 26877
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26908 19671 26911
rect 20254 26908 20260 26920
rect 19659 26880 20260 26908
rect 19659 26877 19671 26880
rect 19613 26871 19671 26877
rect 20254 26868 20260 26880
rect 20312 26908 20318 26920
rect 21361 26911 21419 26917
rect 21361 26908 21373 26911
rect 20312 26880 21373 26908
rect 20312 26868 20318 26880
rect 21361 26877 21373 26880
rect 21407 26908 21419 26911
rect 21407 26880 22094 26908
rect 21407 26877 21419 26880
rect 21361 26871 21419 26877
rect 18233 26775 18291 26781
rect 18233 26741 18245 26775
rect 18279 26772 18291 26775
rect 18506 26772 18512 26784
rect 18279 26744 18512 26772
rect 18279 26741 18291 26744
rect 18233 26735 18291 26741
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 19794 26732 19800 26784
rect 19852 26732 19858 26784
rect 22066 26772 22094 26880
rect 22204 26840 22232 26939
rect 23382 26936 23388 26988
rect 23440 26976 23446 26988
rect 23477 26979 23535 26985
rect 23477 26976 23489 26979
rect 23440 26948 23489 26976
rect 23440 26936 23446 26948
rect 23477 26945 23489 26948
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 23658 26936 23664 26988
rect 23716 26936 23722 26988
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24820 26948 24869 26976
rect 24820 26936 24826 26948
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 26326 26936 26332 26988
rect 26384 26976 26390 26988
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26384 26948 27169 26976
rect 26384 26936 26390 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27246 26936 27252 26988
rect 27304 26976 27310 26988
rect 27341 26979 27399 26985
rect 27341 26976 27353 26979
rect 27304 26948 27353 26976
rect 27304 26936 27310 26948
rect 27341 26945 27353 26948
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 22370 26868 22376 26920
rect 22428 26868 22434 26920
rect 25038 26868 25044 26920
rect 25096 26868 25102 26920
rect 26142 26868 26148 26920
rect 26200 26868 26206 26920
rect 26234 26868 26240 26920
rect 26292 26868 26298 26920
rect 28092 26908 28120 26939
rect 28166 26936 28172 26988
rect 28224 26936 28230 26988
rect 28368 26985 28396 27016
rect 28534 27004 28540 27016
rect 28592 27004 28598 27056
rect 29687 27047 29745 27053
rect 29687 27013 29699 27047
rect 29733 27044 29745 27047
rect 29822 27044 29828 27056
rect 29733 27016 29828 27044
rect 29733 27013 29745 27016
rect 29687 27007 29745 27013
rect 29822 27004 29828 27016
rect 29880 27004 29886 27056
rect 31386 27004 31392 27056
rect 31444 27004 31450 27056
rect 31938 27004 31944 27056
rect 31996 27044 32002 27056
rect 32674 27044 32680 27056
rect 31996 27016 32680 27044
rect 31996 27004 32002 27016
rect 28353 26979 28411 26985
rect 28353 26945 28365 26979
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 28442 26936 28448 26988
rect 28500 26936 28506 26988
rect 29362 26976 29368 26988
rect 28966 26948 29368 26976
rect 28966 26908 28994 26948
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 29454 26936 29460 26988
rect 29512 26936 29518 26988
rect 29546 26936 29552 26988
rect 29604 26936 29610 26988
rect 30285 26979 30343 26985
rect 30285 26976 30297 26979
rect 29840 26948 30297 26976
rect 29840 26920 29868 26948
rect 30285 26945 30297 26948
rect 30331 26945 30343 26979
rect 30285 26939 30343 26945
rect 31573 26979 31631 26985
rect 31573 26945 31585 26979
rect 31619 26976 31631 26979
rect 31662 26976 31668 26988
rect 31619 26948 31668 26976
rect 31619 26945 31631 26948
rect 31573 26939 31631 26945
rect 31662 26936 31668 26948
rect 31720 26936 31726 26988
rect 32324 26985 32352 27016
rect 32674 27004 32680 27016
rect 32732 27004 32738 27056
rect 33962 27044 33968 27056
rect 33060 27016 33968 27044
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 32493 26979 32551 26985
rect 32493 26945 32505 26979
rect 32539 26976 32551 26979
rect 33060 26976 33088 27016
rect 33962 27004 33968 27016
rect 34020 27044 34026 27056
rect 34698 27044 34704 27056
rect 34020 27016 34704 27044
rect 34020 27004 34026 27016
rect 34698 27004 34704 27016
rect 34756 27004 34762 27056
rect 37090 27004 37096 27056
rect 37148 27044 37154 27056
rect 38378 27044 38384 27056
rect 37148 27016 37872 27044
rect 37148 27004 37154 27016
rect 32539 26948 33088 26976
rect 33137 26979 33195 26985
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 33137 26945 33149 26979
rect 33183 26945 33195 26979
rect 33137 26939 33195 26945
rect 33321 26979 33379 26985
rect 33321 26945 33333 26979
rect 33367 26976 33379 26979
rect 33502 26976 33508 26988
rect 33367 26948 33508 26976
rect 33367 26945 33379 26948
rect 33321 26939 33379 26945
rect 28092 26880 28994 26908
rect 28092 26840 28120 26880
rect 29822 26868 29828 26920
rect 29880 26868 29886 26920
rect 33152 26908 33180 26939
rect 33502 26936 33508 26948
rect 33560 26936 33566 26988
rect 34238 26936 34244 26988
rect 34296 26936 34302 26988
rect 34790 26936 34796 26988
rect 34848 26976 34854 26988
rect 35069 26979 35127 26985
rect 35069 26976 35081 26979
rect 34848 26948 35081 26976
rect 34848 26936 34854 26948
rect 35069 26945 35081 26948
rect 35115 26945 35127 26979
rect 35069 26939 35127 26945
rect 35158 26936 35164 26988
rect 35216 26936 35222 26988
rect 36354 26936 36360 26988
rect 36412 26936 36418 26988
rect 36725 26979 36783 26985
rect 36725 26976 36737 26979
rect 36464 26948 36737 26976
rect 34057 26911 34115 26917
rect 34057 26908 34069 26911
rect 33152 26880 33916 26908
rect 33888 26852 33916 26880
rect 33980 26880 34069 26908
rect 22204 26812 28120 26840
rect 32398 26800 32404 26852
rect 32456 26840 32462 26852
rect 33042 26840 33048 26852
rect 32456 26812 33048 26840
rect 32456 26800 32462 26812
rect 33042 26800 33048 26812
rect 33100 26840 33106 26852
rect 33100 26812 33824 26840
rect 33100 26800 33106 26812
rect 22738 26772 22744 26784
rect 22066 26744 22744 26772
rect 22738 26732 22744 26744
rect 22796 26732 22802 26784
rect 23474 26732 23480 26784
rect 23532 26732 23538 26784
rect 23845 26775 23903 26781
rect 23845 26741 23857 26775
rect 23891 26772 23903 26775
rect 24486 26772 24492 26784
rect 23891 26744 24492 26772
rect 23891 26741 23903 26744
rect 23845 26735 23903 26741
rect 24486 26732 24492 26744
rect 24544 26732 24550 26784
rect 27062 26732 27068 26784
rect 27120 26772 27126 26784
rect 27157 26775 27215 26781
rect 27157 26772 27169 26775
rect 27120 26744 27169 26772
rect 27120 26732 27126 26744
rect 27157 26741 27169 26744
rect 27203 26741 27215 26775
rect 27157 26735 27215 26741
rect 27798 26732 27804 26784
rect 27856 26772 27862 26784
rect 27893 26775 27951 26781
rect 27893 26772 27905 26775
rect 27856 26744 27905 26772
rect 27856 26732 27862 26744
rect 27893 26741 27905 26744
rect 27939 26741 27951 26775
rect 27893 26735 27951 26741
rect 33134 26732 33140 26784
rect 33192 26732 33198 26784
rect 33796 26772 33824 26812
rect 33870 26800 33876 26852
rect 33928 26800 33934 26852
rect 33980 26840 34008 26880
rect 34057 26877 34069 26880
rect 34103 26877 34115 26911
rect 34057 26871 34115 26877
rect 34149 26911 34207 26917
rect 34149 26877 34161 26911
rect 34195 26908 34207 26911
rect 34330 26908 34336 26920
rect 34195 26880 34336 26908
rect 34195 26877 34207 26880
rect 34149 26871 34207 26877
rect 34330 26868 34336 26880
rect 34388 26868 34394 26920
rect 36170 26868 36176 26920
rect 36228 26908 36234 26920
rect 36464 26908 36492 26948
rect 36725 26945 36737 26948
rect 36771 26945 36783 26979
rect 36725 26939 36783 26945
rect 37734 26936 37740 26988
rect 37792 26936 37798 26988
rect 37844 26985 37872 27016
rect 38120 27016 38384 27044
rect 37829 26979 37887 26985
rect 37829 26945 37841 26979
rect 37875 26945 37887 26979
rect 37829 26939 37887 26945
rect 37918 26936 37924 26988
rect 37976 26936 37982 26988
rect 38120 26985 38148 27016
rect 38378 27004 38384 27016
rect 38436 27004 38442 27056
rect 39390 27004 39396 27056
rect 39448 27004 39454 27056
rect 39485 27047 39543 27053
rect 39485 27013 39497 27047
rect 39531 27044 39543 27047
rect 39850 27044 39856 27056
rect 39531 27016 39856 27044
rect 39531 27013 39543 27016
rect 39485 27007 39543 27013
rect 39850 27004 39856 27016
rect 39908 27004 39914 27056
rect 41969 27047 42027 27053
rect 41969 27044 41981 27047
rect 41248 27016 41981 27044
rect 38105 26979 38163 26985
rect 38105 26945 38117 26979
rect 38151 26945 38163 26979
rect 38105 26939 38163 26945
rect 38286 26936 38292 26988
rect 38344 26976 38350 26988
rect 38933 26979 38991 26985
rect 38933 26976 38945 26979
rect 38344 26948 38945 26976
rect 38344 26936 38350 26948
rect 38933 26945 38945 26948
rect 38979 26945 38991 26979
rect 38933 26939 38991 26945
rect 39761 26979 39819 26985
rect 39761 26945 39773 26979
rect 39807 26976 39819 26979
rect 40034 26976 40040 26988
rect 39807 26948 40040 26976
rect 39807 26945 39819 26948
rect 39761 26939 39819 26945
rect 40034 26936 40040 26948
rect 40092 26936 40098 26988
rect 40218 26936 40224 26988
rect 40276 26976 40282 26988
rect 40954 26976 40960 26988
rect 40276 26948 40960 26976
rect 40276 26936 40282 26948
rect 40954 26936 40960 26948
rect 41012 26976 41018 26988
rect 41141 26979 41199 26985
rect 41141 26976 41153 26979
rect 41012 26948 41153 26976
rect 41012 26936 41018 26948
rect 41141 26945 41153 26948
rect 41187 26945 41199 26979
rect 41141 26939 41199 26945
rect 36228 26880 36492 26908
rect 36228 26868 36234 26880
rect 36630 26868 36636 26920
rect 36688 26908 36694 26920
rect 36817 26911 36875 26917
rect 36817 26908 36829 26911
rect 36688 26880 36829 26908
rect 36688 26868 36694 26880
rect 36817 26877 36829 26880
rect 36863 26877 36875 26911
rect 36817 26871 36875 26877
rect 36924 26880 38332 26908
rect 34422 26840 34428 26852
rect 33980 26812 34428 26840
rect 33980 26772 34008 26812
rect 34422 26800 34428 26812
rect 34480 26800 34486 26852
rect 35802 26800 35808 26852
rect 35860 26840 35866 26852
rect 36924 26840 36952 26880
rect 35860 26812 36952 26840
rect 35860 26800 35866 26812
rect 36998 26800 37004 26852
rect 37056 26840 37062 26852
rect 37734 26840 37740 26852
rect 37056 26812 37740 26840
rect 37056 26800 37062 26812
rect 37734 26800 37740 26812
rect 37792 26800 37798 26852
rect 38304 26840 38332 26880
rect 38470 26868 38476 26920
rect 38528 26908 38534 26920
rect 38746 26908 38752 26920
rect 38528 26880 38752 26908
rect 38528 26868 38534 26880
rect 38746 26868 38752 26880
rect 38804 26908 38810 26920
rect 38841 26911 38899 26917
rect 38841 26908 38853 26911
rect 38804 26880 38853 26908
rect 38804 26868 38810 26880
rect 38841 26877 38853 26880
rect 38887 26877 38899 26911
rect 38841 26871 38899 26877
rect 39206 26868 39212 26920
rect 39264 26908 39270 26920
rect 39853 26911 39911 26917
rect 39853 26908 39865 26911
rect 39264 26880 39865 26908
rect 39264 26868 39270 26880
rect 39853 26877 39865 26880
rect 39899 26877 39911 26911
rect 39853 26871 39911 26877
rect 40310 26868 40316 26920
rect 40368 26908 40374 26920
rect 40862 26908 40868 26920
rect 40368 26880 40868 26908
rect 40368 26868 40374 26880
rect 40862 26868 40868 26880
rect 40920 26908 40926 26920
rect 41049 26911 41107 26917
rect 41049 26908 41061 26911
rect 40920 26880 41061 26908
rect 40920 26868 40926 26880
rect 41049 26877 41061 26880
rect 41095 26877 41107 26911
rect 41049 26871 41107 26877
rect 39114 26840 39120 26852
rect 38304 26812 39120 26840
rect 39114 26800 39120 26812
rect 39172 26800 39178 26852
rect 39574 26800 39580 26852
rect 39632 26840 39638 26852
rect 41248 26840 41276 27016
rect 41969 27013 41981 27016
rect 42015 27044 42027 27047
rect 43346 27044 43352 27056
rect 42015 27016 43352 27044
rect 42015 27013 42027 27016
rect 41969 27007 42027 27013
rect 43346 27004 43352 27016
rect 43404 27004 43410 27056
rect 41506 26936 41512 26988
rect 41564 26976 41570 26988
rect 41564 26948 42472 26976
rect 41564 26936 41570 26948
rect 41414 26868 41420 26920
rect 41472 26908 41478 26920
rect 41601 26911 41659 26917
rect 41601 26908 41613 26911
rect 41472 26880 41613 26908
rect 41472 26868 41478 26880
rect 41601 26877 41613 26880
rect 41647 26877 41659 26911
rect 41601 26871 41659 26877
rect 39632 26812 41276 26840
rect 39632 26800 39638 26812
rect 42444 26784 42472 26948
rect 43070 26936 43076 26988
rect 43128 26936 43134 26988
rect 33796 26744 34008 26772
rect 34054 26732 34060 26784
rect 34112 26732 34118 26784
rect 34698 26732 34704 26784
rect 34756 26772 34762 26784
rect 35069 26775 35127 26781
rect 35069 26772 35081 26775
rect 34756 26744 35081 26772
rect 34756 26732 34762 26744
rect 35069 26741 35081 26744
rect 35115 26741 35127 26775
rect 35069 26735 35127 26741
rect 36357 26775 36415 26781
rect 36357 26741 36369 26775
rect 36403 26772 36415 26775
rect 36446 26772 36452 26784
rect 36403 26744 36452 26772
rect 36403 26741 36415 26744
rect 36357 26735 36415 26741
rect 36446 26732 36452 26744
rect 36504 26732 36510 26784
rect 37274 26732 37280 26784
rect 37332 26772 37338 26784
rect 37461 26775 37519 26781
rect 37461 26772 37473 26775
rect 37332 26744 37473 26772
rect 37332 26732 37338 26744
rect 37461 26741 37473 26744
rect 37507 26741 37519 26775
rect 37461 26735 37519 26741
rect 38102 26732 38108 26784
rect 38160 26772 38166 26784
rect 38565 26775 38623 26781
rect 38565 26772 38577 26775
rect 38160 26744 38577 26772
rect 38160 26732 38166 26744
rect 38565 26741 38577 26744
rect 38611 26741 38623 26775
rect 38565 26735 38623 26741
rect 38838 26732 38844 26784
rect 38896 26732 38902 26784
rect 40037 26775 40095 26781
rect 40037 26741 40049 26775
rect 40083 26772 40095 26775
rect 40218 26772 40224 26784
rect 40083 26744 40224 26772
rect 40083 26741 40095 26744
rect 40037 26735 40095 26741
rect 40218 26732 40224 26744
rect 40276 26732 40282 26784
rect 41230 26732 41236 26784
rect 41288 26772 41294 26784
rect 41509 26775 41567 26781
rect 41509 26772 41521 26775
rect 41288 26744 41521 26772
rect 41288 26732 41294 26744
rect 41509 26741 41521 26744
rect 41555 26741 41567 26775
rect 41509 26735 41567 26741
rect 42426 26732 42432 26784
rect 42484 26772 42490 26784
rect 42797 26775 42855 26781
rect 42797 26772 42809 26775
rect 42484 26744 42809 26772
rect 42484 26732 42490 26744
rect 42797 26741 42809 26744
rect 42843 26741 42855 26775
rect 42797 26735 42855 26741
rect 1104 26682 43884 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 43884 26682
rect 1104 26608 43884 26630
rect 21637 26571 21695 26577
rect 21637 26537 21649 26571
rect 21683 26568 21695 26571
rect 22830 26568 22836 26580
rect 21683 26540 22836 26568
rect 21683 26537 21695 26540
rect 21637 26531 21695 26537
rect 22830 26528 22836 26540
rect 22888 26528 22894 26580
rect 23566 26528 23572 26580
rect 23624 26568 23630 26580
rect 25777 26571 25835 26577
rect 25777 26568 25789 26571
rect 23624 26540 25789 26568
rect 23624 26528 23630 26540
rect 25777 26537 25789 26540
rect 25823 26568 25835 26571
rect 25866 26568 25872 26580
rect 25823 26540 25872 26568
rect 25823 26537 25835 26540
rect 25777 26531 25835 26537
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 26142 26528 26148 26580
rect 26200 26568 26206 26580
rect 26697 26571 26755 26577
rect 26697 26568 26709 26571
rect 26200 26540 26709 26568
rect 26200 26528 26206 26540
rect 26697 26537 26709 26540
rect 26743 26537 26755 26571
rect 26697 26531 26755 26537
rect 29546 26528 29552 26580
rect 29604 26568 29610 26580
rect 29825 26571 29883 26577
rect 29825 26568 29837 26571
rect 29604 26540 29837 26568
rect 29604 26528 29610 26540
rect 29825 26537 29837 26540
rect 29871 26537 29883 26571
rect 29825 26531 29883 26537
rect 30558 26528 30564 26580
rect 30616 26528 30622 26580
rect 31478 26528 31484 26580
rect 31536 26568 31542 26580
rect 32769 26571 32827 26577
rect 32769 26568 32781 26571
rect 31536 26540 32781 26568
rect 31536 26528 31542 26540
rect 32769 26537 32781 26540
rect 32815 26537 32827 26571
rect 32769 26531 32827 26537
rect 34514 26528 34520 26580
rect 34572 26568 34578 26580
rect 35713 26571 35771 26577
rect 35713 26568 35725 26571
rect 34572 26540 35725 26568
rect 34572 26528 34578 26540
rect 35713 26537 35725 26540
rect 35759 26537 35771 26571
rect 35713 26531 35771 26537
rect 36817 26571 36875 26577
rect 36817 26537 36829 26571
rect 36863 26568 36875 26571
rect 37090 26568 37096 26580
rect 36863 26540 37096 26568
rect 36863 26537 36875 26540
rect 36817 26531 36875 26537
rect 37090 26528 37096 26540
rect 37148 26528 37154 26580
rect 41325 26571 41383 26577
rect 41325 26568 41337 26571
rect 37844 26540 41337 26568
rect 15657 26503 15715 26509
rect 15657 26469 15669 26503
rect 15703 26469 15715 26503
rect 15657 26463 15715 26469
rect 20073 26503 20131 26509
rect 20073 26469 20085 26503
rect 20119 26500 20131 26503
rect 20346 26500 20352 26512
rect 20119 26472 20352 26500
rect 20119 26469 20131 26472
rect 20073 26463 20131 26469
rect 15672 26432 15700 26463
rect 20346 26460 20352 26472
rect 20404 26460 20410 26512
rect 20622 26460 20628 26512
rect 20680 26500 20686 26512
rect 20993 26503 21051 26509
rect 20993 26500 21005 26503
rect 20680 26472 21005 26500
rect 20680 26460 20686 26472
rect 20993 26469 21005 26472
rect 21039 26500 21051 26503
rect 26050 26500 26056 26512
rect 21039 26472 26056 26500
rect 21039 26469 21051 26472
rect 20993 26463 21051 26469
rect 15672 26404 17540 26432
rect 14274 26324 14280 26376
rect 14332 26364 14338 26376
rect 15286 26364 15292 26376
rect 14332 26336 15292 26364
rect 14332 26324 14338 26336
rect 15286 26324 15292 26336
rect 15344 26364 15350 26376
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 15344 26336 17417 26364
rect 15344 26324 15350 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 17512 26364 17540 26404
rect 19794 26392 19800 26444
rect 19852 26392 19858 26444
rect 22557 26435 22615 26441
rect 22557 26401 22569 26435
rect 22603 26432 22615 26435
rect 23382 26432 23388 26444
rect 22603 26404 23388 26432
rect 22603 26401 22615 26404
rect 22557 26395 22615 26401
rect 23382 26392 23388 26404
rect 23440 26432 23446 26444
rect 23569 26435 23627 26441
rect 23569 26432 23581 26435
rect 23440 26404 23581 26432
rect 23440 26392 23446 26404
rect 23569 26401 23581 26404
rect 23615 26401 23627 26435
rect 23569 26395 23627 26401
rect 17512 26336 19288 26364
rect 17405 26327 17463 26333
rect 14292 26296 14320 26324
rect 13740 26268 14320 26296
rect 13262 26188 13268 26240
rect 13320 26228 13326 26240
rect 13740 26228 13768 26268
rect 14366 26256 14372 26308
rect 14424 26296 14430 26308
rect 14522 26299 14580 26305
rect 14522 26296 14534 26299
rect 14424 26268 14534 26296
rect 14424 26256 14430 26268
rect 14522 26265 14534 26268
rect 14568 26265 14580 26299
rect 14522 26259 14580 26265
rect 17672 26299 17730 26305
rect 17672 26265 17684 26299
rect 17718 26296 17730 26299
rect 17770 26296 17776 26308
rect 17718 26268 17776 26296
rect 17718 26265 17730 26268
rect 17672 26259 17730 26265
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 19260 26296 19288 26336
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19705 26367 19763 26373
rect 19705 26364 19717 26367
rect 19392 26336 19717 26364
rect 19392 26324 19398 26336
rect 19705 26333 19717 26336
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 22462 26324 22468 26376
rect 22520 26324 22526 26376
rect 22649 26367 22707 26373
rect 22649 26333 22661 26367
rect 22695 26364 22707 26367
rect 22738 26364 22744 26376
rect 22695 26336 22744 26364
rect 22695 26333 22707 26336
rect 22649 26327 22707 26333
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23676 26373 23704 26472
rect 26050 26460 26056 26472
rect 26108 26460 26114 26512
rect 26237 26503 26295 26509
rect 26237 26469 26249 26503
rect 26283 26500 26295 26503
rect 26326 26500 26332 26512
rect 26283 26472 26332 26500
rect 26283 26469 26295 26472
rect 26237 26463 26295 26469
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 27893 26503 27951 26509
rect 27893 26500 27905 26503
rect 27172 26472 27905 26500
rect 24854 26392 24860 26444
rect 24912 26432 24918 26444
rect 25958 26432 25964 26444
rect 24912 26404 25964 26432
rect 24912 26392 24918 26404
rect 25958 26392 25964 26404
rect 26016 26392 26022 26444
rect 27172 26441 27200 26472
rect 27893 26469 27905 26472
rect 27939 26469 27951 26503
rect 27893 26463 27951 26469
rect 31726 26472 33824 26500
rect 27157 26435 27215 26441
rect 27157 26401 27169 26435
rect 27203 26401 27215 26435
rect 27157 26395 27215 26401
rect 27338 26392 27344 26444
rect 27396 26392 27402 26444
rect 27982 26392 27988 26444
rect 28040 26432 28046 26444
rect 28442 26432 28448 26444
rect 28040 26404 28448 26432
rect 28040 26392 28046 26404
rect 28442 26392 28448 26404
rect 28500 26392 28506 26444
rect 29086 26392 29092 26444
rect 29144 26432 29150 26444
rect 29144 26404 30052 26432
rect 29144 26392 29150 26404
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26333 23719 26367
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 23661 26327 23719 26333
rect 24596 26336 24961 26364
rect 21266 26296 21272 26308
rect 19260 26268 21272 26296
rect 21266 26256 21272 26268
rect 21324 26296 21330 26308
rect 21605 26299 21663 26305
rect 21605 26296 21617 26299
rect 21324 26268 21617 26296
rect 21324 26256 21330 26268
rect 21605 26265 21617 26268
rect 21651 26265 21663 26299
rect 21605 26259 21663 26265
rect 21821 26299 21879 26305
rect 21821 26265 21833 26299
rect 21867 26296 21879 26299
rect 22370 26296 22376 26308
rect 21867 26268 22376 26296
rect 21867 26265 21879 26268
rect 21821 26259 21879 26265
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 24596 26240 24624 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 25133 26367 25191 26373
rect 25133 26333 25145 26367
rect 25179 26364 25191 26367
rect 25222 26364 25228 26376
rect 25179 26336 25228 26364
rect 25179 26333 25191 26336
rect 25133 26327 25191 26333
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 26053 26367 26111 26373
rect 26053 26364 26065 26367
rect 25648 26336 26065 26364
rect 25648 26324 25654 26336
rect 26053 26333 26065 26336
rect 26099 26364 26111 26367
rect 26142 26364 26148 26376
rect 26099 26336 26148 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 27062 26324 27068 26376
rect 27120 26324 27126 26376
rect 29270 26324 29276 26376
rect 29328 26364 29334 26376
rect 29914 26364 29920 26376
rect 29328 26336 29920 26364
rect 29328 26324 29334 26336
rect 29914 26324 29920 26336
rect 29972 26324 29978 26376
rect 30024 26364 30052 26404
rect 30926 26392 30932 26444
rect 30984 26432 30990 26444
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30984 26404 31125 26432
rect 30984 26392 30990 26404
rect 31113 26401 31125 26404
rect 31159 26432 31171 26435
rect 31726 26432 31754 26472
rect 33134 26432 33140 26444
rect 31159 26404 31754 26432
rect 32968 26404 33140 26432
rect 31159 26401 31171 26404
rect 31113 26395 31171 26401
rect 32968 26373 32996 26404
rect 33134 26392 33140 26404
rect 33192 26392 33198 26444
rect 33796 26432 33824 26472
rect 33870 26460 33876 26512
rect 33928 26500 33934 26512
rect 37844 26500 37872 26540
rect 41325 26537 41337 26540
rect 41371 26537 41383 26571
rect 41325 26531 41383 26537
rect 33928 26472 37872 26500
rect 33928 26460 33934 26472
rect 35728 26444 35756 26472
rect 33796 26404 34928 26432
rect 31757 26367 31815 26373
rect 31757 26364 31769 26367
rect 30024 26336 31769 26364
rect 31757 26333 31769 26336
rect 31803 26333 31815 26367
rect 31757 26327 31815 26333
rect 32953 26367 33011 26373
rect 32953 26333 32965 26367
rect 32999 26333 33011 26367
rect 33597 26367 33655 26373
rect 33597 26364 33609 26367
rect 32953 26327 33011 26333
rect 33060 26336 33609 26364
rect 25774 26256 25780 26308
rect 25832 26256 25838 26308
rect 25866 26256 25872 26308
rect 25924 26296 25930 26308
rect 28261 26299 28319 26305
rect 28261 26296 28273 26299
rect 25924 26268 28273 26296
rect 25924 26256 25930 26268
rect 28261 26265 28273 26268
rect 28307 26296 28319 26299
rect 29086 26296 29092 26308
rect 28307 26268 29092 26296
rect 28307 26265 28319 26268
rect 28261 26259 28319 26265
rect 29086 26256 29092 26268
rect 29144 26256 29150 26308
rect 29178 26256 29184 26308
rect 29236 26256 29242 26308
rect 30650 26256 30656 26308
rect 30708 26296 30714 26308
rect 30929 26299 30987 26305
rect 30929 26296 30941 26299
rect 30708 26268 30941 26296
rect 30708 26256 30714 26268
rect 30929 26265 30941 26268
rect 30975 26265 30987 26299
rect 30929 26259 30987 26265
rect 32674 26256 32680 26308
rect 32732 26296 32738 26308
rect 33060 26296 33088 26336
rect 33597 26333 33609 26336
rect 33643 26333 33655 26367
rect 33597 26327 33655 26333
rect 33778 26324 33784 26376
rect 33836 26324 33842 26376
rect 33873 26367 33931 26373
rect 33873 26333 33885 26367
rect 33919 26333 33931 26367
rect 33873 26327 33931 26333
rect 32732 26268 33088 26296
rect 33137 26299 33195 26305
rect 32732 26256 32738 26268
rect 33137 26265 33149 26299
rect 33183 26296 33195 26299
rect 33226 26296 33232 26308
rect 33183 26268 33232 26296
rect 33183 26265 33195 26268
rect 33137 26259 33195 26265
rect 13320 26200 13768 26228
rect 13320 26188 13326 26200
rect 18598 26188 18604 26240
rect 18656 26228 18662 26240
rect 18785 26231 18843 26237
rect 18785 26228 18797 26231
rect 18656 26200 18797 26228
rect 18656 26188 18662 26200
rect 18785 26197 18797 26200
rect 18831 26197 18843 26231
rect 18785 26191 18843 26197
rect 21450 26188 21456 26240
rect 21508 26188 21514 26240
rect 24029 26231 24087 26237
rect 24029 26197 24041 26231
rect 24075 26228 24087 26231
rect 24578 26228 24584 26240
rect 24075 26200 24584 26228
rect 24075 26197 24087 26200
rect 24029 26191 24087 26197
rect 24578 26188 24584 26200
rect 24636 26188 24642 26240
rect 25041 26231 25099 26237
rect 25041 26197 25053 26231
rect 25087 26228 25099 26231
rect 25682 26228 25688 26240
rect 25087 26200 25688 26228
rect 25087 26197 25099 26200
rect 25041 26191 25099 26197
rect 25682 26188 25688 26200
rect 25740 26188 25746 26240
rect 26050 26188 26056 26240
rect 26108 26228 26114 26240
rect 28353 26231 28411 26237
rect 28353 26228 28365 26231
rect 26108 26200 28365 26228
rect 26108 26188 26114 26200
rect 28353 26197 28365 26200
rect 28399 26228 28411 26231
rect 28994 26228 29000 26240
rect 28399 26200 29000 26228
rect 28399 26197 28411 26200
rect 28353 26191 28411 26197
rect 28994 26188 29000 26200
rect 29052 26188 29058 26240
rect 31018 26188 31024 26240
rect 31076 26188 31082 26240
rect 32306 26188 32312 26240
rect 32364 26228 32370 26240
rect 33152 26228 33180 26259
rect 33226 26256 33232 26268
rect 33284 26256 33290 26308
rect 33502 26256 33508 26308
rect 33560 26296 33566 26308
rect 33888 26296 33916 26327
rect 34054 26324 34060 26376
rect 34112 26364 34118 26376
rect 34606 26364 34612 26376
rect 34112 26336 34612 26364
rect 34112 26324 34118 26336
rect 34606 26324 34612 26336
rect 34664 26324 34670 26376
rect 34900 26373 34928 26404
rect 35710 26392 35716 26444
rect 35768 26392 35774 26444
rect 36909 26435 36967 26441
rect 36909 26401 36921 26435
rect 36955 26432 36967 26435
rect 36998 26432 37004 26444
rect 36955 26404 37004 26432
rect 36955 26401 36967 26404
rect 36909 26395 36967 26401
rect 36998 26392 37004 26404
rect 37056 26392 37062 26444
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26364 34943 26367
rect 36170 26364 36176 26376
rect 34931 26336 36176 26364
rect 34931 26333 34943 26336
rect 34885 26327 34943 26333
rect 36170 26324 36176 26336
rect 36228 26324 36234 26376
rect 36630 26324 36636 26376
rect 36688 26324 36694 26376
rect 35069 26299 35127 26305
rect 35069 26296 35081 26299
rect 33560 26268 35081 26296
rect 33560 26256 33566 26268
rect 35069 26265 35081 26268
rect 35115 26265 35127 26299
rect 35069 26259 35127 26265
rect 34514 26228 34520 26240
rect 32364 26200 34520 26228
rect 32364 26188 32370 26200
rect 34514 26188 34520 26200
rect 34572 26188 34578 26240
rect 35084 26228 35112 26259
rect 35250 26256 35256 26308
rect 35308 26256 35314 26308
rect 36648 26296 36676 26324
rect 37369 26299 37427 26305
rect 37369 26296 37381 26299
rect 36648 26268 37381 26296
rect 37369 26265 37381 26268
rect 37415 26265 37427 26299
rect 37369 26259 37427 26265
rect 37458 26256 37464 26308
rect 37516 26296 37522 26308
rect 37553 26299 37611 26305
rect 37553 26296 37565 26299
rect 37516 26268 37565 26296
rect 37516 26256 37522 26268
rect 37553 26265 37565 26268
rect 37599 26265 37611 26299
rect 37553 26259 37611 26265
rect 37737 26299 37795 26305
rect 37737 26265 37749 26299
rect 37783 26296 37795 26299
rect 37844 26296 37872 26472
rect 38378 26460 38384 26512
rect 38436 26500 38442 26512
rect 38436 26472 38654 26500
rect 38436 26460 38442 26472
rect 38626 26432 38654 26472
rect 38948 26472 40172 26500
rect 38948 26441 38976 26472
rect 38933 26435 38991 26441
rect 38933 26432 38945 26435
rect 38626 26404 38945 26432
rect 38933 26401 38945 26404
rect 38979 26401 38991 26435
rect 38933 26395 38991 26401
rect 39114 26392 39120 26444
rect 39172 26432 39178 26444
rect 39301 26435 39359 26441
rect 39301 26432 39313 26435
rect 39172 26404 39313 26432
rect 39172 26392 39178 26404
rect 39301 26401 39313 26404
rect 39347 26401 39359 26435
rect 39301 26395 39359 26401
rect 38378 26324 38384 26376
rect 38436 26364 38442 26376
rect 38562 26364 38568 26376
rect 38436 26336 38568 26364
rect 38436 26324 38442 26336
rect 38562 26324 38568 26336
rect 38620 26364 38626 26376
rect 39025 26367 39083 26373
rect 39025 26364 39037 26367
rect 38620 26336 39037 26364
rect 38620 26324 38626 26336
rect 39025 26333 39037 26336
rect 39071 26333 39083 26367
rect 39316 26364 39344 26395
rect 39390 26392 39396 26444
rect 39448 26392 39454 26444
rect 40034 26392 40040 26444
rect 40092 26392 40098 26444
rect 40144 26432 40172 26472
rect 40144 26404 40632 26432
rect 39666 26364 39672 26376
rect 39316 26336 39672 26364
rect 39025 26327 39083 26333
rect 39666 26324 39672 26336
rect 39724 26324 39730 26376
rect 39942 26324 39948 26376
rect 40000 26364 40006 26376
rect 40313 26367 40371 26373
rect 40313 26364 40325 26367
rect 40000 26336 40325 26364
rect 40000 26324 40006 26336
rect 40313 26333 40325 26336
rect 40359 26333 40371 26367
rect 40313 26327 40371 26333
rect 40402 26324 40408 26376
rect 40460 26324 40466 26376
rect 40494 26324 40500 26376
rect 40552 26364 40558 26376
rect 40604 26364 40632 26404
rect 41046 26392 41052 26444
rect 41104 26432 41110 26444
rect 41874 26432 41880 26444
rect 41104 26404 41880 26432
rect 41104 26392 41110 26404
rect 41874 26392 41880 26404
rect 41932 26432 41938 26444
rect 43070 26432 43076 26444
rect 41932 26404 43076 26432
rect 41932 26392 41938 26404
rect 40552 26336 40632 26364
rect 40552 26324 40558 26336
rect 40678 26324 40684 26376
rect 40736 26324 40742 26376
rect 40954 26324 40960 26376
rect 41012 26364 41018 26376
rect 41417 26367 41475 26373
rect 41417 26364 41429 26367
rect 41012 26336 41429 26364
rect 41012 26324 41018 26336
rect 41417 26333 41429 26336
rect 41463 26333 41475 26367
rect 41417 26327 41475 26333
rect 37783 26268 37872 26296
rect 41432 26296 41460 26327
rect 41782 26324 41788 26376
rect 41840 26324 41846 26376
rect 42904 26373 42932 26404
rect 43070 26392 43076 26404
rect 43128 26392 43134 26444
rect 42061 26367 42119 26373
rect 42061 26333 42073 26367
rect 42107 26333 42119 26367
rect 42061 26327 42119 26333
rect 42889 26367 42947 26373
rect 42889 26333 42901 26367
rect 42935 26333 42947 26367
rect 42889 26327 42947 26333
rect 41966 26296 41972 26308
rect 41432 26268 41972 26296
rect 37783 26265 37795 26268
rect 37737 26259 37795 26265
rect 41966 26256 41972 26268
rect 42024 26256 42030 26308
rect 35802 26228 35808 26240
rect 35084 26200 35808 26228
rect 35802 26188 35808 26200
rect 35860 26188 35866 26240
rect 35894 26188 35900 26240
rect 35952 26228 35958 26240
rect 36449 26231 36507 26237
rect 36449 26228 36461 26231
rect 35952 26200 36461 26228
rect 35952 26188 35958 26200
rect 36449 26197 36461 26200
rect 36495 26228 36507 26231
rect 37918 26228 37924 26240
rect 36495 26200 37924 26228
rect 36495 26197 36507 26200
rect 36449 26191 36507 26197
rect 37918 26188 37924 26200
rect 37976 26228 37982 26240
rect 38197 26231 38255 26237
rect 38197 26228 38209 26231
rect 37976 26200 38209 26228
rect 37976 26188 37982 26200
rect 38197 26197 38209 26200
rect 38243 26197 38255 26231
rect 38197 26191 38255 26197
rect 38746 26188 38752 26240
rect 38804 26188 38810 26240
rect 41230 26188 41236 26240
rect 41288 26228 41294 26240
rect 42076 26228 42104 26327
rect 41288 26200 42104 26228
rect 41288 26188 41294 26200
rect 1104 26138 43884 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 43884 26138
rect 1104 26064 43884 26086
rect 19613 26027 19671 26033
rect 19613 25993 19625 26027
rect 19659 26024 19671 26027
rect 20530 26024 20536 26036
rect 19659 25996 20536 26024
rect 19659 25993 19671 25996
rect 19613 25987 19671 25993
rect 20530 25984 20536 25996
rect 20588 25984 20594 26036
rect 22005 26027 22063 26033
rect 22005 25993 22017 26027
rect 22051 26024 22063 26027
rect 22462 26024 22468 26036
rect 22051 25996 22468 26024
rect 22051 25993 22063 25996
rect 22005 25987 22063 25993
rect 20438 25916 20444 25968
rect 20496 25916 20502 25968
rect 13716 25891 13774 25897
rect 13716 25857 13728 25891
rect 13762 25888 13774 25891
rect 14274 25888 14280 25900
rect 13762 25860 14280 25888
rect 13762 25857 13774 25860
rect 13716 25851 13774 25857
rect 14274 25848 14280 25860
rect 14332 25848 14338 25900
rect 15838 25848 15844 25900
rect 15896 25848 15902 25900
rect 18506 25848 18512 25900
rect 18564 25848 18570 25900
rect 21266 25848 21272 25900
rect 21324 25848 21330 25900
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 22020 25888 22048 25987
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 25130 25984 25136 26036
rect 25188 26024 25194 26036
rect 25866 26024 25872 26036
rect 25188 25996 25872 26024
rect 25188 25984 25194 25996
rect 25866 25984 25872 25996
rect 25924 26024 25930 26036
rect 26050 26024 26056 26036
rect 25924 25996 26056 26024
rect 25924 25984 25930 25996
rect 26050 25984 26056 25996
rect 26108 25984 26114 26036
rect 26234 25984 26240 26036
rect 26292 26024 26298 26036
rect 27341 26027 27399 26033
rect 27341 26024 27353 26027
rect 26292 25996 27353 26024
rect 26292 25984 26298 25996
rect 27341 25993 27353 25996
rect 27387 25993 27399 26027
rect 27341 25987 27399 25993
rect 28534 25984 28540 26036
rect 28592 26024 28598 26036
rect 28592 25996 30972 26024
rect 28592 25984 28598 25996
rect 24673 25959 24731 25965
rect 24673 25925 24685 25959
rect 24719 25956 24731 25959
rect 25222 25956 25228 25968
rect 24719 25928 25228 25956
rect 24719 25925 24731 25928
rect 24673 25919 24731 25925
rect 25222 25916 25228 25928
rect 25280 25916 25286 25968
rect 27154 25916 27160 25968
rect 27212 25956 27218 25968
rect 28353 25959 28411 25965
rect 28353 25956 28365 25959
rect 27212 25928 28365 25956
rect 27212 25916 27218 25928
rect 28353 25925 28365 25928
rect 28399 25956 28411 25959
rect 30006 25956 30012 25968
rect 28399 25928 30012 25956
rect 28399 25925 28411 25928
rect 28353 25919 28411 25925
rect 30006 25916 30012 25928
rect 30064 25916 30070 25968
rect 30101 25959 30159 25965
rect 30101 25925 30113 25959
rect 30147 25925 30159 25959
rect 30944 25956 30972 25996
rect 31018 25984 31024 26036
rect 31076 25984 31082 26036
rect 31294 26024 31300 26036
rect 31128 25996 31300 26024
rect 31128 25956 31156 25996
rect 31294 25984 31300 25996
rect 31352 26024 31358 26036
rect 31938 26024 31944 26036
rect 31352 25996 31944 26024
rect 31352 25984 31358 25996
rect 31938 25984 31944 25996
rect 31996 26024 32002 26036
rect 32306 26024 32312 26036
rect 31996 25996 32312 26024
rect 31996 25984 32002 25996
rect 32306 25984 32312 25996
rect 32364 25984 32370 26036
rect 32401 26027 32459 26033
rect 32401 25993 32413 26027
rect 32447 26024 32459 26027
rect 32490 26024 32496 26036
rect 32447 25996 32496 26024
rect 32447 25993 32459 25996
rect 32401 25987 32459 25993
rect 32490 25984 32496 25996
rect 32548 25984 32554 26036
rect 33226 25984 33232 26036
rect 33284 26024 33290 26036
rect 33321 26027 33379 26033
rect 33321 26024 33333 26027
rect 33284 25996 33333 26024
rect 33284 25984 33290 25996
rect 33321 25993 33333 25996
rect 33367 26024 33379 26027
rect 33686 26024 33692 26036
rect 33367 25996 33692 26024
rect 33367 25993 33379 25996
rect 33321 25987 33379 25993
rect 33686 25984 33692 25996
rect 33744 25984 33750 26036
rect 34054 25984 34060 26036
rect 34112 25984 34118 26036
rect 38102 26024 38108 26036
rect 35820 25996 38108 26024
rect 33042 25956 33048 25968
rect 30944 25928 31156 25956
rect 31220 25928 33048 25956
rect 30101 25919 30159 25925
rect 21499 25860 22048 25888
rect 22465 25891 22523 25897
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 22465 25857 22477 25891
rect 22511 25888 22523 25891
rect 22830 25888 22836 25900
rect 22511 25860 22836 25888
rect 22511 25857 22523 25860
rect 22465 25851 22523 25857
rect 22830 25848 22836 25860
rect 22888 25848 22894 25900
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 23474 25888 23480 25900
rect 23339 25860 23480 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25888 23627 25891
rect 23658 25888 23664 25900
rect 23615 25860 23664 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 23658 25848 23664 25860
rect 23716 25848 23722 25900
rect 24578 25848 24584 25900
rect 24636 25848 24642 25900
rect 24854 25848 24860 25900
rect 24912 25848 24918 25900
rect 25682 25848 25688 25900
rect 25740 25848 25746 25900
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25888 26203 25891
rect 27246 25888 27252 25900
rect 26191 25860 27252 25888
rect 26191 25857 26203 25860
rect 26145 25851 26203 25857
rect 27246 25848 27252 25860
rect 27304 25848 27310 25900
rect 27522 25848 27528 25900
rect 27580 25848 27586 25900
rect 27617 25891 27675 25897
rect 27617 25857 27629 25891
rect 27663 25857 27675 25891
rect 27617 25851 27675 25857
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25888 27951 25891
rect 27982 25888 27988 25900
rect 27939 25860 27988 25888
rect 27939 25857 27951 25860
rect 27893 25851 27951 25857
rect 13262 25780 13268 25832
rect 13320 25820 13326 25832
rect 13449 25823 13507 25829
rect 13449 25820 13461 25823
rect 13320 25792 13461 25820
rect 13320 25780 13326 25792
rect 13449 25789 13461 25792
rect 13495 25789 13507 25823
rect 13449 25783 13507 25789
rect 18598 25780 18604 25832
rect 18656 25780 18662 25832
rect 18877 25823 18935 25829
rect 18877 25789 18889 25823
rect 18923 25820 18935 25823
rect 19334 25820 19340 25832
rect 18923 25792 19340 25820
rect 18923 25789 18935 25792
rect 18877 25783 18935 25789
rect 19334 25780 19340 25792
rect 19392 25780 19398 25832
rect 20717 25823 20775 25829
rect 20717 25789 20729 25823
rect 20763 25820 20775 25823
rect 20990 25820 20996 25832
rect 20763 25792 20996 25820
rect 20763 25789 20775 25792
rect 20717 25783 20775 25789
rect 20990 25780 20996 25792
rect 21048 25780 21054 25832
rect 23382 25780 23388 25832
rect 23440 25780 23446 25832
rect 25041 25823 25099 25829
rect 25041 25789 25053 25823
rect 25087 25820 25099 25823
rect 25869 25823 25927 25829
rect 25869 25820 25881 25823
rect 25087 25792 25881 25820
rect 25087 25789 25099 25792
rect 25041 25783 25099 25789
rect 25869 25789 25881 25792
rect 25915 25789 25927 25823
rect 25869 25783 25927 25789
rect 25961 25823 26019 25829
rect 25961 25789 25973 25823
rect 26007 25789 26019 25823
rect 25961 25783 26019 25789
rect 25976 25752 26004 25783
rect 26050 25780 26056 25832
rect 26108 25780 26114 25832
rect 27632 25820 27660 25851
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 28166 25820 28172 25832
rect 27632 25792 28172 25820
rect 28166 25780 28172 25792
rect 28224 25820 28230 25832
rect 28442 25820 28448 25832
rect 28224 25792 28448 25820
rect 28224 25780 28230 25792
rect 28442 25780 28448 25792
rect 28500 25780 28506 25832
rect 30116 25820 30144 25919
rect 31220 25820 31248 25928
rect 33042 25916 33048 25928
rect 33100 25916 33106 25968
rect 34609 25959 34667 25965
rect 34609 25925 34621 25959
rect 34655 25956 34667 25959
rect 34698 25956 34704 25968
rect 34655 25928 34704 25956
rect 34655 25925 34667 25928
rect 34609 25919 34667 25925
rect 34698 25916 34704 25928
rect 34756 25916 34762 25968
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25888 31447 25891
rect 31754 25888 31760 25900
rect 31435 25860 31760 25888
rect 31435 25857 31447 25860
rect 31389 25851 31447 25857
rect 31754 25848 31760 25860
rect 31812 25848 31818 25900
rect 32398 25848 32404 25900
rect 32456 25848 32462 25900
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 30116 25792 31248 25820
rect 31478 25780 31484 25832
rect 31536 25780 31542 25832
rect 31573 25823 31631 25829
rect 31573 25789 31585 25823
rect 31619 25789 31631 25823
rect 32508 25820 32536 25851
rect 33134 25848 33140 25900
rect 33192 25848 33198 25900
rect 34149 25891 34207 25897
rect 34149 25857 34161 25891
rect 34195 25888 34207 25891
rect 35713 25891 35771 25897
rect 35713 25888 35725 25891
rect 34195 25860 35725 25888
rect 34195 25857 34207 25860
rect 34149 25851 34207 25857
rect 35713 25857 35725 25860
rect 35759 25888 35771 25891
rect 35820 25888 35848 25996
rect 38102 25984 38108 25996
rect 38160 25984 38166 26036
rect 38289 26027 38347 26033
rect 38289 25993 38301 26027
rect 38335 26024 38347 26027
rect 39206 26024 39212 26036
rect 38335 25996 39212 26024
rect 38335 25993 38347 25996
rect 38289 25987 38347 25993
rect 39206 25984 39212 25996
rect 39264 26024 39270 26036
rect 39390 26024 39396 26036
rect 39264 25996 39396 26024
rect 39264 25984 39270 25996
rect 39390 25984 39396 25996
rect 39448 26024 39454 26036
rect 40034 26024 40040 26036
rect 39448 25996 40040 26024
rect 39448 25984 39454 25996
rect 40034 25984 40040 25996
rect 40092 25984 40098 26036
rect 40310 25984 40316 26036
rect 40368 25984 40374 26036
rect 41230 25984 41236 26036
rect 41288 26024 41294 26036
rect 41288 25996 42932 26024
rect 41288 25984 41294 25996
rect 35986 25916 35992 25968
rect 36044 25916 36050 25968
rect 36446 25916 36452 25968
rect 36504 25956 36510 25968
rect 38749 25959 38807 25965
rect 38749 25956 38761 25959
rect 36504 25928 38761 25956
rect 36504 25916 36510 25928
rect 38749 25925 38761 25928
rect 38795 25925 38807 25959
rect 38749 25919 38807 25925
rect 39482 25916 39488 25968
rect 39540 25956 39546 25968
rect 41046 25956 41052 25968
rect 39540 25928 41052 25956
rect 39540 25916 39546 25928
rect 41046 25916 41052 25928
rect 41104 25916 41110 25968
rect 41690 25916 41696 25968
rect 41748 25916 41754 25968
rect 41898 25959 41956 25965
rect 41898 25925 41910 25959
rect 41944 25956 41956 25959
rect 41944 25928 42012 25956
rect 41944 25925 41956 25928
rect 41898 25919 41956 25925
rect 35759 25860 35848 25888
rect 36004 25888 36032 25916
rect 36173 25891 36231 25897
rect 36173 25888 36185 25891
rect 36004 25860 36185 25888
rect 35759 25857 35771 25860
rect 35713 25851 35771 25857
rect 36173 25857 36185 25860
rect 36219 25857 36231 25891
rect 36173 25851 36231 25857
rect 37366 25848 37372 25900
rect 37424 25888 37430 25900
rect 37645 25891 37703 25897
rect 37645 25888 37657 25891
rect 37424 25860 37657 25888
rect 37424 25848 37430 25860
rect 37645 25857 37657 25860
rect 37691 25857 37703 25891
rect 37645 25851 37703 25857
rect 37737 25891 37795 25897
rect 37737 25857 37749 25891
rect 37783 25888 37795 25891
rect 37826 25888 37832 25900
rect 37783 25860 37832 25888
rect 37783 25857 37795 25860
rect 37737 25851 37795 25857
rect 37826 25848 37832 25860
rect 37884 25848 37890 25900
rect 38286 25848 38292 25900
rect 38344 25888 38350 25900
rect 38933 25891 38991 25897
rect 38933 25888 38945 25891
rect 38344 25860 38945 25888
rect 38344 25848 38350 25860
rect 38933 25857 38945 25860
rect 38979 25857 38991 25891
rect 38933 25851 38991 25857
rect 39114 25848 39120 25900
rect 39172 25848 39178 25900
rect 39206 25848 39212 25900
rect 39264 25848 39270 25900
rect 40494 25848 40500 25900
rect 40552 25848 40558 25900
rect 31573 25783 31631 25789
rect 32416 25792 35388 25820
rect 27246 25752 27252 25764
rect 25976 25724 27252 25752
rect 27246 25712 27252 25724
rect 27304 25752 27310 25764
rect 27304 25724 27936 25752
rect 27304 25712 27310 25724
rect 14826 25644 14832 25696
rect 14884 25644 14890 25696
rect 15562 25644 15568 25696
rect 15620 25684 15626 25696
rect 15657 25687 15715 25693
rect 15657 25684 15669 25687
rect 15620 25656 15669 25684
rect 15620 25644 15626 25656
rect 15657 25653 15669 25656
rect 15703 25653 15715 25687
rect 15657 25647 15715 25653
rect 16022 25644 16028 25696
rect 16080 25684 16086 25696
rect 20073 25687 20131 25693
rect 20073 25684 20085 25687
rect 16080 25656 20085 25684
rect 16080 25644 16086 25656
rect 20073 25653 20085 25656
rect 20119 25653 20131 25687
rect 20073 25647 20131 25653
rect 21358 25644 21364 25696
rect 21416 25684 21422 25696
rect 21453 25687 21511 25693
rect 21453 25684 21465 25687
rect 21416 25656 21465 25684
rect 21416 25644 21422 25656
rect 21453 25653 21465 25656
rect 21499 25653 21511 25687
rect 21453 25647 21511 25653
rect 22370 25644 22376 25696
rect 22428 25684 22434 25696
rect 23014 25684 23020 25696
rect 22428 25656 23020 25684
rect 22428 25644 22434 25656
rect 23014 25644 23020 25656
rect 23072 25644 23078 25696
rect 23750 25644 23756 25696
rect 23808 25644 23814 25696
rect 26329 25687 26387 25693
rect 26329 25653 26341 25687
rect 26375 25684 26387 25687
rect 26970 25684 26976 25696
rect 26375 25656 26976 25684
rect 26375 25653 26387 25656
rect 26329 25647 26387 25653
rect 26970 25644 26976 25656
rect 27028 25644 27034 25696
rect 27706 25644 27712 25696
rect 27764 25684 27770 25696
rect 27801 25687 27859 25693
rect 27801 25684 27813 25687
rect 27764 25656 27813 25684
rect 27764 25644 27770 25656
rect 27801 25653 27813 25656
rect 27847 25653 27859 25687
rect 27908 25684 27936 25724
rect 31386 25712 31392 25764
rect 31444 25752 31450 25764
rect 31588 25752 31616 25783
rect 31444 25724 31616 25752
rect 31444 25712 31450 25724
rect 32416 25684 32444 25792
rect 34164 25764 34192 25792
rect 34146 25712 34152 25764
rect 34204 25712 34210 25764
rect 34606 25712 34612 25764
rect 34664 25712 34670 25764
rect 35360 25752 35388 25792
rect 35802 25780 35808 25832
rect 35860 25780 35866 25832
rect 35989 25823 36047 25829
rect 35989 25789 36001 25823
rect 36035 25820 36047 25823
rect 37461 25823 37519 25829
rect 37461 25820 37473 25823
rect 36035 25792 37473 25820
rect 36035 25789 36047 25792
rect 35989 25783 36047 25789
rect 37461 25789 37473 25792
rect 37507 25820 37519 25823
rect 37550 25820 37556 25832
rect 37507 25792 37556 25820
rect 37507 25789 37519 25792
rect 37461 25783 37519 25789
rect 37550 25780 37556 25792
rect 37608 25820 37614 25832
rect 41233 25823 41291 25829
rect 41233 25820 41245 25823
rect 37608 25792 41245 25820
rect 37608 25780 37614 25792
rect 41233 25789 41245 25792
rect 41279 25820 41291 25823
rect 41506 25820 41512 25832
rect 41279 25792 41512 25820
rect 41279 25789 41291 25792
rect 41233 25783 41291 25789
rect 41506 25780 41512 25792
rect 41564 25780 41570 25832
rect 36633 25755 36691 25761
rect 36633 25752 36645 25755
rect 35360 25724 36645 25752
rect 36633 25721 36645 25724
rect 36679 25752 36691 25755
rect 37826 25752 37832 25764
rect 36679 25724 37832 25752
rect 36679 25721 36691 25724
rect 36633 25715 36691 25721
rect 37826 25712 37832 25724
rect 37884 25712 37890 25764
rect 27908 25656 32444 25684
rect 27801 25647 27859 25653
rect 33410 25644 33416 25696
rect 33468 25684 33474 25696
rect 33873 25687 33931 25693
rect 33873 25684 33885 25687
rect 33468 25656 33885 25684
rect 33468 25644 33474 25656
rect 33873 25653 33885 25656
rect 33919 25653 33931 25687
rect 33873 25647 33931 25653
rect 35342 25644 35348 25696
rect 35400 25684 35406 25696
rect 35437 25687 35495 25693
rect 35437 25684 35449 25687
rect 35400 25656 35449 25684
rect 35400 25644 35406 25656
rect 35437 25653 35449 25656
rect 35483 25653 35495 25687
rect 35437 25647 35495 25653
rect 35897 25687 35955 25693
rect 35897 25653 35909 25687
rect 35943 25684 35955 25687
rect 36354 25684 36360 25696
rect 35943 25656 36360 25684
rect 35943 25653 35955 25656
rect 35897 25647 35955 25653
rect 36354 25644 36360 25656
rect 36412 25644 36418 25696
rect 37734 25644 37740 25696
rect 37792 25644 37798 25696
rect 37844 25684 37872 25712
rect 39482 25684 39488 25696
rect 37844 25656 39488 25684
rect 39482 25644 39488 25656
rect 39540 25684 39546 25696
rect 39669 25687 39727 25693
rect 39669 25684 39681 25687
rect 39540 25656 39681 25684
rect 39540 25644 39546 25656
rect 39669 25653 39681 25656
rect 39715 25653 39727 25687
rect 39669 25647 39727 25653
rect 41690 25644 41696 25696
rect 41748 25684 41754 25696
rect 41877 25687 41935 25693
rect 41877 25684 41889 25687
rect 41748 25656 41889 25684
rect 41748 25644 41754 25656
rect 41877 25653 41889 25656
rect 41923 25653 41935 25687
rect 41984 25684 42012 25928
rect 42518 25848 42524 25900
rect 42576 25888 42582 25900
rect 42904 25897 42932 25996
rect 42797 25891 42855 25897
rect 42797 25888 42809 25891
rect 42576 25860 42809 25888
rect 42576 25848 42582 25860
rect 42797 25857 42809 25860
rect 42843 25857 42855 25891
rect 42797 25851 42855 25857
rect 42889 25891 42947 25897
rect 42889 25857 42901 25891
rect 42935 25857 42947 25891
rect 42889 25851 42947 25857
rect 42061 25755 42119 25761
rect 42061 25721 42073 25755
rect 42107 25752 42119 25755
rect 42794 25752 42800 25764
rect 42107 25724 42800 25752
rect 42107 25721 42119 25724
rect 42061 25715 42119 25721
rect 42794 25712 42800 25724
rect 42852 25712 42858 25764
rect 42613 25687 42671 25693
rect 42613 25684 42625 25687
rect 41984 25656 42625 25684
rect 41877 25647 41935 25653
rect 42613 25653 42625 25656
rect 42659 25684 42671 25687
rect 42978 25684 42984 25696
rect 42659 25656 42984 25684
rect 42659 25653 42671 25656
rect 42613 25647 42671 25653
rect 42978 25644 42984 25656
rect 43036 25644 43042 25696
rect 1104 25594 43884 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 43884 25594
rect 1104 25520 43884 25542
rect 14274 25440 14280 25492
rect 14332 25440 14338 25492
rect 19426 25440 19432 25492
rect 19484 25480 19490 25492
rect 19613 25483 19671 25489
rect 19613 25480 19625 25483
rect 19484 25452 19625 25480
rect 19484 25440 19490 25452
rect 19613 25449 19625 25452
rect 19659 25449 19671 25483
rect 19613 25443 19671 25449
rect 22925 25483 22983 25489
rect 22925 25449 22937 25483
rect 22971 25480 22983 25483
rect 23014 25480 23020 25492
rect 22971 25452 23020 25480
rect 22971 25449 22983 25452
rect 22925 25443 22983 25449
rect 23014 25440 23020 25452
rect 23072 25440 23078 25492
rect 23109 25483 23167 25489
rect 23109 25449 23121 25483
rect 23155 25480 23167 25483
rect 23474 25480 23480 25492
rect 23155 25452 23480 25480
rect 23155 25449 23167 25452
rect 23109 25443 23167 25449
rect 23474 25440 23480 25452
rect 23532 25440 23538 25492
rect 23842 25440 23848 25492
rect 23900 25480 23906 25492
rect 24946 25480 24952 25492
rect 23900 25452 24952 25480
rect 23900 25440 23906 25452
rect 24946 25440 24952 25452
rect 25004 25440 25010 25492
rect 25222 25440 25228 25492
rect 25280 25440 25286 25492
rect 27338 25440 27344 25492
rect 27396 25480 27402 25492
rect 27525 25483 27583 25489
rect 27525 25480 27537 25483
rect 27396 25452 27537 25480
rect 27396 25440 27402 25452
rect 27525 25449 27537 25452
rect 27571 25449 27583 25483
rect 27525 25443 27583 25449
rect 27982 25440 27988 25492
rect 28040 25480 28046 25492
rect 29086 25480 29092 25492
rect 28040 25452 29092 25480
rect 28040 25440 28046 25452
rect 29086 25440 29092 25452
rect 29144 25480 29150 25492
rect 29144 25452 30236 25480
rect 29144 25440 29150 25452
rect 18138 25372 18144 25424
rect 18196 25412 18202 25424
rect 20165 25415 20223 25421
rect 20165 25412 20177 25415
rect 18196 25384 20177 25412
rect 18196 25372 18202 25384
rect 20165 25381 20177 25384
rect 20211 25412 20223 25415
rect 20898 25412 20904 25424
rect 20211 25384 20904 25412
rect 20211 25381 20223 25384
rect 20165 25375 20223 25381
rect 20898 25372 20904 25384
rect 20956 25372 20962 25424
rect 22066 25384 26004 25412
rect 15286 25304 15292 25356
rect 15344 25304 15350 25356
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 15562 25285 15568 25288
rect 15556 25276 15568 25285
rect 15523 25248 15568 25276
rect 15556 25239 15568 25248
rect 15562 25236 15568 25239
rect 15620 25236 15626 25288
rect 17678 25236 17684 25288
rect 17736 25236 17742 25288
rect 20806 25236 20812 25288
rect 20864 25276 20870 25288
rect 21085 25279 21143 25285
rect 21085 25276 21097 25279
rect 20864 25248 21097 25276
rect 20864 25236 20870 25248
rect 21085 25245 21097 25248
rect 21131 25276 21143 25279
rect 21450 25276 21456 25288
rect 21131 25248 21456 25276
rect 21131 25245 21143 25248
rect 21085 25239 21143 25245
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 22066 25276 22094 25384
rect 25976 25356 26004 25384
rect 26050 25372 26056 25424
rect 26108 25412 26114 25424
rect 29178 25412 29184 25424
rect 26108 25384 29184 25412
rect 26108 25372 26114 25384
rect 29178 25372 29184 25384
rect 29236 25372 29242 25424
rect 30208 25412 30236 25452
rect 30282 25440 30288 25492
rect 30340 25480 30346 25492
rect 30377 25483 30435 25489
rect 30377 25480 30389 25483
rect 30340 25452 30389 25480
rect 30340 25440 30346 25452
rect 30377 25449 30389 25452
rect 30423 25449 30435 25483
rect 30377 25443 30435 25449
rect 30742 25440 30748 25492
rect 30800 25480 30806 25492
rect 31205 25483 31263 25489
rect 31205 25480 31217 25483
rect 30800 25452 31217 25480
rect 30800 25440 30806 25452
rect 31205 25449 31217 25452
rect 31251 25449 31263 25483
rect 31205 25443 31263 25449
rect 31478 25440 31484 25492
rect 31536 25480 31542 25492
rect 32309 25483 32367 25489
rect 32309 25480 32321 25483
rect 31536 25452 32321 25480
rect 31536 25440 31542 25452
rect 32309 25449 32321 25452
rect 32355 25449 32367 25483
rect 32309 25443 32367 25449
rect 32398 25440 32404 25492
rect 32456 25480 32462 25492
rect 32766 25480 32772 25492
rect 32456 25452 32772 25480
rect 32456 25440 32462 25452
rect 32766 25440 32772 25452
rect 32824 25440 32830 25492
rect 34054 25440 34060 25492
rect 34112 25480 34118 25492
rect 34241 25483 34299 25489
rect 34241 25480 34253 25483
rect 34112 25452 34253 25480
rect 34112 25440 34118 25452
rect 34241 25449 34253 25452
rect 34287 25449 34299 25483
rect 34241 25443 34299 25449
rect 35713 25483 35771 25489
rect 35713 25449 35725 25483
rect 35759 25480 35771 25483
rect 37366 25480 37372 25492
rect 35759 25452 37372 25480
rect 35759 25449 35771 25452
rect 35713 25443 35771 25449
rect 37366 25440 37372 25452
rect 37424 25440 37430 25492
rect 39114 25440 39120 25492
rect 39172 25480 39178 25492
rect 42610 25480 42616 25492
rect 39172 25452 42616 25480
rect 39172 25440 39178 25452
rect 42610 25440 42616 25452
rect 42668 25480 42674 25492
rect 42981 25483 43039 25489
rect 42981 25480 42993 25483
rect 42668 25452 42993 25480
rect 42668 25440 42674 25452
rect 42981 25449 42993 25452
rect 43027 25449 43039 25483
rect 42981 25443 43039 25449
rect 31573 25415 31631 25421
rect 31573 25412 31585 25415
rect 29288 25384 30144 25412
rect 30208 25384 31585 25412
rect 23750 25304 23756 25356
rect 23808 25344 23814 25356
rect 24762 25344 24768 25356
rect 23808 25316 24768 25344
rect 23808 25304 23814 25316
rect 24762 25304 24768 25316
rect 24820 25344 24826 25356
rect 24946 25344 24952 25356
rect 24820 25316 24952 25344
rect 24820 25304 24826 25316
rect 24946 25304 24952 25316
rect 25004 25304 25010 25356
rect 25958 25304 25964 25356
rect 26016 25344 26022 25356
rect 26329 25347 26387 25353
rect 26329 25344 26341 25347
rect 26016 25316 26341 25344
rect 26016 25304 26022 25316
rect 26329 25313 26341 25316
rect 26375 25344 26387 25347
rect 29288 25344 29316 25384
rect 26375 25316 29316 25344
rect 26375 25313 26387 25316
rect 26329 25307 26387 25313
rect 29454 25304 29460 25356
rect 29512 25344 29518 25356
rect 30116 25344 30144 25384
rect 31573 25381 31585 25384
rect 31619 25412 31631 25415
rect 32674 25412 32680 25424
rect 31619 25384 32680 25412
rect 31619 25381 31631 25384
rect 31573 25375 31631 25381
rect 32674 25372 32680 25384
rect 32732 25372 32738 25424
rect 35526 25372 35532 25424
rect 35584 25412 35590 25424
rect 35894 25412 35900 25424
rect 35584 25384 35900 25412
rect 35584 25372 35590 25384
rect 35894 25372 35900 25384
rect 35952 25372 35958 25424
rect 39206 25412 39212 25424
rect 39040 25384 39212 25412
rect 30374 25344 30380 25356
rect 29512 25316 30052 25344
rect 30116 25316 30380 25344
rect 29512 25304 29518 25316
rect 21560 25248 22094 25276
rect 22281 25279 22339 25285
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 20901 25211 20959 25217
rect 20901 25208 20913 25211
rect 19484 25180 20913 25208
rect 19484 25168 19490 25180
rect 20901 25177 20913 25180
rect 20947 25208 20959 25211
rect 21560 25208 21588 25248
rect 22281 25245 22293 25279
rect 22327 25276 22339 25279
rect 22327 25248 23152 25276
rect 22327 25245 22339 25248
rect 22281 25239 22339 25245
rect 23124 25220 23152 25248
rect 23474 25236 23480 25288
rect 23532 25276 23538 25288
rect 23661 25279 23719 25285
rect 23661 25276 23673 25279
rect 23532 25248 23673 25276
rect 23532 25236 23538 25248
rect 23661 25245 23673 25248
rect 23707 25245 23719 25279
rect 23661 25239 23719 25245
rect 23842 25236 23848 25288
rect 23900 25236 23906 25288
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 25041 25279 25099 25285
rect 25041 25245 25053 25279
rect 25087 25276 25099 25279
rect 25130 25276 25136 25288
rect 25087 25248 25136 25276
rect 25087 25245 25099 25248
rect 25041 25239 25099 25245
rect 20947 25180 21588 25208
rect 21729 25211 21787 25217
rect 20947 25177 20959 25180
rect 20901 25171 20959 25177
rect 21729 25177 21741 25211
rect 21775 25208 21787 25211
rect 22738 25208 22744 25220
rect 21775 25180 22744 25208
rect 21775 25177 21787 25180
rect 21729 25171 21787 25177
rect 22738 25168 22744 25180
rect 22796 25208 22802 25220
rect 22796 25180 23060 25208
rect 22796 25168 22802 25180
rect 16669 25143 16727 25149
rect 16669 25109 16681 25143
rect 16715 25140 16727 25143
rect 17034 25140 17040 25152
rect 16715 25112 17040 25140
rect 16715 25109 16727 25112
rect 16669 25103 16727 25109
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 17494 25100 17500 25152
rect 17552 25100 17558 25152
rect 20714 25100 20720 25152
rect 20772 25100 20778 25152
rect 22830 25100 22836 25152
rect 22888 25140 22894 25152
rect 22941 25143 22999 25149
rect 22941 25140 22953 25143
rect 22888 25112 22953 25140
rect 22888 25100 22894 25112
rect 22941 25109 22953 25112
rect 22987 25109 22999 25143
rect 23032 25140 23060 25180
rect 23106 25168 23112 25220
rect 23164 25208 23170 25220
rect 23860 25208 23888 25236
rect 23164 25180 23888 25208
rect 23164 25168 23170 25180
rect 23934 25168 23940 25220
rect 23992 25208 23998 25220
rect 24029 25211 24087 25217
rect 24029 25208 24041 25211
rect 23992 25180 24041 25208
rect 23992 25168 23998 25180
rect 24029 25177 24041 25180
rect 24075 25208 24087 25211
rect 25056 25208 25084 25239
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 27614 25236 27620 25288
rect 27672 25276 27678 25288
rect 27709 25279 27767 25285
rect 27709 25276 27721 25279
rect 27672 25248 27721 25276
rect 27672 25236 27678 25248
rect 27709 25245 27721 25248
rect 27755 25245 27767 25279
rect 27709 25239 27767 25245
rect 27982 25236 27988 25288
rect 28040 25236 28046 25288
rect 28166 25236 28172 25288
rect 28224 25236 28230 25288
rect 28626 25236 28632 25288
rect 28684 25236 28690 25288
rect 29546 25236 29552 25288
rect 29604 25276 29610 25288
rect 30024 25285 30052 25316
rect 30374 25304 30380 25316
rect 30432 25304 30438 25356
rect 31294 25304 31300 25356
rect 31352 25344 31358 25356
rect 31481 25347 31539 25353
rect 31481 25344 31493 25347
rect 31352 25316 31493 25344
rect 31352 25304 31358 25316
rect 31481 25313 31493 25316
rect 31527 25313 31539 25347
rect 31481 25307 31539 25313
rect 34514 25304 34520 25356
rect 34572 25344 34578 25356
rect 35066 25344 35072 25356
rect 34572 25316 35072 25344
rect 34572 25304 34578 25316
rect 35066 25304 35072 25316
rect 35124 25344 35130 25356
rect 36357 25347 36415 25353
rect 36357 25344 36369 25347
rect 35124 25316 36369 25344
rect 35124 25304 35130 25316
rect 36357 25313 36369 25316
rect 36403 25313 36415 25347
rect 36357 25307 36415 25313
rect 36814 25304 36820 25356
rect 36872 25344 36878 25356
rect 36872 25316 38654 25344
rect 36872 25304 36878 25316
rect 29733 25279 29791 25285
rect 29733 25276 29745 25279
rect 29604 25248 29745 25276
rect 29604 25236 29610 25248
rect 29733 25245 29745 25248
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 30009 25279 30067 25285
rect 30009 25245 30021 25279
rect 30055 25245 30067 25279
rect 30009 25239 30067 25245
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25276 30251 25279
rect 30834 25276 30840 25288
rect 30239 25248 30840 25276
rect 30239 25245 30251 25248
rect 30193 25239 30251 25245
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 31386 25236 31392 25288
rect 31444 25236 31450 25288
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25276 31723 25279
rect 32306 25276 32312 25288
rect 31711 25248 32312 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 32306 25236 32312 25248
rect 32364 25236 32370 25288
rect 32398 25236 32404 25288
rect 32456 25236 32462 25288
rect 32674 25236 32680 25288
rect 32732 25276 32738 25288
rect 32861 25279 32919 25285
rect 32861 25276 32873 25279
rect 32732 25248 32873 25276
rect 32732 25236 32738 25248
rect 32861 25245 32873 25248
rect 32907 25245 32919 25279
rect 32861 25239 32919 25245
rect 33045 25279 33103 25285
rect 33045 25245 33057 25279
rect 33091 25276 33103 25279
rect 33502 25276 33508 25288
rect 33091 25248 33508 25276
rect 33091 25245 33103 25248
rect 33045 25239 33103 25245
rect 33502 25236 33508 25248
rect 33560 25276 33566 25288
rect 33778 25276 33784 25288
rect 33560 25248 33784 25276
rect 33560 25236 33566 25248
rect 33778 25236 33784 25248
rect 33836 25276 33842 25288
rect 34057 25279 34115 25285
rect 34057 25276 34069 25279
rect 33836 25248 34069 25276
rect 33836 25236 33842 25248
rect 34057 25245 34069 25248
rect 34103 25245 34115 25279
rect 34057 25239 34115 25245
rect 34974 25236 34980 25288
rect 35032 25236 35038 25288
rect 35161 25279 35219 25285
rect 35161 25245 35173 25279
rect 35207 25276 35219 25279
rect 35250 25276 35256 25288
rect 35207 25248 35256 25276
rect 35207 25245 35219 25248
rect 35161 25239 35219 25245
rect 35250 25236 35256 25248
rect 35308 25236 35314 25288
rect 35621 25279 35679 25285
rect 35621 25245 35633 25279
rect 35667 25245 35679 25279
rect 35621 25239 35679 25245
rect 35805 25279 35863 25285
rect 35805 25245 35817 25279
rect 35851 25276 35863 25279
rect 36262 25276 36268 25288
rect 35851 25248 36268 25276
rect 35851 25245 35863 25248
rect 35805 25239 35863 25245
rect 27430 25208 27436 25220
rect 24075 25180 25084 25208
rect 25148 25180 27436 25208
rect 24075 25177 24087 25180
rect 24029 25171 24087 25177
rect 25148 25140 25176 25180
rect 27430 25168 27436 25180
rect 27488 25208 27494 25220
rect 28994 25208 29000 25220
rect 27488 25180 29000 25208
rect 27488 25168 27494 25180
rect 28994 25168 29000 25180
rect 29052 25168 29058 25220
rect 29362 25168 29368 25220
rect 29420 25208 29426 25220
rect 29871 25211 29929 25217
rect 29871 25208 29883 25211
rect 29420 25180 29883 25208
rect 29420 25168 29426 25180
rect 29871 25177 29883 25180
rect 29917 25177 29929 25211
rect 29871 25171 29929 25177
rect 30101 25211 30159 25217
rect 30101 25177 30113 25211
rect 30147 25177 30159 25211
rect 31404 25208 31432 25236
rect 32953 25211 33011 25217
rect 32953 25208 32965 25211
rect 31404 25180 32965 25208
rect 30101 25171 30159 25177
rect 32953 25177 32965 25180
rect 32999 25177 33011 25211
rect 32953 25171 33011 25177
rect 23032 25112 25176 25140
rect 22941 25103 22999 25109
rect 25682 25100 25688 25152
rect 25740 25100 25746 25152
rect 26142 25100 26148 25152
rect 26200 25140 26206 25152
rect 26878 25140 26884 25152
rect 26200 25112 26884 25140
rect 26200 25100 26206 25112
rect 26878 25100 26884 25112
rect 26936 25100 26942 25152
rect 28810 25100 28816 25152
rect 28868 25100 28874 25152
rect 29638 25100 29644 25152
rect 29696 25140 29702 25152
rect 30116 25140 30144 25171
rect 33686 25168 33692 25220
rect 33744 25208 33750 25220
rect 33873 25211 33931 25217
rect 33873 25208 33885 25211
rect 33744 25180 33885 25208
rect 33744 25168 33750 25180
rect 33873 25177 33885 25180
rect 33919 25177 33931 25211
rect 33873 25171 33931 25177
rect 34606 25168 34612 25220
rect 34664 25208 34670 25220
rect 35342 25208 35348 25220
rect 34664 25180 35348 25208
rect 34664 25168 34670 25180
rect 35342 25168 35348 25180
rect 35400 25208 35406 25220
rect 35636 25208 35664 25239
rect 36262 25236 36268 25248
rect 36320 25236 36326 25288
rect 36630 25236 36636 25288
rect 36688 25276 36694 25288
rect 37277 25279 37335 25285
rect 37277 25276 37289 25279
rect 36688 25248 37289 25276
rect 36688 25236 36694 25248
rect 37277 25245 37289 25248
rect 37323 25245 37335 25279
rect 37277 25239 37335 25245
rect 37826 25236 37832 25288
rect 37884 25276 37890 25288
rect 38197 25279 38255 25285
rect 38197 25276 38209 25279
rect 37884 25248 38209 25276
rect 37884 25236 37890 25248
rect 38197 25245 38209 25248
rect 38243 25245 38255 25279
rect 38197 25239 38255 25245
rect 38378 25236 38384 25288
rect 38436 25236 38442 25288
rect 35400 25180 35664 25208
rect 35400 25168 35406 25180
rect 36722 25168 36728 25220
rect 36780 25208 36786 25220
rect 37093 25211 37151 25217
rect 37093 25208 37105 25211
rect 36780 25180 37105 25208
rect 36780 25168 36786 25180
rect 37093 25177 37105 25180
rect 37139 25177 37151 25211
rect 37093 25171 37151 25177
rect 37366 25168 37372 25220
rect 37424 25208 37430 25220
rect 38286 25208 38292 25220
rect 37424 25180 38292 25208
rect 37424 25168 37430 25180
rect 38286 25168 38292 25180
rect 38344 25168 38350 25220
rect 38626 25208 38654 25316
rect 39040 25270 39068 25384
rect 39206 25372 39212 25384
rect 39264 25372 39270 25424
rect 40034 25372 40040 25424
rect 40092 25412 40098 25424
rect 40092 25384 40264 25412
rect 40092 25372 40098 25384
rect 39117 25279 39175 25285
rect 39117 25270 39129 25279
rect 39040 25245 39129 25270
rect 39163 25245 39175 25279
rect 39040 25242 39175 25245
rect 39117 25239 39175 25242
rect 39206 25236 39212 25288
rect 39264 25236 39270 25288
rect 39298 25236 39304 25288
rect 39356 25276 39362 25288
rect 39393 25279 39451 25285
rect 39393 25276 39405 25279
rect 39356 25248 39405 25276
rect 39356 25236 39362 25248
rect 39393 25245 39405 25248
rect 39439 25245 39451 25279
rect 39393 25239 39451 25245
rect 39485 25279 39543 25285
rect 39485 25245 39497 25279
rect 39531 25276 39543 25279
rect 39531 25248 39712 25276
rect 39531 25245 39543 25248
rect 39485 25239 39543 25245
rect 39408 25208 39436 25239
rect 39574 25208 39580 25220
rect 38626 25180 39344 25208
rect 39408 25180 39580 25208
rect 29696 25112 30144 25140
rect 35069 25143 35127 25149
rect 29696 25100 29702 25112
rect 35069 25109 35081 25143
rect 35115 25140 35127 25143
rect 35434 25140 35440 25152
rect 35115 25112 35440 25140
rect 35115 25109 35127 25112
rect 35069 25103 35127 25109
rect 35434 25100 35440 25112
rect 35492 25100 35498 25152
rect 37458 25100 37464 25152
rect 37516 25100 37522 25152
rect 38933 25143 38991 25149
rect 38933 25109 38945 25143
rect 38979 25140 38991 25143
rect 39114 25140 39120 25152
rect 38979 25112 39120 25140
rect 38979 25109 38991 25112
rect 38933 25103 38991 25109
rect 39114 25100 39120 25112
rect 39172 25100 39178 25152
rect 39316 25140 39344 25180
rect 39574 25168 39580 25180
rect 39632 25168 39638 25220
rect 39684 25140 39712 25248
rect 40034 25236 40040 25288
rect 40092 25276 40098 25288
rect 40236 25285 40264 25384
rect 40494 25372 40500 25424
rect 40552 25412 40558 25424
rect 41325 25415 41383 25421
rect 41325 25412 41337 25415
rect 40552 25384 41337 25412
rect 40552 25372 40558 25384
rect 40221 25279 40279 25285
rect 40092 25248 40172 25276
rect 40092 25236 40098 25248
rect 40144 25208 40172 25248
rect 40221 25245 40233 25279
rect 40267 25245 40279 25279
rect 41156 25276 41184 25384
rect 41325 25381 41337 25384
rect 41371 25381 41383 25415
rect 41325 25375 41383 25381
rect 41874 25372 41880 25424
rect 41932 25412 41938 25424
rect 41932 25384 42865 25412
rect 41932 25372 41938 25384
rect 41230 25304 41236 25356
rect 41288 25344 41294 25356
rect 42837 25353 42865 25384
rect 42337 25347 42395 25353
rect 42337 25344 42349 25347
rect 41288 25316 42349 25344
rect 41288 25304 41294 25316
rect 42337 25313 42349 25316
rect 42383 25313 42395 25347
rect 42337 25307 42395 25313
rect 42822 25347 42880 25353
rect 42822 25313 42834 25347
rect 42868 25313 42880 25347
rect 42822 25307 42880 25313
rect 41156 25248 41414 25276
rect 40221 25239 40279 25245
rect 40865 25211 40923 25217
rect 40865 25208 40877 25211
rect 40144 25180 40877 25208
rect 40865 25177 40877 25180
rect 40911 25177 40923 25211
rect 40865 25171 40923 25177
rect 40129 25143 40187 25149
rect 40129 25140 40141 25143
rect 39316 25112 40141 25140
rect 40129 25109 40141 25112
rect 40175 25109 40187 25143
rect 41386 25140 41414 25248
rect 41506 25236 41512 25288
rect 41564 25276 41570 25288
rect 41693 25279 41751 25285
rect 41693 25276 41705 25279
rect 41564 25248 41705 25276
rect 41564 25236 41570 25248
rect 41693 25245 41705 25248
rect 41739 25245 41751 25279
rect 41693 25239 41751 25245
rect 41785 25279 41843 25285
rect 41785 25245 41797 25279
rect 41831 25276 41843 25279
rect 42058 25276 42064 25288
rect 41831 25248 42064 25276
rect 41831 25245 41843 25248
rect 41785 25239 41843 25245
rect 42058 25236 42064 25248
rect 42116 25236 42122 25288
rect 42426 25168 42432 25220
rect 42484 25208 42490 25220
rect 42484 25180 42748 25208
rect 42484 25168 42490 25180
rect 41966 25140 41972 25152
rect 41386 25112 41972 25140
rect 40129 25103 40187 25109
rect 41966 25100 41972 25112
rect 42024 25140 42030 25152
rect 42518 25140 42524 25152
rect 42024 25112 42524 25140
rect 42024 25100 42030 25112
rect 42518 25100 42524 25112
rect 42576 25140 42582 25152
rect 42720 25149 42748 25180
rect 42613 25143 42671 25149
rect 42613 25140 42625 25143
rect 42576 25112 42625 25140
rect 42576 25100 42582 25112
rect 42613 25109 42625 25112
rect 42659 25109 42671 25143
rect 42613 25103 42671 25109
rect 42705 25143 42763 25149
rect 42705 25109 42717 25143
rect 42751 25109 42763 25143
rect 42705 25103 42763 25109
rect 1104 25050 43884 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 43884 25050
rect 1104 24976 43884 24998
rect 15565 24939 15623 24945
rect 15565 24905 15577 24939
rect 15611 24936 15623 24939
rect 15838 24936 15844 24948
rect 15611 24908 15844 24936
rect 15611 24905 15623 24908
rect 15565 24899 15623 24905
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 19426 24896 19432 24948
rect 19484 24896 19490 24948
rect 20898 24896 20904 24948
rect 20956 24936 20962 24948
rect 21910 24936 21916 24948
rect 20956 24908 21916 24936
rect 20956 24896 20962 24908
rect 21910 24896 21916 24908
rect 21968 24936 21974 24948
rect 21968 24908 22140 24936
rect 21968 24896 21974 24908
rect 15933 24871 15991 24877
rect 15933 24837 15945 24871
rect 15979 24868 15991 24871
rect 17034 24868 17040 24880
rect 15979 24840 17040 24868
rect 15979 24837 15991 24840
rect 15933 24831 15991 24837
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 17494 24877 17500 24880
rect 17488 24868 17500 24877
rect 17455 24840 17500 24868
rect 17488 24831 17500 24840
rect 17494 24828 17500 24831
rect 17552 24828 17558 24880
rect 12894 24760 12900 24812
rect 12952 24760 12958 24812
rect 13797 24803 13855 24809
rect 13797 24800 13809 24803
rect 13096 24772 13809 24800
rect 13096 24673 13124 24772
rect 13797 24769 13809 24772
rect 13843 24769 13855 24803
rect 13797 24763 13855 24769
rect 16022 24760 16028 24812
rect 16080 24760 16086 24812
rect 18322 24800 18328 24812
rect 16224 24772 18328 24800
rect 13262 24692 13268 24744
rect 13320 24732 13326 24744
rect 16224 24741 16252 24772
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 19444 24800 19472 24896
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19444 24772 19993 24800
rect 19981 24769 19993 24772
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24800 20223 24803
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20211 24772 20637 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20625 24769 20637 24772
rect 20671 24800 20683 24803
rect 20806 24800 20812 24812
rect 20671 24772 20812 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 20806 24760 20812 24772
rect 20864 24760 20870 24812
rect 20898 24760 20904 24812
rect 20956 24760 20962 24812
rect 22112 24809 22140 24908
rect 24026 24896 24032 24948
rect 24084 24936 24090 24948
rect 24578 24936 24584 24948
rect 24084 24908 24584 24936
rect 24084 24896 24090 24908
rect 24578 24896 24584 24908
rect 24636 24896 24642 24948
rect 24765 24939 24823 24945
rect 24765 24905 24777 24939
rect 24811 24905 24823 24939
rect 24765 24899 24823 24905
rect 23474 24868 23480 24880
rect 23216 24840 23480 24868
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 23017 24803 23075 24809
rect 23017 24769 23029 24803
rect 23063 24800 23075 24803
rect 23106 24800 23112 24812
rect 23063 24772 23112 24800
rect 23063 24769 23075 24772
rect 23017 24763 23075 24769
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 13320 24704 13553 24732
rect 13320 24692 13326 24704
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 16209 24735 16267 24741
rect 16209 24701 16221 24735
rect 16255 24701 16267 24735
rect 16209 24695 16267 24701
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24701 17279 24735
rect 21358 24732 21364 24744
rect 17221 24695 17279 24701
rect 20824 24704 21364 24732
rect 13081 24667 13139 24673
rect 13081 24633 13093 24667
rect 13127 24633 13139 24667
rect 13081 24627 13139 24633
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 14921 24599 14979 24605
rect 14921 24596 14933 24599
rect 14700 24568 14933 24596
rect 14700 24556 14706 24568
rect 14921 24565 14933 24568
rect 14967 24565 14979 24599
rect 17236 24596 17264 24695
rect 20824 24608 20852 24704
rect 21358 24692 21364 24704
rect 21416 24732 21422 24744
rect 22020 24732 22048 24763
rect 21416 24704 22048 24732
rect 22112 24732 22140 24763
rect 23106 24760 23112 24772
rect 23164 24760 23170 24812
rect 23216 24809 23244 24840
rect 23474 24828 23480 24840
rect 23532 24828 23538 24880
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23201 24763 23259 24769
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24780 24800 24808 24899
rect 24946 24896 24952 24948
rect 25004 24896 25010 24948
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 31389 24939 31447 24945
rect 31389 24936 31401 24939
rect 27672 24908 31401 24936
rect 27672 24896 27678 24908
rect 31389 24905 31401 24908
rect 31435 24936 31447 24939
rect 31570 24936 31576 24948
rect 31435 24908 31576 24936
rect 31435 24905 31447 24908
rect 31389 24899 31447 24905
rect 31570 24896 31576 24908
rect 31628 24896 31634 24948
rect 31754 24936 31760 24948
rect 31726 24896 31760 24936
rect 31812 24896 31818 24948
rect 32306 24896 32312 24948
rect 32364 24896 32370 24948
rect 34698 24896 34704 24948
rect 34756 24936 34762 24948
rect 34756 24908 36768 24936
rect 34756 24896 34762 24908
rect 24964 24868 24992 24896
rect 24964 24840 25176 24868
rect 25148 24809 25176 24840
rect 28810 24828 28816 24880
rect 28868 24868 28874 24880
rect 28914 24871 28972 24877
rect 28914 24868 28926 24871
rect 28868 24840 28926 24868
rect 28868 24828 28874 24840
rect 28914 24837 28926 24840
rect 28960 24837 28972 24871
rect 28914 24831 28972 24837
rect 29086 24828 29092 24880
rect 29144 24868 29150 24880
rect 29144 24840 30052 24868
rect 29144 24828 29150 24840
rect 23983 24772 24808 24800
rect 24949 24803 25007 24809
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 25133 24803 25191 24809
rect 25133 24769 25145 24803
rect 25179 24769 25191 24803
rect 25133 24763 25191 24769
rect 26513 24803 26571 24809
rect 26513 24769 26525 24803
rect 26559 24800 26571 24803
rect 26694 24800 26700 24812
rect 26559 24772 26700 24800
rect 26559 24769 26571 24772
rect 26513 24763 26571 24769
rect 23566 24732 23572 24744
rect 22112 24704 23572 24732
rect 21416 24692 21422 24704
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 23842 24692 23848 24744
rect 23900 24692 23906 24744
rect 24210 24692 24216 24744
rect 24268 24692 24274 24744
rect 24305 24735 24363 24741
rect 24305 24701 24317 24735
rect 24351 24701 24363 24735
rect 24305 24695 24363 24701
rect 23109 24667 23167 24673
rect 23109 24633 23121 24667
rect 23155 24664 23167 24667
rect 24026 24664 24032 24676
rect 23155 24636 24032 24664
rect 23155 24633 23167 24636
rect 23109 24627 23167 24633
rect 24026 24624 24032 24636
rect 24084 24624 24090 24676
rect 24320 24664 24348 24695
rect 24578 24692 24584 24744
rect 24636 24732 24642 24744
rect 24964 24732 24992 24763
rect 26694 24760 26700 24772
rect 26752 24800 26758 24812
rect 27154 24800 27160 24812
rect 26752 24772 27160 24800
rect 26752 24760 26758 24772
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 27246 24760 27252 24812
rect 27304 24760 27310 24812
rect 28166 24760 28172 24812
rect 28224 24800 28230 24812
rect 29181 24803 29239 24809
rect 28224 24772 29132 24800
rect 28224 24760 28230 24772
rect 24636 24704 24992 24732
rect 25041 24735 25099 24741
rect 24636 24692 24642 24704
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 25087 24704 25176 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 25148 24676 25176 24704
rect 25222 24692 25228 24744
rect 25280 24692 25286 24744
rect 29104 24732 29132 24772
rect 29181 24769 29193 24803
rect 29227 24800 29239 24803
rect 29362 24800 29368 24812
rect 29227 24772 29368 24800
rect 29227 24769 29239 24772
rect 29181 24763 29239 24769
rect 29362 24760 29368 24772
rect 29420 24800 29426 24812
rect 29730 24800 29736 24812
rect 29420 24772 29736 24800
rect 29420 24760 29426 24772
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 29914 24760 29920 24812
rect 29972 24760 29978 24812
rect 30024 24809 30052 24840
rect 30374 24828 30380 24880
rect 30432 24868 30438 24880
rect 31726 24868 31754 24896
rect 35894 24868 35900 24880
rect 30432 24840 31754 24868
rect 32876 24840 35900 24868
rect 30432 24828 30438 24840
rect 30009 24803 30067 24809
rect 30009 24769 30021 24803
rect 30055 24769 30067 24803
rect 30009 24763 30067 24769
rect 30098 24760 30104 24812
rect 30156 24800 30162 24812
rect 30285 24803 30343 24809
rect 30285 24800 30297 24803
rect 30156 24772 30297 24800
rect 30156 24760 30162 24772
rect 30285 24769 30297 24772
rect 30331 24769 30343 24803
rect 30285 24763 30343 24769
rect 30834 24760 30840 24812
rect 30892 24760 30898 24812
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31386 24800 31392 24812
rect 30975 24772 31392 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 31386 24760 31392 24772
rect 31444 24760 31450 24812
rect 32122 24760 32128 24812
rect 32180 24800 32186 24812
rect 32398 24800 32404 24812
rect 32180 24772 32404 24800
rect 32180 24760 32186 24772
rect 32398 24760 32404 24772
rect 32456 24800 32462 24812
rect 32493 24803 32551 24809
rect 32493 24800 32505 24803
rect 32456 24772 32505 24800
rect 32456 24760 32462 24772
rect 32493 24769 32505 24772
rect 32539 24769 32551 24803
rect 32769 24803 32827 24809
rect 32769 24800 32781 24803
rect 32493 24763 32551 24769
rect 32600 24772 32781 24800
rect 30852 24732 30880 24760
rect 32600 24732 32628 24772
rect 32769 24769 32781 24772
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 29104 24704 32628 24732
rect 32674 24692 32680 24744
rect 32732 24732 32738 24744
rect 32876 24732 32904 24840
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24800 33011 24803
rect 33689 24803 33747 24809
rect 32999 24772 33548 24800
rect 32999 24769 33011 24772
rect 32953 24763 33011 24769
rect 32732 24704 32904 24732
rect 32732 24692 32738 24704
rect 24320 24636 24992 24664
rect 18414 24596 18420 24608
rect 17236 24568 18420 24596
rect 14921 24559 14979 24565
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 18598 24556 18604 24608
rect 18656 24556 18662 24608
rect 20070 24556 20076 24608
rect 20128 24556 20134 24608
rect 20717 24599 20775 24605
rect 20717 24565 20729 24599
rect 20763 24596 20775 24599
rect 20806 24596 20812 24608
rect 20763 24568 20812 24596
rect 20763 24565 20775 24568
rect 20717 24559 20775 24565
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 21082 24556 21088 24608
rect 21140 24556 21146 24608
rect 21450 24556 21456 24608
rect 21508 24596 21514 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21508 24568 22017 24596
rect 21508 24556 21514 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22005 24559 22063 24565
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 23658 24556 23664 24608
rect 23716 24556 23722 24608
rect 24210 24556 24216 24608
rect 24268 24596 24274 24608
rect 24854 24596 24860 24608
rect 24268 24568 24860 24596
rect 24268 24556 24274 24568
rect 24854 24556 24860 24568
rect 24912 24556 24918 24608
rect 24964 24596 24992 24636
rect 25130 24624 25136 24676
rect 25188 24624 25194 24676
rect 27801 24667 27859 24673
rect 27801 24633 27813 24667
rect 27847 24664 27859 24667
rect 28074 24664 28080 24676
rect 27847 24636 28080 24664
rect 27847 24633 27859 24636
rect 27801 24627 27859 24633
rect 28074 24624 28080 24636
rect 28132 24624 28138 24676
rect 29454 24624 29460 24676
rect 29512 24664 29518 24676
rect 30837 24667 30895 24673
rect 30837 24664 30849 24667
rect 29512 24636 30849 24664
rect 29512 24624 29518 24636
rect 30837 24633 30849 24636
rect 30883 24633 30895 24667
rect 30837 24627 30895 24633
rect 32582 24624 32588 24676
rect 32640 24624 32646 24676
rect 33520 24664 33548 24772
rect 33689 24769 33701 24803
rect 33735 24800 33747 24803
rect 33778 24800 33784 24812
rect 33735 24772 33784 24800
rect 33735 24769 33747 24772
rect 33689 24763 33747 24769
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 33873 24803 33931 24809
rect 33873 24769 33885 24803
rect 33919 24769 33931 24803
rect 33873 24763 33931 24769
rect 33594 24692 33600 24744
rect 33652 24732 33658 24744
rect 33888 24732 33916 24763
rect 34514 24760 34520 24812
rect 34572 24760 34578 24812
rect 34716 24809 34744 24840
rect 35894 24828 35900 24840
rect 35952 24828 35958 24880
rect 35989 24871 36047 24877
rect 35989 24837 36001 24871
rect 36035 24868 36047 24871
rect 36740 24868 36768 24908
rect 37826 24896 37832 24948
rect 37884 24936 37890 24948
rect 38473 24939 38531 24945
rect 38473 24936 38485 24939
rect 37884 24908 38485 24936
rect 37884 24896 37890 24908
rect 38473 24905 38485 24908
rect 38519 24905 38531 24939
rect 38473 24899 38531 24905
rect 36035 24840 36676 24868
rect 36740 24840 40264 24868
rect 36035 24837 36047 24840
rect 35989 24831 36047 24837
rect 36648 24812 36676 24840
rect 34701 24803 34759 24809
rect 34701 24769 34713 24803
rect 34747 24769 34759 24803
rect 34701 24763 34759 24769
rect 34974 24760 34980 24812
rect 35032 24800 35038 24812
rect 35342 24800 35348 24812
rect 35032 24772 35348 24800
rect 35032 24760 35038 24772
rect 35342 24760 35348 24772
rect 35400 24800 35406 24812
rect 35618 24800 35624 24812
rect 35400 24772 35624 24800
rect 35400 24760 35406 24772
rect 35618 24760 35624 24772
rect 35676 24800 35682 24812
rect 35713 24803 35771 24809
rect 35713 24800 35725 24803
rect 35676 24772 35725 24800
rect 35676 24760 35682 24772
rect 35713 24769 35725 24772
rect 35759 24769 35771 24803
rect 35713 24763 35771 24769
rect 36449 24803 36507 24809
rect 36449 24769 36461 24803
rect 36495 24800 36507 24803
rect 36538 24800 36544 24812
rect 36495 24772 36544 24800
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 36630 24760 36636 24812
rect 36688 24760 36694 24812
rect 36725 24803 36783 24809
rect 36725 24769 36737 24803
rect 36771 24800 36783 24803
rect 37734 24800 37740 24812
rect 36771 24772 37740 24800
rect 36771 24769 36783 24772
rect 36725 24763 36783 24769
rect 37734 24760 37740 24772
rect 37792 24760 37798 24812
rect 39301 24803 39359 24809
rect 39301 24769 39313 24803
rect 39347 24800 39359 24803
rect 40034 24800 40040 24812
rect 39347 24772 40040 24800
rect 39347 24769 39359 24772
rect 39301 24763 39359 24769
rect 33652 24704 35296 24732
rect 33652 24692 33658 24704
rect 35268 24676 35296 24704
rect 35986 24692 35992 24744
rect 36044 24692 36050 24744
rect 37090 24692 37096 24744
rect 37148 24732 37154 24744
rect 37461 24735 37519 24741
rect 37461 24732 37473 24735
rect 37148 24704 37473 24732
rect 37148 24692 37154 24704
rect 37461 24701 37473 24704
rect 37507 24701 37519 24735
rect 39316 24732 39344 24763
rect 40034 24760 40040 24772
rect 40092 24760 40098 24812
rect 40126 24760 40132 24812
rect 40184 24760 40190 24812
rect 37461 24695 37519 24701
rect 37568 24704 39344 24732
rect 39393 24735 39451 24741
rect 34422 24664 34428 24676
rect 33520 24636 34428 24664
rect 34422 24624 34428 24636
rect 34480 24624 34486 24676
rect 35066 24624 35072 24676
rect 35124 24664 35130 24676
rect 35161 24667 35219 24673
rect 35161 24664 35173 24667
rect 35124 24636 35173 24664
rect 35124 24624 35130 24636
rect 35161 24633 35173 24636
rect 35207 24633 35219 24667
rect 35161 24627 35219 24633
rect 35250 24624 35256 24676
rect 35308 24664 35314 24676
rect 35618 24664 35624 24676
rect 35308 24636 35624 24664
rect 35308 24624 35314 24636
rect 35618 24624 35624 24636
rect 35676 24664 35682 24676
rect 37568 24664 37596 24704
rect 39393 24701 39405 24735
rect 39439 24701 39451 24735
rect 39393 24695 39451 24701
rect 35676 24636 37596 24664
rect 35676 24624 35682 24636
rect 37734 24624 37740 24676
rect 37792 24624 37798 24676
rect 37826 24624 37832 24676
rect 37884 24664 37890 24676
rect 37921 24667 37979 24673
rect 37921 24664 37933 24667
rect 37884 24636 37933 24664
rect 37884 24624 37890 24636
rect 37921 24633 37933 24636
rect 37967 24633 37979 24667
rect 37921 24627 37979 24633
rect 38010 24624 38016 24676
rect 38068 24664 38074 24676
rect 39408 24664 39436 24695
rect 39482 24692 39488 24744
rect 39540 24692 39546 24744
rect 39577 24735 39635 24741
rect 39577 24701 39589 24735
rect 39623 24732 39635 24735
rect 39666 24732 39672 24744
rect 39623 24704 39672 24732
rect 39623 24701 39635 24704
rect 39577 24695 39635 24701
rect 39666 24692 39672 24704
rect 39724 24692 39730 24744
rect 40236 24732 40264 24840
rect 41782 24828 41788 24880
rect 41840 24868 41846 24880
rect 42751 24871 42809 24877
rect 42751 24868 42763 24871
rect 41840 24840 42763 24868
rect 41840 24828 41846 24840
rect 42751 24837 42763 24840
rect 42797 24837 42809 24871
rect 42751 24831 42809 24837
rect 42978 24828 42984 24880
rect 43036 24828 43042 24880
rect 40310 24760 40316 24812
rect 40368 24760 40374 24812
rect 40494 24760 40500 24812
rect 40552 24800 40558 24812
rect 40773 24803 40831 24809
rect 40773 24800 40785 24803
rect 40552 24772 40785 24800
rect 40552 24760 40558 24772
rect 40773 24769 40785 24772
rect 40819 24769 40831 24803
rect 40773 24763 40831 24769
rect 40865 24803 40923 24809
rect 40865 24769 40877 24803
rect 40911 24800 40923 24803
rect 41138 24800 41144 24812
rect 40911 24772 41144 24800
rect 40911 24769 40923 24772
rect 40865 24763 40923 24769
rect 41138 24760 41144 24772
rect 41196 24760 41202 24812
rect 41693 24803 41751 24809
rect 41693 24769 41705 24803
rect 41739 24800 41751 24803
rect 41739 24772 41920 24800
rect 41739 24769 41751 24772
rect 41693 24763 41751 24769
rect 40236 24704 40448 24732
rect 38068 24636 39436 24664
rect 38068 24624 38074 24636
rect 25777 24599 25835 24605
rect 25777 24596 25789 24599
rect 24964 24568 25789 24596
rect 25777 24565 25789 24568
rect 25823 24596 25835 24599
rect 28258 24596 28264 24608
rect 25823 24568 28264 24596
rect 25823 24565 25835 24568
rect 25777 24559 25835 24565
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 29730 24556 29736 24608
rect 29788 24556 29794 24608
rect 30193 24599 30251 24605
rect 30193 24565 30205 24599
rect 30239 24596 30251 24599
rect 30742 24596 30748 24608
rect 30239 24568 30748 24596
rect 30239 24565 30251 24568
rect 30193 24559 30251 24565
rect 30742 24556 30748 24568
rect 30800 24556 30806 24608
rect 31662 24556 31668 24608
rect 31720 24596 31726 24608
rect 33873 24599 33931 24605
rect 33873 24596 33885 24599
rect 31720 24568 33885 24596
rect 31720 24556 31726 24568
rect 33873 24565 33885 24568
rect 33919 24596 33931 24599
rect 34514 24596 34520 24608
rect 33919 24568 34520 24596
rect 33919 24565 33931 24568
rect 33873 24559 33931 24565
rect 34514 24556 34520 24568
rect 34572 24556 34578 24608
rect 34698 24556 34704 24608
rect 34756 24556 34762 24608
rect 35710 24556 35716 24608
rect 35768 24596 35774 24608
rect 35805 24599 35863 24605
rect 35805 24596 35817 24599
rect 35768 24568 35817 24596
rect 35768 24556 35774 24568
rect 35805 24565 35817 24568
rect 35851 24565 35863 24599
rect 35805 24559 35863 24565
rect 36446 24556 36452 24608
rect 36504 24556 36510 24608
rect 36906 24556 36912 24608
rect 36964 24556 36970 24608
rect 39022 24556 39028 24608
rect 39080 24596 39086 24608
rect 39117 24599 39175 24605
rect 39117 24596 39129 24599
rect 39080 24568 39129 24596
rect 39080 24556 39086 24568
rect 39117 24565 39129 24568
rect 39163 24565 39175 24599
rect 39117 24559 39175 24565
rect 39482 24556 39488 24608
rect 39540 24596 39546 24608
rect 40313 24599 40371 24605
rect 40313 24596 40325 24599
rect 39540 24568 40325 24596
rect 39540 24556 39546 24568
rect 40313 24565 40325 24568
rect 40359 24565 40371 24599
rect 40420 24596 40448 24704
rect 41230 24692 41236 24744
rect 41288 24732 41294 24744
rect 41785 24735 41843 24741
rect 41785 24732 41797 24735
rect 41288 24704 41797 24732
rect 41288 24692 41294 24704
rect 41785 24701 41797 24704
rect 41831 24701 41843 24735
rect 41892 24732 41920 24772
rect 41966 24760 41972 24812
rect 42024 24760 42030 24812
rect 42610 24760 42616 24812
rect 42668 24760 42674 24812
rect 42886 24760 42892 24812
rect 42944 24760 42950 24812
rect 43070 24760 43076 24812
rect 43128 24760 43134 24812
rect 42426 24732 42432 24744
rect 41892 24704 42432 24732
rect 41785 24695 41843 24701
rect 42426 24692 42432 24704
rect 42484 24692 42490 24744
rect 40494 24624 40500 24676
rect 40552 24664 40558 24676
rect 41509 24667 41567 24673
rect 41509 24664 41521 24667
rect 40552 24636 41521 24664
rect 40552 24624 40558 24636
rect 41509 24633 41521 24636
rect 41555 24633 41567 24667
rect 43257 24667 43315 24673
rect 43257 24664 43269 24667
rect 41509 24627 41567 24633
rect 41616 24636 43269 24664
rect 41616 24596 41644 24636
rect 43257 24633 43269 24636
rect 43303 24633 43315 24667
rect 43257 24627 43315 24633
rect 40420 24568 41644 24596
rect 40313 24559 40371 24565
rect 41874 24556 41880 24608
rect 41932 24556 41938 24608
rect 1104 24506 43884 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 43884 24506
rect 1104 24432 43884 24454
rect 12894 24352 12900 24404
rect 12952 24392 12958 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 12952 24364 14289 24392
rect 12952 24352 12958 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 17678 24352 17684 24404
rect 17736 24352 17742 24404
rect 20346 24352 20352 24404
rect 20404 24392 20410 24404
rect 20404 24364 21680 24392
rect 20404 24352 20410 24364
rect 19797 24327 19855 24333
rect 19797 24293 19809 24327
rect 19843 24324 19855 24327
rect 20622 24324 20628 24336
rect 19843 24296 20628 24324
rect 19843 24293 19855 24296
rect 19797 24287 19855 24293
rect 20622 24284 20628 24296
rect 20680 24284 20686 24336
rect 14921 24259 14979 24265
rect 14921 24225 14933 24259
rect 14967 24256 14979 24259
rect 15102 24256 15108 24268
rect 14967 24228 15108 24256
rect 14967 24225 14979 24228
rect 14921 24219 14979 24225
rect 15102 24216 15108 24228
rect 15160 24256 15166 24268
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 15160 24228 15485 24256
rect 15160 24216 15166 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 15473 24219 15531 24225
rect 18322 24216 18328 24268
rect 18380 24216 18386 24268
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24256 20315 24259
rect 21545 24259 21603 24265
rect 21545 24256 21557 24259
rect 20303 24228 21557 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 21545 24225 21557 24228
rect 21591 24225 21603 24259
rect 21652 24256 21680 24364
rect 21726 24352 21732 24404
rect 21784 24392 21790 24404
rect 23658 24392 23664 24404
rect 21784 24364 23664 24392
rect 21784 24352 21790 24364
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 23753 24395 23811 24401
rect 23753 24361 23765 24395
rect 23799 24392 23811 24395
rect 23842 24392 23848 24404
rect 23799 24364 23848 24392
rect 23799 24361 23811 24364
rect 23753 24355 23811 24361
rect 23842 24352 23848 24364
rect 23900 24352 23906 24404
rect 24762 24352 24768 24404
rect 24820 24352 24826 24404
rect 24854 24352 24860 24404
rect 24912 24392 24918 24404
rect 25685 24395 25743 24401
rect 25685 24392 25697 24395
rect 24912 24364 25697 24392
rect 24912 24352 24918 24364
rect 25685 24361 25697 24364
rect 25731 24361 25743 24395
rect 25685 24355 25743 24361
rect 28445 24395 28503 24401
rect 28445 24361 28457 24395
rect 28491 24392 28503 24395
rect 28626 24392 28632 24404
rect 28491 24364 28632 24392
rect 28491 24361 28503 24364
rect 28445 24355 28503 24361
rect 28626 24352 28632 24364
rect 28684 24352 28690 24404
rect 29914 24352 29920 24404
rect 29972 24392 29978 24404
rect 30929 24395 30987 24401
rect 30929 24392 30941 24395
rect 29972 24364 30941 24392
rect 29972 24352 29978 24364
rect 30929 24361 30941 24364
rect 30975 24361 30987 24395
rect 30929 24355 30987 24361
rect 32953 24395 33011 24401
rect 32953 24361 32965 24395
rect 32999 24392 33011 24395
rect 33042 24392 33048 24404
rect 32999 24364 33048 24392
rect 32999 24361 33011 24364
rect 32953 24355 33011 24361
rect 33042 24352 33048 24364
rect 33100 24352 33106 24404
rect 35069 24395 35127 24401
rect 35069 24361 35081 24395
rect 35115 24392 35127 24395
rect 35342 24392 35348 24404
rect 35115 24364 35348 24392
rect 35115 24361 35127 24364
rect 35069 24355 35127 24361
rect 35342 24352 35348 24364
rect 35400 24392 35406 24404
rect 35802 24392 35808 24404
rect 35400 24364 35808 24392
rect 35400 24352 35406 24364
rect 35802 24352 35808 24364
rect 35860 24352 35866 24404
rect 35894 24352 35900 24404
rect 35952 24392 35958 24404
rect 36538 24392 36544 24404
rect 35952 24364 36544 24392
rect 35952 24352 35958 24364
rect 36538 24352 36544 24364
rect 36596 24352 36602 24404
rect 36725 24395 36783 24401
rect 36725 24361 36737 24395
rect 36771 24392 36783 24395
rect 36771 24364 37320 24392
rect 36771 24361 36783 24364
rect 36725 24355 36783 24361
rect 21818 24284 21824 24336
rect 21876 24324 21882 24336
rect 22554 24324 22560 24336
rect 21876 24296 22560 24324
rect 21876 24284 21882 24296
rect 22554 24284 22560 24296
rect 22612 24284 22618 24336
rect 23106 24284 23112 24336
rect 23164 24284 23170 24336
rect 32490 24324 32496 24336
rect 26804 24296 32496 24324
rect 21652 24228 26740 24256
rect 21545 24219 21603 24225
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 16022 24188 16028 24200
rect 14783 24160 16028 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 19521 24191 19579 24197
rect 19521 24157 19533 24191
rect 19567 24188 19579 24191
rect 20070 24188 20076 24200
rect 19567 24160 20076 24188
rect 19567 24157 19579 24160
rect 19521 24151 19579 24157
rect 20070 24148 20076 24160
rect 20128 24188 20134 24200
rect 20272 24188 20300 24219
rect 20128 24160 20300 24188
rect 20625 24191 20683 24197
rect 20128 24148 20134 24160
rect 20625 24157 20637 24191
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 18049 24123 18107 24129
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 18598 24120 18604 24132
rect 18095 24092 18604 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18598 24080 18604 24092
rect 18656 24080 18662 24132
rect 19797 24123 19855 24129
rect 19797 24089 19809 24123
rect 19843 24120 19855 24123
rect 20640 24120 20668 24151
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 21637 24191 21695 24197
rect 21637 24188 21649 24191
rect 20772 24160 21649 24188
rect 20772 24148 20778 24160
rect 21637 24157 21649 24160
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 21729 24191 21787 24197
rect 21729 24157 21741 24191
rect 21775 24157 21787 24191
rect 21729 24151 21787 24157
rect 21082 24120 21088 24132
rect 19843 24092 21088 24120
rect 19843 24089 19855 24092
rect 19797 24083 19855 24089
rect 21082 24080 21088 24092
rect 21140 24120 21146 24132
rect 21744 24120 21772 24151
rect 21818 24148 21824 24200
rect 21876 24148 21882 24200
rect 22373 24191 22431 24197
rect 22373 24188 22385 24191
rect 22066 24160 22385 24188
rect 22066 24120 22094 24160
rect 22373 24157 22385 24160
rect 22419 24157 22431 24191
rect 22373 24151 22431 24157
rect 22554 24148 22560 24200
rect 22612 24148 22618 24200
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 24026 24148 24032 24200
rect 24084 24148 24090 24200
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 24544 24160 24593 24188
rect 24544 24148 24550 24160
rect 24581 24157 24593 24160
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 24949 24191 25007 24197
rect 24949 24157 24961 24191
rect 24995 24188 25007 24191
rect 25222 24188 25228 24200
rect 24995 24160 25228 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25222 24148 25228 24160
rect 25280 24188 25286 24200
rect 25869 24191 25927 24197
rect 25869 24188 25881 24191
rect 25280 24160 25881 24188
rect 25280 24148 25286 24160
rect 25869 24157 25881 24160
rect 25915 24157 25927 24191
rect 25869 24151 25927 24157
rect 21140 24092 22094 24120
rect 22572 24120 22600 24148
rect 22922 24120 22928 24132
rect 22572 24092 22928 24120
rect 21140 24080 21146 24092
rect 22922 24080 22928 24092
rect 22980 24120 22986 24132
rect 24210 24120 24216 24132
rect 22980 24092 24216 24120
rect 22980 24080 22986 24092
rect 24210 24080 24216 24092
rect 24268 24080 24274 24132
rect 25884 24120 25912 24151
rect 26602 24148 26608 24200
rect 26660 24148 26666 24200
rect 26712 24197 26740 24228
rect 26698 24191 26756 24197
rect 26698 24157 26710 24191
rect 26744 24157 26756 24191
rect 26698 24151 26756 24157
rect 26804 24120 26832 24296
rect 32490 24284 32496 24296
rect 32548 24284 32554 24336
rect 33502 24284 33508 24336
rect 33560 24324 33566 24336
rect 35710 24324 35716 24336
rect 33560 24296 35716 24324
rect 33560 24284 33566 24296
rect 27801 24259 27859 24265
rect 27801 24256 27813 24259
rect 26896 24228 27813 24256
rect 26896 24197 26924 24228
rect 27801 24225 27813 24228
rect 27847 24225 27859 24259
rect 28166 24256 28172 24268
rect 27801 24219 27859 24225
rect 27908 24228 28172 24256
rect 27908 24200 27936 24228
rect 28166 24216 28172 24228
rect 28224 24216 28230 24268
rect 29089 24259 29147 24265
rect 29089 24225 29101 24259
rect 29135 24256 29147 24259
rect 29730 24256 29736 24268
rect 29135 24228 29736 24256
rect 29135 24225 29147 24228
rect 29089 24219 29147 24225
rect 29730 24216 29736 24228
rect 29788 24216 29794 24268
rect 30285 24259 30343 24265
rect 30285 24256 30297 24259
rect 30024 24228 30297 24256
rect 27154 24197 27160 24200
rect 26881 24191 26939 24197
rect 26881 24157 26893 24191
rect 26927 24157 26939 24191
rect 26881 24151 26939 24157
rect 27111 24191 27160 24197
rect 27111 24157 27123 24191
rect 27157 24157 27160 24191
rect 27111 24151 27160 24157
rect 27154 24148 27160 24151
rect 27212 24148 27218 24200
rect 27706 24148 27712 24200
rect 27764 24148 27770 24200
rect 27890 24148 27896 24200
rect 27948 24148 27954 24200
rect 28074 24148 28080 24200
rect 28132 24188 28138 24200
rect 28813 24191 28871 24197
rect 28813 24188 28825 24191
rect 28132 24160 28825 24188
rect 28132 24148 28138 24160
rect 28813 24157 28825 24160
rect 28859 24157 28871 24191
rect 28813 24151 28871 24157
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 30024 24188 30052 24228
rect 30285 24225 30297 24228
rect 30331 24256 30343 24259
rect 30926 24256 30932 24268
rect 30331 24228 30932 24256
rect 30331 24225 30343 24228
rect 30285 24219 30343 24225
rect 30926 24216 30932 24228
rect 30984 24216 30990 24268
rect 31113 24259 31171 24265
rect 31113 24225 31125 24259
rect 31159 24256 31171 24259
rect 31478 24256 31484 24268
rect 31159 24228 31484 24256
rect 31159 24225 31171 24228
rect 31113 24219 31171 24225
rect 31478 24216 31484 24228
rect 31536 24216 31542 24268
rect 31570 24216 31576 24268
rect 31628 24256 31634 24268
rect 33226 24256 33232 24268
rect 31628 24228 33232 24256
rect 31628 24216 31634 24228
rect 33226 24216 33232 24228
rect 33284 24216 33290 24268
rect 33520 24228 33824 24256
rect 29512 24160 30052 24188
rect 30101 24191 30159 24197
rect 29512 24148 29518 24160
rect 30101 24157 30113 24191
rect 30147 24188 30159 24191
rect 30190 24188 30196 24200
rect 30147 24160 30196 24188
rect 30147 24157 30159 24160
rect 30101 24151 30159 24157
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 31205 24191 31263 24197
rect 31205 24157 31217 24191
rect 31251 24188 31263 24191
rect 31294 24188 31300 24200
rect 31251 24160 31300 24188
rect 31251 24157 31263 24160
rect 31205 24151 31263 24157
rect 31294 24148 31300 24160
rect 31352 24148 31358 24200
rect 32401 24191 32459 24197
rect 32401 24157 32413 24191
rect 32447 24188 32459 24191
rect 32766 24188 32772 24200
rect 32447 24160 32772 24188
rect 32447 24157 32459 24160
rect 32401 24151 32459 24157
rect 32766 24148 32772 24160
rect 32824 24188 32830 24200
rect 33520 24188 33548 24228
rect 32824 24160 33548 24188
rect 32824 24148 32830 24160
rect 33594 24148 33600 24200
rect 33652 24148 33658 24200
rect 33796 24197 33824 24228
rect 33870 24216 33876 24268
rect 33928 24216 33934 24268
rect 34072 24197 34100 24296
rect 35710 24284 35716 24296
rect 35768 24284 35774 24336
rect 37090 24284 37096 24336
rect 37148 24324 37154 24336
rect 37185 24327 37243 24333
rect 37185 24324 37197 24327
rect 37148 24296 37197 24324
rect 37148 24284 37154 24296
rect 37185 24293 37197 24296
rect 37231 24293 37243 24327
rect 37292 24324 37320 24364
rect 37366 24352 37372 24404
rect 37424 24352 37430 24404
rect 37458 24352 37464 24404
rect 37516 24392 37522 24404
rect 38105 24395 38163 24401
rect 38105 24392 38117 24395
rect 37516 24364 38117 24392
rect 37516 24352 37522 24364
rect 38105 24361 38117 24364
rect 38151 24361 38163 24395
rect 38105 24355 38163 24361
rect 40034 24352 40040 24404
rect 40092 24352 40098 24404
rect 40402 24352 40408 24404
rect 40460 24352 40466 24404
rect 41230 24352 41236 24404
rect 41288 24352 41294 24404
rect 42058 24352 42064 24404
rect 42116 24352 42122 24404
rect 37292 24296 38332 24324
rect 37185 24287 37243 24293
rect 34330 24216 34336 24268
rect 34388 24256 34394 24268
rect 37553 24259 37611 24265
rect 34388 24228 37136 24256
rect 34388 24216 34394 24228
rect 33781 24191 33839 24197
rect 33781 24157 33793 24191
rect 33827 24157 33839 24191
rect 33781 24151 33839 24157
rect 34057 24191 34115 24197
rect 34057 24157 34069 24191
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34238 24148 34244 24200
rect 34296 24148 34302 24200
rect 34422 24148 34428 24200
rect 34480 24188 34486 24200
rect 35069 24191 35127 24197
rect 35069 24188 35081 24191
rect 34480 24160 35081 24188
rect 34480 24148 34486 24160
rect 35069 24157 35081 24160
rect 35115 24188 35127 24191
rect 35437 24191 35495 24197
rect 35115 24160 35388 24188
rect 35115 24157 35127 24160
rect 35069 24151 35127 24157
rect 25884 24092 26832 24120
rect 26973 24123 27031 24129
rect 26973 24089 26985 24123
rect 27019 24120 27031 24123
rect 27908 24120 27936 24148
rect 27019 24092 27936 24120
rect 27019 24089 27031 24092
rect 26973 24083 27031 24089
rect 29178 24080 29184 24132
rect 29236 24120 29242 24132
rect 29236 24092 30420 24120
rect 29236 24080 29242 24092
rect 14642 24012 14648 24064
rect 14700 24012 14706 24064
rect 18138 24012 18144 24064
rect 18196 24012 18202 24064
rect 19613 24055 19671 24061
rect 19613 24021 19625 24055
rect 19659 24052 19671 24055
rect 20714 24052 20720 24064
rect 19659 24024 20720 24052
rect 19659 24021 19671 24024
rect 19613 24015 19671 24021
rect 20714 24012 20720 24024
rect 20772 24012 20778 24064
rect 20898 24012 20904 24064
rect 20956 24012 20962 24064
rect 21358 24012 21364 24064
rect 21416 24012 21422 24064
rect 22465 24055 22523 24061
rect 22465 24021 22477 24055
rect 22511 24052 22523 24055
rect 22554 24052 22560 24064
rect 22511 24024 22560 24052
rect 22511 24021 22523 24024
rect 22465 24015 22523 24021
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 25130 24012 25136 24064
rect 25188 24012 25194 24064
rect 27249 24055 27307 24061
rect 27249 24021 27261 24055
rect 27295 24052 27307 24055
rect 27338 24052 27344 24064
rect 27295 24024 27344 24052
rect 27295 24021 27307 24024
rect 27249 24015 27307 24021
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 28905 24055 28963 24061
rect 28905 24021 28917 24055
rect 28951 24052 28963 24055
rect 29733 24055 29791 24061
rect 29733 24052 29745 24055
rect 28951 24024 29745 24052
rect 28951 24021 28963 24024
rect 28905 24015 28963 24021
rect 29733 24021 29745 24024
rect 29779 24021 29791 24055
rect 29733 24015 29791 24021
rect 30193 24055 30251 24061
rect 30193 24021 30205 24055
rect 30239 24052 30251 24055
rect 30282 24052 30288 24064
rect 30239 24024 30288 24052
rect 30239 24021 30251 24024
rect 30193 24015 30251 24021
rect 30282 24012 30288 24024
rect 30340 24012 30346 24064
rect 30392 24052 30420 24092
rect 31386 24080 31392 24132
rect 31444 24120 31450 24132
rect 31481 24123 31539 24129
rect 31481 24120 31493 24123
rect 31444 24092 31493 24120
rect 31444 24080 31450 24092
rect 31481 24089 31493 24092
rect 31527 24089 31539 24123
rect 31481 24083 31539 24089
rect 32217 24055 32275 24061
rect 32217 24052 32229 24055
rect 30392 24024 32229 24052
rect 32217 24021 32229 24024
rect 32263 24052 32275 24055
rect 34146 24052 34152 24064
rect 32263 24024 34152 24052
rect 32263 24021 32275 24024
rect 32217 24015 32275 24021
rect 34146 24012 34152 24024
rect 34204 24012 34210 24064
rect 35250 24012 35256 24064
rect 35308 24012 35314 24064
rect 35360 24052 35388 24160
rect 35437 24157 35449 24191
rect 35483 24188 35495 24191
rect 36262 24188 36268 24200
rect 35483 24160 36268 24188
rect 35483 24157 35495 24160
rect 35437 24151 35495 24157
rect 36262 24148 36268 24160
rect 36320 24148 36326 24200
rect 36354 24148 36360 24200
rect 36412 24148 36418 24200
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24188 36599 24191
rect 36998 24188 37004 24200
rect 36587 24160 37004 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36998 24148 37004 24160
rect 37056 24148 37062 24200
rect 37108 24188 37136 24228
rect 37553 24225 37565 24259
rect 37599 24225 37611 24259
rect 37553 24219 37611 24225
rect 37200 24197 37412 24198
rect 37200 24191 37427 24197
rect 37200 24188 37381 24191
rect 37108 24170 37381 24188
rect 37108 24160 37228 24170
rect 37369 24157 37381 24170
rect 37415 24157 37427 24191
rect 37369 24151 37427 24157
rect 37568 24120 37596 24219
rect 37642 24148 37648 24200
rect 37700 24148 37706 24200
rect 38010 24148 38016 24200
rect 38068 24188 38074 24200
rect 38304 24197 38332 24296
rect 41322 24256 41328 24268
rect 38948 24228 41328 24256
rect 38105 24191 38163 24197
rect 38105 24188 38117 24191
rect 38068 24160 38117 24188
rect 38068 24148 38074 24160
rect 38105 24157 38117 24160
rect 38151 24157 38163 24191
rect 38105 24151 38163 24157
rect 38289 24191 38347 24197
rect 38289 24157 38301 24191
rect 38335 24188 38347 24191
rect 38378 24188 38384 24200
rect 38335 24160 38384 24188
rect 38335 24157 38347 24160
rect 38289 24151 38347 24157
rect 38378 24148 38384 24160
rect 38436 24148 38442 24200
rect 38948 24197 38976 24228
rect 41322 24216 41328 24228
rect 41380 24216 41386 24268
rect 41690 24216 41696 24268
rect 41748 24256 41754 24268
rect 42886 24256 42892 24268
rect 41748 24228 42892 24256
rect 41748 24216 41754 24228
rect 42886 24216 42892 24228
rect 42944 24216 42950 24268
rect 38933 24191 38991 24197
rect 38933 24157 38945 24191
rect 38979 24157 38991 24191
rect 38933 24151 38991 24157
rect 39117 24191 39175 24197
rect 39117 24157 39129 24191
rect 39163 24188 39175 24191
rect 39390 24188 39396 24200
rect 39163 24160 39396 24188
rect 39163 24157 39175 24160
rect 39117 24151 39175 24157
rect 39390 24148 39396 24160
rect 39448 24148 39454 24200
rect 39666 24148 39672 24200
rect 39724 24188 39730 24200
rect 40037 24191 40095 24197
rect 40037 24188 40049 24191
rect 39724 24160 40049 24188
rect 39724 24148 39730 24160
rect 40037 24157 40049 24160
rect 40083 24157 40095 24191
rect 40037 24151 40095 24157
rect 40126 24148 40132 24200
rect 40184 24148 40190 24200
rect 41417 24191 41475 24197
rect 41417 24157 41429 24191
rect 41463 24188 41475 24191
rect 41782 24188 41788 24200
rect 41463 24160 41788 24188
rect 41463 24157 41475 24160
rect 41417 24151 41475 24157
rect 41782 24148 41788 24160
rect 41840 24148 41846 24200
rect 41877 24191 41935 24197
rect 41877 24157 41889 24191
rect 41923 24188 41935 24191
rect 42426 24188 42432 24200
rect 41923 24160 42432 24188
rect 41923 24157 41935 24160
rect 41877 24151 41935 24157
rect 42426 24148 42432 24160
rect 42484 24148 42490 24200
rect 43257 24191 43315 24197
rect 43257 24157 43269 24191
rect 43303 24188 43315 24191
rect 43346 24188 43352 24200
rect 43303 24160 43352 24188
rect 43303 24157 43315 24160
rect 43257 24151 43315 24157
rect 43346 24148 43352 24160
rect 43404 24188 43410 24200
rect 43990 24188 43996 24200
rect 43404 24160 43996 24188
rect 43404 24148 43410 24160
rect 43990 24148 43996 24160
rect 44048 24148 44054 24200
rect 37568 24092 37688 24120
rect 36446 24052 36452 24064
rect 35360 24024 36452 24052
rect 36446 24012 36452 24024
rect 36504 24012 36510 24064
rect 37660 24052 37688 24092
rect 37826 24080 37832 24132
rect 37884 24120 37890 24132
rect 41690 24120 41696 24132
rect 37884 24092 41696 24120
rect 37884 24080 37890 24092
rect 41690 24080 41696 24092
rect 41748 24080 41754 24132
rect 41984 24092 43208 24120
rect 38010 24052 38016 24064
rect 37660 24024 38016 24052
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 38470 24012 38476 24064
rect 38528 24012 38534 24064
rect 38562 24012 38568 24064
rect 38620 24052 38626 24064
rect 39025 24055 39083 24061
rect 39025 24052 39037 24055
rect 38620 24024 39037 24052
rect 38620 24012 38626 24024
rect 39025 24021 39037 24024
rect 39071 24021 39083 24055
rect 39025 24015 39083 24021
rect 40954 24012 40960 24064
rect 41012 24052 41018 24064
rect 41984 24052 42012 24092
rect 43180 24064 43208 24092
rect 41012 24024 42012 24052
rect 41012 24012 41018 24024
rect 42334 24012 42340 24064
rect 42392 24052 42398 24064
rect 42518 24052 42524 24064
rect 42392 24024 42524 24052
rect 42392 24012 42398 24024
rect 42518 24012 42524 24024
rect 42576 24052 42582 24064
rect 42978 24052 42984 24064
rect 42576 24024 42984 24052
rect 42576 24012 42582 24024
rect 42978 24012 42984 24024
rect 43036 24012 43042 24064
rect 43162 24012 43168 24064
rect 43220 24012 43226 24064
rect 1104 23962 43884 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 43884 23962
rect 1104 23888 43884 23910
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14458 23848 14464 23860
rect 14139 23820 14464 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 14553 23851 14611 23857
rect 14553 23817 14565 23851
rect 14599 23848 14611 23851
rect 14734 23848 14740 23860
rect 14599 23820 14740 23848
rect 14599 23817 14611 23820
rect 14553 23811 14611 23817
rect 14734 23808 14740 23820
rect 14792 23848 14798 23860
rect 18138 23848 18144 23860
rect 14792 23820 18144 23848
rect 14792 23808 14798 23820
rect 18138 23808 18144 23820
rect 18196 23848 18202 23860
rect 21726 23848 21732 23860
rect 18196 23820 21732 23848
rect 18196 23808 18202 23820
rect 21726 23808 21732 23820
rect 21784 23808 21790 23860
rect 23661 23851 23719 23857
rect 23661 23848 23673 23851
rect 22296 23820 23673 23848
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 14700 23752 15700 23780
rect 14700 23740 14706 23752
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 14826 23712 14832 23724
rect 14507 23684 14832 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 15672 23721 15700 23752
rect 17862 23740 17868 23792
rect 17920 23780 17926 23792
rect 17920 23752 18920 23780
rect 17920 23740 17926 23752
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 15657 23715 15715 23721
rect 15657 23681 15669 23715
rect 15703 23681 15715 23715
rect 15657 23675 15715 23681
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23644 14795 23647
rect 15102 23644 15108 23656
rect 14783 23616 15108 23644
rect 14783 23613 14795 23616
rect 14737 23607 14795 23613
rect 13633 23579 13691 23585
rect 13633 23545 13645 23579
rect 13679 23576 13691 23579
rect 14752 23576 14780 23607
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 15580 23644 15608 23675
rect 17678 23672 17684 23724
rect 17736 23672 17742 23724
rect 18892 23721 18920 23752
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21818 23780 21824 23792
rect 21048 23752 21824 23780
rect 21048 23740 21054 23752
rect 21818 23740 21824 23752
rect 21876 23780 21882 23792
rect 22296 23789 22324 23820
rect 23661 23817 23673 23820
rect 23707 23848 23719 23851
rect 25866 23848 25872 23860
rect 23707 23820 25872 23848
rect 23707 23817 23719 23820
rect 23661 23811 23719 23817
rect 25866 23808 25872 23820
rect 25924 23808 25930 23860
rect 26418 23808 26424 23860
rect 26476 23848 26482 23860
rect 26605 23851 26663 23857
rect 26605 23848 26617 23851
rect 26476 23820 26617 23848
rect 26476 23808 26482 23820
rect 26605 23817 26617 23820
rect 26651 23817 26663 23851
rect 26605 23811 26663 23817
rect 29089 23851 29147 23857
rect 29089 23817 29101 23851
rect 29135 23848 29147 23851
rect 29135 23820 29776 23848
rect 29135 23817 29147 23820
rect 29089 23811 29147 23817
rect 22281 23783 22339 23789
rect 21876 23752 22232 23780
rect 21876 23740 21882 23752
rect 18509 23715 18567 23721
rect 18509 23681 18521 23715
rect 18555 23681 18567 23715
rect 18509 23675 18567 23681
rect 18877 23715 18935 23721
rect 18877 23681 18889 23715
rect 18923 23681 18935 23715
rect 18877 23675 18935 23681
rect 15436 23616 15608 23644
rect 15436 23604 15442 23616
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 18524 23644 18552 23675
rect 18966 23672 18972 23724
rect 19024 23672 19030 23724
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 20717 23715 20775 23721
rect 20717 23681 20729 23715
rect 20763 23712 20775 23715
rect 21358 23712 21364 23724
rect 20763 23684 21364 23712
rect 20763 23681 20775 23684
rect 20717 23675 20775 23681
rect 21358 23672 21364 23684
rect 21416 23672 21422 23724
rect 22204 23721 22232 23752
rect 22281 23749 22293 23783
rect 22327 23749 22339 23783
rect 22281 23743 22339 23749
rect 22370 23740 22376 23792
rect 22428 23740 22434 23792
rect 24302 23780 24308 23792
rect 22940 23752 24308 23780
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 22554 23672 22560 23724
rect 22612 23672 22618 23724
rect 17276 23616 18552 23644
rect 17276 23604 17282 23616
rect 18598 23604 18604 23656
rect 18656 23604 18662 23656
rect 21085 23647 21143 23653
rect 21085 23613 21097 23647
rect 21131 23644 21143 23647
rect 21266 23644 21272 23656
rect 21131 23616 21272 23644
rect 21131 23613 21143 23616
rect 21085 23607 21143 23613
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 22940 23644 22968 23752
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 24946 23740 24952 23792
rect 25004 23780 25010 23792
rect 25470 23783 25528 23789
rect 25470 23780 25482 23783
rect 25004 23752 25482 23780
rect 25004 23740 25010 23752
rect 25470 23749 25482 23752
rect 25516 23749 25528 23783
rect 25470 23743 25528 23749
rect 27614 23740 27620 23792
rect 27672 23780 27678 23792
rect 27672 23752 28028 23780
rect 27672 23740 27678 23752
rect 23017 23715 23075 23721
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 24486 23712 24492 23724
rect 23063 23684 24492 23712
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 24486 23672 24492 23684
rect 24544 23672 24550 23724
rect 24581 23715 24639 23721
rect 24581 23681 24593 23715
rect 24627 23712 24639 23715
rect 25958 23712 25964 23724
rect 24627 23684 25964 23712
rect 24627 23681 24639 23684
rect 24581 23675 24639 23681
rect 25958 23672 25964 23684
rect 26016 23672 26022 23724
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23712 27491 23715
rect 27798 23712 27804 23724
rect 27479 23684 27804 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 27890 23672 27896 23724
rect 27948 23672 27954 23724
rect 21324 23616 22968 23644
rect 21324 23604 21330 23616
rect 23750 23604 23756 23656
rect 23808 23644 23814 23656
rect 25225 23647 25283 23653
rect 25225 23644 25237 23647
rect 23808 23616 25237 23644
rect 23808 23604 23814 23616
rect 25225 23613 25237 23616
rect 25271 23613 25283 23647
rect 25225 23607 25283 23613
rect 27617 23647 27675 23653
rect 27617 23613 27629 23647
rect 27663 23644 27675 23647
rect 27706 23644 27712 23656
rect 27663 23616 27712 23644
rect 27663 23613 27675 23616
rect 27617 23607 27675 23613
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 28000 23644 28028 23752
rect 29178 23740 29184 23792
rect 29236 23780 29242 23792
rect 29454 23780 29460 23792
rect 29236 23752 29460 23780
rect 29236 23740 29242 23752
rect 29454 23740 29460 23752
rect 29512 23740 29518 23792
rect 29748 23780 29776 23820
rect 30282 23808 30288 23860
rect 30340 23808 30346 23860
rect 30742 23808 30748 23860
rect 30800 23808 30806 23860
rect 34330 23808 34336 23860
rect 34388 23808 34394 23860
rect 34790 23808 34796 23860
rect 34848 23848 34854 23860
rect 35253 23851 35311 23857
rect 35253 23848 35265 23851
rect 34848 23820 35265 23848
rect 34848 23808 34854 23820
rect 35253 23817 35265 23820
rect 35299 23817 35311 23851
rect 35253 23811 35311 23817
rect 35342 23808 35348 23860
rect 35400 23848 35406 23860
rect 35400 23820 39620 23848
rect 35400 23808 35406 23820
rect 30098 23780 30104 23792
rect 29748 23752 30104 23780
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23712 28779 23715
rect 28902 23712 28908 23724
rect 28767 23684 28908 23712
rect 28767 23681 28779 23684
rect 28721 23675 28779 23681
rect 28902 23672 28908 23684
rect 28960 23672 28966 23724
rect 28626 23644 28632 23656
rect 28000 23616 28632 23644
rect 28626 23604 28632 23616
rect 28684 23644 28690 23656
rect 29748 23653 29776 23752
rect 30098 23740 30104 23752
rect 30156 23740 30162 23792
rect 30190 23740 30196 23792
rect 30248 23780 30254 23792
rect 31757 23783 31815 23789
rect 31757 23780 31769 23783
rect 30248 23752 31769 23780
rect 30248 23740 30254 23752
rect 31757 23749 31769 23752
rect 31803 23780 31815 23783
rect 31846 23780 31852 23792
rect 31803 23752 31852 23780
rect 31803 23749 31815 23752
rect 31757 23743 31815 23749
rect 31846 23740 31852 23752
rect 31904 23740 31910 23792
rect 32309 23783 32367 23789
rect 32309 23749 32321 23783
rect 32355 23780 32367 23783
rect 32490 23780 32496 23792
rect 32355 23752 32496 23780
rect 32355 23749 32367 23752
rect 32309 23743 32367 23749
rect 32490 23740 32496 23752
rect 32548 23740 32554 23792
rect 33597 23783 33655 23789
rect 33597 23749 33609 23783
rect 33643 23780 33655 23783
rect 33686 23780 33692 23792
rect 33643 23752 33692 23780
rect 33643 23749 33655 23752
rect 33597 23743 33655 23749
rect 33686 23740 33692 23752
rect 33744 23780 33750 23792
rect 33744 23752 34468 23780
rect 33744 23740 33750 23752
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23712 29975 23715
rect 30374 23712 30380 23724
rect 29963 23684 30380 23712
rect 29963 23681 29975 23684
rect 29917 23675 29975 23681
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30834 23672 30840 23724
rect 30892 23712 30898 23724
rect 30929 23715 30987 23721
rect 30929 23712 30941 23715
rect 30892 23684 30941 23712
rect 30892 23672 30898 23684
rect 30929 23681 30941 23684
rect 30975 23681 30987 23715
rect 30929 23675 30987 23681
rect 31202 23672 31208 23724
rect 31260 23672 31266 23724
rect 32585 23715 32643 23721
rect 32585 23681 32597 23715
rect 32631 23712 32643 23715
rect 32674 23712 32680 23724
rect 32631 23684 32680 23712
rect 32631 23681 32643 23684
rect 32585 23675 32643 23681
rect 32674 23672 32680 23684
rect 32732 23672 32738 23724
rect 33502 23672 33508 23724
rect 33560 23672 33566 23724
rect 33781 23715 33839 23721
rect 33781 23681 33793 23715
rect 33827 23712 33839 23715
rect 34146 23712 34152 23724
rect 33827 23684 34152 23712
rect 33827 23681 33839 23684
rect 33781 23675 33839 23681
rect 34146 23672 34152 23684
rect 34204 23672 34210 23724
rect 34238 23672 34244 23724
rect 34296 23672 34302 23724
rect 34440 23721 34468 23752
rect 34698 23740 34704 23792
rect 34756 23780 34762 23792
rect 34885 23783 34943 23789
rect 34885 23780 34897 23783
rect 34756 23752 34897 23780
rect 34756 23740 34762 23752
rect 34885 23749 34897 23752
rect 34931 23749 34943 23783
rect 37826 23780 37832 23792
rect 34885 23743 34943 23749
rect 37660 23752 37832 23780
rect 34425 23715 34483 23721
rect 34425 23681 34437 23715
rect 34471 23712 34483 23715
rect 35069 23715 35127 23721
rect 34471 23684 35020 23712
rect 34471 23681 34483 23684
rect 34425 23675 34483 23681
rect 28813 23647 28871 23653
rect 28813 23644 28825 23647
rect 28684 23616 28825 23644
rect 28684 23604 28690 23616
rect 28813 23613 28825 23616
rect 28859 23613 28871 23647
rect 28813 23607 28871 23613
rect 29733 23647 29791 23653
rect 29733 23613 29745 23647
rect 29779 23613 29791 23647
rect 29733 23607 29791 23613
rect 29825 23647 29883 23653
rect 29825 23613 29837 23647
rect 29871 23644 29883 23647
rect 30282 23644 30288 23656
rect 29871 23616 30288 23644
rect 29871 23613 29883 23616
rect 29825 23607 29883 23613
rect 13679 23548 14780 23576
rect 17957 23579 18015 23585
rect 13679 23545 13691 23548
rect 13633 23539 13691 23545
rect 17957 23545 17969 23579
rect 18003 23576 18015 23579
rect 24765 23579 24823 23585
rect 18003 23548 24348 23576
rect 18003 23545 18015 23548
rect 17957 23539 18015 23545
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16298 23508 16304 23520
rect 15979 23480 16304 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16298 23468 16304 23480
rect 16356 23468 16362 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20441 23511 20499 23517
rect 20441 23508 20453 23511
rect 20128 23480 20453 23508
rect 20128 23468 20134 23480
rect 20441 23477 20453 23480
rect 20487 23477 20499 23511
rect 20441 23471 20499 23477
rect 22005 23511 22063 23517
rect 22005 23477 22017 23511
rect 22051 23508 22063 23511
rect 22554 23508 22560 23520
rect 22051 23480 22560 23508
rect 22051 23477 22063 23480
rect 22005 23471 22063 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 23201 23511 23259 23517
rect 23201 23477 23213 23511
rect 23247 23508 23259 23511
rect 23474 23508 23480 23520
rect 23247 23480 23480 23508
rect 23247 23477 23259 23480
rect 23201 23471 23259 23477
rect 23474 23468 23480 23480
rect 23532 23468 23538 23520
rect 24320 23508 24348 23548
rect 24765 23545 24777 23579
rect 24811 23576 24823 23579
rect 24946 23576 24952 23588
rect 24811 23548 24952 23576
rect 24811 23545 24823 23548
rect 24765 23539 24823 23545
rect 24946 23536 24952 23548
rect 25004 23536 25010 23588
rect 26602 23536 26608 23588
rect 26660 23576 26666 23588
rect 26660 23548 27292 23576
rect 26660 23536 26666 23548
rect 27264 23520 27292 23548
rect 27430 23536 27436 23588
rect 27488 23576 27494 23588
rect 27488 23548 27844 23576
rect 27488 23536 27494 23548
rect 26694 23508 26700 23520
rect 24320 23480 26700 23508
rect 26694 23468 26700 23480
rect 26752 23468 26758 23520
rect 27154 23468 27160 23520
rect 27212 23468 27218 23520
rect 27246 23468 27252 23520
rect 27304 23508 27310 23520
rect 27525 23511 27583 23517
rect 27525 23508 27537 23511
rect 27304 23480 27537 23508
rect 27304 23468 27310 23480
rect 27525 23477 27537 23480
rect 27571 23477 27583 23511
rect 27525 23471 27583 23477
rect 27614 23468 27620 23520
rect 27672 23508 27678 23520
rect 27709 23511 27767 23517
rect 27709 23508 27721 23511
rect 27672 23480 27721 23508
rect 27672 23468 27678 23480
rect 27709 23477 27721 23480
rect 27755 23477 27767 23511
rect 27816 23508 27844 23548
rect 28994 23536 29000 23588
rect 29052 23576 29058 23588
rect 29840 23576 29868 23607
rect 30282 23604 30288 23616
rect 30340 23604 30346 23656
rect 31110 23604 31116 23656
rect 31168 23604 31174 23656
rect 32030 23604 32036 23656
rect 32088 23644 32094 23656
rect 32493 23647 32551 23653
rect 32493 23644 32505 23647
rect 32088 23616 32505 23644
rect 32088 23604 32094 23616
rect 32493 23613 32505 23616
rect 32539 23613 32551 23647
rect 34992 23644 35020 23684
rect 35069 23681 35081 23715
rect 35115 23712 35127 23715
rect 35434 23712 35440 23724
rect 35115 23684 35440 23712
rect 35115 23681 35127 23684
rect 35069 23675 35127 23681
rect 35434 23672 35440 23684
rect 35492 23712 35498 23724
rect 35710 23712 35716 23724
rect 35492 23684 35716 23712
rect 35492 23672 35498 23684
rect 35710 23672 35716 23684
rect 35768 23672 35774 23724
rect 35897 23715 35955 23721
rect 35897 23681 35909 23715
rect 35943 23712 35955 23715
rect 36262 23712 36268 23724
rect 35943 23684 36268 23712
rect 35943 23681 35955 23684
rect 35897 23675 35955 23681
rect 36262 23672 36268 23684
rect 36320 23672 36326 23724
rect 36357 23715 36415 23721
rect 36357 23681 36369 23715
rect 36403 23712 36415 23715
rect 36538 23712 36544 23724
rect 36403 23684 36544 23712
rect 36403 23681 36415 23684
rect 36357 23675 36415 23681
rect 36538 23672 36544 23684
rect 36596 23672 36602 23724
rect 37660 23721 37688 23752
rect 37826 23740 37832 23752
rect 37884 23740 37890 23792
rect 39022 23740 39028 23792
rect 39080 23740 39086 23792
rect 39206 23740 39212 23792
rect 39264 23780 39270 23792
rect 39264 23752 39344 23780
rect 39264 23740 39270 23752
rect 37645 23715 37703 23721
rect 37645 23681 37657 23715
rect 37691 23681 37703 23715
rect 37645 23675 37703 23681
rect 38105 23715 38163 23721
rect 38105 23681 38117 23715
rect 38151 23712 38163 23715
rect 38286 23712 38292 23724
rect 38151 23684 38292 23712
rect 38151 23681 38163 23684
rect 38105 23675 38163 23681
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 39316 23721 39344 23752
rect 39301 23715 39359 23721
rect 39301 23681 39313 23715
rect 39347 23681 39359 23715
rect 39301 23675 39359 23681
rect 39482 23672 39488 23724
rect 39540 23672 39546 23724
rect 39592 23712 39620 23820
rect 39666 23808 39672 23860
rect 39724 23808 39730 23860
rect 40678 23808 40684 23860
rect 40736 23808 40742 23860
rect 42978 23808 42984 23860
rect 43036 23808 43042 23860
rect 40773 23783 40831 23789
rect 40773 23749 40785 23783
rect 40819 23780 40831 23783
rect 42334 23780 42340 23792
rect 40819 23752 42340 23780
rect 40819 23749 40831 23752
rect 40773 23743 40831 23749
rect 42334 23740 42340 23752
rect 42392 23740 42398 23792
rect 41325 23715 41383 23721
rect 41325 23712 41337 23715
rect 39592 23684 41337 23712
rect 41325 23681 41337 23684
rect 41371 23681 41383 23715
rect 41325 23675 41383 23681
rect 41506 23672 41512 23724
rect 41564 23672 41570 23724
rect 42794 23672 42800 23724
rect 42852 23672 42858 23724
rect 35342 23644 35348 23656
rect 34992 23616 35348 23644
rect 32493 23607 32551 23613
rect 35342 23604 35348 23616
rect 35400 23604 35406 23656
rect 35618 23604 35624 23656
rect 35676 23644 35682 23656
rect 36081 23647 36139 23653
rect 36081 23644 36093 23647
rect 35676 23616 36093 23644
rect 35676 23604 35682 23616
rect 36081 23613 36093 23616
rect 36127 23613 36139 23647
rect 36081 23607 36139 23613
rect 36173 23647 36231 23653
rect 36173 23613 36185 23647
rect 36219 23644 36231 23647
rect 36909 23647 36967 23653
rect 36909 23644 36921 23647
rect 36219 23616 36921 23644
rect 36219 23613 36231 23616
rect 36173 23607 36231 23613
rect 36909 23613 36921 23616
rect 36955 23644 36967 23647
rect 37090 23644 37096 23656
rect 36955 23616 37096 23644
rect 36955 23613 36967 23616
rect 36909 23607 36967 23613
rect 37090 23604 37096 23616
rect 37148 23604 37154 23656
rect 37458 23604 37464 23656
rect 37516 23644 37522 23656
rect 37737 23647 37795 23653
rect 37737 23644 37749 23647
rect 37516 23616 37749 23644
rect 37516 23604 37522 23616
rect 37737 23613 37749 23616
rect 37783 23613 37795 23647
rect 37737 23607 37795 23613
rect 37826 23604 37832 23656
rect 37884 23644 37890 23656
rect 40678 23644 40684 23656
rect 37884 23616 40684 23644
rect 37884 23604 37890 23616
rect 40678 23604 40684 23616
rect 40736 23604 40742 23656
rect 29052 23548 29868 23576
rect 29052 23536 29058 23548
rect 32858 23536 32864 23588
rect 32916 23576 32922 23588
rect 33781 23579 33839 23585
rect 33781 23576 33793 23579
rect 32916 23548 33793 23576
rect 32916 23536 32922 23548
rect 33781 23545 33793 23548
rect 33827 23576 33839 23579
rect 35434 23576 35440 23588
rect 33827 23548 35440 23576
rect 33827 23545 33839 23548
rect 33781 23539 33839 23545
rect 35434 23536 35440 23548
rect 35492 23536 35498 23588
rect 35802 23536 35808 23588
rect 35860 23576 35866 23588
rect 35989 23579 36047 23585
rect 35989 23576 36001 23579
rect 35860 23548 36001 23576
rect 35860 23536 35866 23548
rect 35989 23545 36001 23548
rect 36035 23545 36047 23579
rect 35989 23539 36047 23545
rect 36446 23536 36452 23588
rect 36504 23576 36510 23588
rect 41138 23576 41144 23588
rect 36504 23548 41144 23576
rect 36504 23536 36510 23548
rect 41138 23536 41144 23548
rect 41196 23536 41202 23588
rect 28721 23511 28779 23517
rect 28721 23508 28733 23511
rect 27816 23480 28733 23508
rect 27709 23471 27767 23477
rect 28721 23477 28733 23480
rect 28767 23508 28779 23511
rect 29546 23508 29552 23520
rect 28767 23480 29552 23508
rect 28767 23477 28779 23480
rect 28721 23471 28779 23477
rect 29546 23468 29552 23480
rect 29604 23468 29610 23520
rect 31205 23511 31263 23517
rect 31205 23477 31217 23511
rect 31251 23508 31263 23511
rect 32306 23508 32312 23520
rect 31251 23480 32312 23508
rect 31251 23477 31263 23480
rect 31205 23471 31263 23477
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 32398 23468 32404 23520
rect 32456 23468 32462 23520
rect 35713 23511 35771 23517
rect 35713 23477 35725 23511
rect 35759 23508 35771 23511
rect 35894 23508 35900 23520
rect 35759 23480 35900 23508
rect 35759 23477 35771 23480
rect 35713 23471 35771 23477
rect 35894 23468 35900 23480
rect 35952 23468 35958 23520
rect 37458 23468 37464 23520
rect 37516 23468 37522 23520
rect 37642 23468 37648 23520
rect 37700 23468 37706 23520
rect 38378 23468 38384 23520
rect 38436 23508 38442 23520
rect 39117 23511 39175 23517
rect 39117 23508 39129 23511
rect 38436 23480 39129 23508
rect 38436 23468 38442 23480
rect 39117 23477 39129 23480
rect 39163 23477 39175 23511
rect 39117 23471 39175 23477
rect 1104 23418 43884 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 43884 23418
rect 1104 23344 43884 23366
rect 15749 23307 15807 23313
rect 15749 23273 15761 23307
rect 15795 23304 15807 23307
rect 17678 23304 17684 23316
rect 15795 23276 17684 23304
rect 15795 23273 15807 23276
rect 15749 23267 15807 23273
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 20806 23304 20812 23316
rect 19720 23276 20812 23304
rect 14277 23239 14335 23245
rect 14277 23205 14289 23239
rect 14323 23205 14335 23239
rect 14277 23199 14335 23205
rect 14292 23168 14320 23199
rect 15470 23196 15476 23248
rect 15528 23196 15534 23248
rect 16577 23239 16635 23245
rect 16577 23205 16589 23239
rect 16623 23236 16635 23239
rect 18230 23236 18236 23248
rect 16623 23208 18236 23236
rect 16623 23205 16635 23208
rect 16577 23199 16635 23205
rect 18230 23196 18236 23208
rect 18288 23196 18294 23248
rect 15488 23168 15516 23196
rect 15746 23168 15752 23180
rect 14292 23140 15148 23168
rect 13633 23103 13691 23109
rect 13633 23069 13645 23103
rect 13679 23100 13691 23103
rect 14274 23100 14280 23112
rect 13679 23072 14280 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 15120 23109 15148 23140
rect 15304 23140 15752 23168
rect 15304 23109 15332 23140
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 17034 23128 17040 23180
rect 17092 23128 17098 23180
rect 17862 23128 17868 23180
rect 17920 23128 17926 23180
rect 19720 23177 19748 23276
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 21910 23264 21916 23316
rect 21968 23264 21974 23316
rect 22373 23307 22431 23313
rect 22373 23273 22385 23307
rect 22419 23304 22431 23307
rect 22830 23304 22836 23316
rect 22419 23276 22836 23304
rect 22419 23273 22431 23276
rect 22373 23267 22431 23273
rect 22830 23264 22836 23276
rect 22888 23264 22894 23316
rect 25958 23264 25964 23316
rect 26016 23264 26022 23316
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 31113 23307 31171 23313
rect 31113 23304 31125 23307
rect 28960 23276 31125 23304
rect 28960 23264 28966 23276
rect 31113 23273 31125 23276
rect 31159 23304 31171 23307
rect 31386 23304 31392 23316
rect 31159 23276 31392 23304
rect 31159 23273 31171 23276
rect 31113 23267 31171 23273
rect 31386 23264 31392 23276
rect 31444 23264 31450 23316
rect 33137 23307 33195 23313
rect 33137 23273 33149 23307
rect 33183 23304 33195 23307
rect 33226 23304 33232 23316
rect 33183 23276 33232 23304
rect 33183 23273 33195 23276
rect 33137 23267 33195 23273
rect 33226 23264 33232 23276
rect 33284 23264 33290 23316
rect 33502 23264 33508 23316
rect 33560 23304 33566 23316
rect 33962 23304 33968 23316
rect 33560 23276 33968 23304
rect 33560 23264 33566 23276
rect 33962 23264 33968 23276
rect 34020 23264 34026 23316
rect 35345 23307 35403 23313
rect 35345 23273 35357 23307
rect 35391 23304 35403 23307
rect 36722 23304 36728 23316
rect 35391 23276 36728 23304
rect 35391 23273 35403 23276
rect 35345 23267 35403 23273
rect 36722 23264 36728 23276
rect 36780 23304 36786 23316
rect 36817 23307 36875 23313
rect 36817 23304 36829 23307
rect 36780 23276 36829 23304
rect 36780 23264 36786 23276
rect 36817 23273 36829 23276
rect 36863 23273 36875 23307
rect 36817 23267 36875 23273
rect 38289 23307 38347 23313
rect 38289 23273 38301 23307
rect 38335 23304 38347 23307
rect 38470 23304 38476 23316
rect 38335 23276 38476 23304
rect 38335 23273 38347 23276
rect 38289 23267 38347 23273
rect 38470 23264 38476 23276
rect 38528 23304 38534 23316
rect 38654 23304 38660 23316
rect 38528 23276 38660 23304
rect 38528 23264 38534 23276
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 39206 23264 39212 23316
rect 39264 23304 39270 23316
rect 39301 23307 39359 23313
rect 39301 23304 39313 23307
rect 39264 23276 39313 23304
rect 39264 23264 39270 23276
rect 39301 23273 39313 23276
rect 39347 23273 39359 23307
rect 39301 23267 39359 23273
rect 40218 23264 40224 23316
rect 40276 23264 40282 23316
rect 41506 23264 41512 23316
rect 41564 23304 41570 23316
rect 41693 23307 41751 23313
rect 41693 23304 41705 23307
rect 41564 23276 41705 23304
rect 41564 23264 41570 23276
rect 41693 23273 41705 23276
rect 41739 23273 41751 23307
rect 41693 23267 41751 23273
rect 41782 23264 41788 23316
rect 41840 23304 41846 23316
rect 41877 23307 41935 23313
rect 41877 23304 41889 23307
rect 41840 23276 41889 23304
rect 41840 23264 41846 23276
rect 41877 23273 41889 23276
rect 41923 23273 41935 23307
rect 41877 23267 41935 23273
rect 42797 23307 42855 23313
rect 42797 23273 42809 23307
rect 42843 23304 42855 23307
rect 42886 23304 42892 23316
rect 42843 23276 42892 23304
rect 42843 23273 42855 23276
rect 42797 23267 42855 23273
rect 42886 23264 42892 23276
rect 42944 23264 42950 23316
rect 19981 23239 20039 23245
rect 19981 23205 19993 23239
rect 20027 23236 20039 23239
rect 20027 23208 20576 23236
rect 20027 23205 20039 23208
rect 19981 23199 20039 23205
rect 20548 23177 20576 23208
rect 31294 23196 31300 23248
rect 31352 23236 31358 23248
rect 32585 23239 32643 23245
rect 32585 23236 32597 23239
rect 31352 23208 32597 23236
rect 31352 23196 31358 23208
rect 32585 23205 32597 23208
rect 32631 23236 32643 23239
rect 37090 23236 37096 23248
rect 32631 23208 37096 23236
rect 32631 23205 32643 23208
rect 32585 23199 32643 23205
rect 37090 23196 37096 23208
rect 37148 23196 37154 23248
rect 37277 23239 37335 23245
rect 37277 23205 37289 23239
rect 37323 23236 37335 23239
rect 40497 23239 40555 23245
rect 37323 23208 40172 23236
rect 37323 23205 37335 23208
rect 37277 23199 37335 23205
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23137 20591 23171
rect 20533 23131 20591 23137
rect 23750 23128 23756 23180
rect 23808 23128 23814 23180
rect 24762 23128 24768 23180
rect 24820 23128 24826 23180
rect 25130 23128 25136 23180
rect 25188 23168 25194 23180
rect 25225 23171 25283 23177
rect 25225 23168 25237 23171
rect 25188 23140 25237 23168
rect 25188 23128 25194 23140
rect 25225 23137 25237 23140
rect 25271 23137 25283 23171
rect 25225 23131 25283 23137
rect 26605 23171 26663 23177
rect 26605 23137 26617 23171
rect 26651 23168 26663 23171
rect 27154 23168 27160 23180
rect 26651 23140 27160 23168
rect 26651 23137 26663 23140
rect 26605 23131 26663 23137
rect 27154 23128 27160 23140
rect 27212 23128 27218 23180
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23168 27583 23171
rect 27798 23168 27804 23180
rect 27571 23140 27804 23168
rect 27571 23137 27583 23140
rect 27525 23131 27583 23137
rect 27798 23128 27804 23140
rect 27856 23128 27862 23180
rect 31938 23128 31944 23180
rect 31996 23168 32002 23180
rect 31996 23140 34560 23168
rect 31996 23128 32002 23140
rect 15105 23103 15163 23109
rect 15105 23069 15117 23103
rect 15151 23069 15163 23103
rect 15105 23063 15163 23069
rect 15289 23103 15347 23109
rect 15289 23069 15301 23103
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 15378 23060 15384 23112
rect 15436 23060 15442 23112
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 15519 23072 15700 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 14458 22992 14464 23044
rect 14516 22992 14522 23044
rect 14645 23035 14703 23041
rect 14645 23001 14657 23035
rect 14691 23032 14703 23035
rect 15562 23032 15568 23044
rect 14691 23004 15568 23032
rect 14691 23001 14703 23004
rect 14645 22995 14703 23001
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 13449 22967 13507 22973
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 13538 22964 13544 22976
rect 13495 22936 13544 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 15672 22964 15700 23072
rect 16298 23060 16304 23112
rect 16356 23060 16362 23112
rect 17218 23060 17224 23112
rect 17276 23060 17282 23112
rect 17586 23060 17592 23112
rect 17644 23060 17650 23112
rect 18598 23060 18604 23112
rect 18656 23100 18662 23112
rect 18785 23103 18843 23109
rect 18785 23100 18797 23103
rect 18656 23072 18797 23100
rect 18656 23060 18662 23072
rect 18785 23069 18797 23072
rect 18831 23069 18843 23103
rect 18785 23063 18843 23069
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 19392 23072 19625 23100
rect 19392 23060 19398 23072
rect 19613 23069 19625 23072
rect 19659 23100 19671 23103
rect 19978 23100 19984 23112
rect 19659 23072 19984 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20898 23100 20904 23112
rect 20671 23072 20904 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 23474 23060 23480 23112
rect 23532 23109 23538 23112
rect 23532 23100 23544 23109
rect 23532 23072 23577 23100
rect 23532 23063 23544 23072
rect 23532 23060 23538 23063
rect 24854 23060 24860 23112
rect 24912 23060 24918 23112
rect 26329 23103 26387 23109
rect 26329 23069 26341 23103
rect 26375 23100 26387 23103
rect 26418 23100 26424 23112
rect 26375 23072 26424 23100
rect 26375 23069 26387 23072
rect 26329 23063 26387 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 27338 23060 27344 23112
rect 27396 23060 27402 23112
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 28350 23100 28356 23112
rect 27663 23072 28356 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 28721 23103 28779 23109
rect 28721 23069 28733 23103
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23100 28871 23103
rect 28902 23100 28908 23112
rect 28859 23072 28908 23100
rect 28859 23069 28871 23072
rect 28813 23063 28871 23069
rect 17236 23032 17264 23060
rect 17678 23032 17684 23044
rect 17236 23004 17684 23032
rect 17678 22992 17684 23004
rect 17736 22992 17742 23044
rect 19058 22992 19064 23044
rect 19116 23032 19122 23044
rect 28736 23032 28764 23063
rect 28902 23060 28908 23072
rect 28960 23060 28966 23112
rect 28997 23103 29055 23109
rect 28997 23069 29009 23103
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23100 29791 23103
rect 33134 23100 33140 23112
rect 29779 23072 33140 23100
rect 29779 23069 29791 23072
rect 29733 23063 29791 23069
rect 19116 23004 28764 23032
rect 19116 22992 19122 23004
rect 14884 22936 15700 22964
rect 14884 22924 14890 22936
rect 18506 22924 18512 22976
rect 18564 22964 18570 22976
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 18564 22936 18613 22964
rect 18564 22924 18570 22936
rect 18601 22933 18613 22936
rect 18647 22933 18659 22967
rect 18601 22927 18659 22933
rect 20990 22924 20996 22976
rect 21048 22924 21054 22976
rect 24026 22924 24032 22976
rect 24084 22964 24090 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24084 22936 24593 22964
rect 24084 22924 24090 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 26421 22967 26479 22973
rect 26421 22933 26433 22967
rect 26467 22964 26479 22967
rect 27157 22967 27215 22973
rect 27157 22964 27169 22967
rect 26467 22936 27169 22964
rect 26467 22933 26479 22936
rect 26421 22927 26479 22933
rect 27157 22933 27169 22936
rect 27203 22933 27215 22967
rect 27157 22927 27215 22933
rect 28166 22924 28172 22976
rect 28224 22924 28230 22976
rect 28736 22964 28764 23004
rect 28902 22964 28908 22976
rect 28736 22936 28908 22964
rect 28902 22924 28908 22936
rect 28960 22924 28966 22976
rect 29012 22964 29040 23063
rect 33134 23060 33140 23072
rect 33192 23100 33198 23112
rect 33870 23100 33876 23112
rect 33192 23072 33876 23100
rect 33192 23060 33198 23072
rect 33870 23060 33876 23072
rect 33928 23060 33934 23112
rect 34532 23100 34560 23140
rect 34698 23128 34704 23180
rect 34756 23168 34762 23180
rect 37001 23171 37059 23177
rect 34756 23140 35204 23168
rect 34756 23128 34762 23140
rect 34790 23100 34796 23112
rect 34532 23072 34796 23100
rect 34790 23060 34796 23072
rect 34848 23060 34854 23112
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23069 34943 23103
rect 34885 23063 34943 23069
rect 29181 23035 29239 23041
rect 29181 23001 29193 23035
rect 29227 23032 29239 23035
rect 29978 23035 30036 23041
rect 29978 23032 29990 23035
rect 29227 23004 29990 23032
rect 29227 23001 29239 23004
rect 29181 22995 29239 23001
rect 29978 23001 29990 23004
rect 30024 23001 30036 23035
rect 29978 22995 30036 23001
rect 30282 22992 30288 23044
rect 30340 23032 30346 23044
rect 30340 23004 31892 23032
rect 30340 22992 30346 23004
rect 30190 22964 30196 22976
rect 29012 22936 30196 22964
rect 30190 22924 30196 22936
rect 30248 22924 30254 22976
rect 31662 22924 31668 22976
rect 31720 22924 31726 22976
rect 31864 22964 31892 23004
rect 31938 22992 31944 23044
rect 31996 22992 32002 23044
rect 32416 23004 33548 23032
rect 32416 22964 32444 23004
rect 31864 22936 32444 22964
rect 33520 22964 33548 23004
rect 33594 22992 33600 23044
rect 33652 22992 33658 23044
rect 33778 22992 33784 23044
rect 33836 22992 33842 23044
rect 34900 23032 34928 23063
rect 34974 23060 34980 23112
rect 35032 23060 35038 23112
rect 35176 23109 35204 23140
rect 37001 23137 37013 23171
rect 37047 23168 37059 23171
rect 37826 23168 37832 23180
rect 37047 23140 37832 23168
rect 37047 23137 37059 23140
rect 37001 23131 37059 23137
rect 37826 23128 37832 23140
rect 37884 23168 37890 23180
rect 38105 23171 38163 23177
rect 37884 23140 38056 23168
rect 37884 23128 37890 23140
rect 35161 23103 35219 23109
rect 35161 23069 35173 23103
rect 35207 23069 35219 23103
rect 35161 23063 35219 23069
rect 35986 23060 35992 23112
rect 36044 23100 36050 23112
rect 37093 23103 37151 23109
rect 36044 23072 37044 23100
rect 36044 23060 36050 23072
rect 35618 23032 35624 23044
rect 33888 23004 35624 23032
rect 33888 22964 33916 23004
rect 35618 22992 35624 23004
rect 35676 22992 35682 23044
rect 36814 22992 36820 23044
rect 36872 22992 36878 23044
rect 37016 23032 37044 23072
rect 37093 23069 37105 23103
rect 37139 23100 37151 23103
rect 37182 23100 37188 23112
rect 37139 23072 37188 23100
rect 37139 23069 37151 23072
rect 37093 23063 37151 23069
rect 37182 23060 37188 23072
rect 37240 23060 37246 23112
rect 37550 23060 37556 23112
rect 37608 23100 37614 23112
rect 37921 23103 37979 23109
rect 37921 23100 37933 23103
rect 37608 23072 37933 23100
rect 37608 23060 37614 23072
rect 37921 23069 37933 23072
rect 37967 23069 37979 23103
rect 38028 23100 38056 23140
rect 38105 23137 38117 23171
rect 38151 23168 38163 23171
rect 38746 23168 38752 23180
rect 38151 23140 38752 23168
rect 38151 23137 38163 23140
rect 38105 23131 38163 23137
rect 38746 23128 38752 23140
rect 38804 23128 38810 23180
rect 38838 23128 38844 23180
rect 38896 23168 38902 23180
rect 39298 23168 39304 23180
rect 38896 23140 39304 23168
rect 38896 23128 38902 23140
rect 39298 23128 39304 23140
rect 39356 23128 39362 23180
rect 40144 23177 40172 23208
rect 40497 23205 40509 23239
rect 40543 23236 40555 23239
rect 43070 23236 43076 23248
rect 40543 23208 43076 23236
rect 40543 23205 40555 23208
rect 40497 23199 40555 23205
rect 43070 23196 43076 23208
rect 43128 23196 43134 23248
rect 40129 23171 40187 23177
rect 40129 23137 40141 23171
rect 40175 23137 40187 23171
rect 40129 23131 40187 23137
rect 41966 23128 41972 23180
rect 42024 23168 42030 23180
rect 42061 23171 42119 23177
rect 42061 23168 42073 23171
rect 42024 23140 42073 23168
rect 42024 23128 42030 23140
rect 42061 23137 42073 23140
rect 42107 23168 42119 23171
rect 42886 23168 42892 23180
rect 42107 23140 42892 23168
rect 42107 23137 42119 23140
rect 42061 23131 42119 23137
rect 42886 23128 42892 23140
rect 42944 23128 42950 23180
rect 38562 23100 38568 23112
rect 38028 23072 38568 23100
rect 37921 23063 37979 23069
rect 38562 23060 38568 23072
rect 38620 23060 38626 23112
rect 39206 23060 39212 23112
rect 39264 23060 39270 23112
rect 39393 23103 39451 23109
rect 39393 23069 39405 23103
rect 39439 23069 39451 23103
rect 39393 23063 39451 23069
rect 37016 23004 38240 23032
rect 33520 22936 33916 22964
rect 35897 22967 35955 22973
rect 35897 22933 35909 22967
rect 35943 22964 35955 22967
rect 36262 22964 36268 22976
rect 35943 22936 36268 22964
rect 35943 22933 35955 22936
rect 35897 22927 35955 22933
rect 36262 22924 36268 22936
rect 36320 22964 36326 22976
rect 37550 22964 37556 22976
rect 36320 22936 37556 22964
rect 36320 22924 36326 22936
rect 37550 22924 37556 22936
rect 37608 22924 37614 22976
rect 37642 22924 37648 22976
rect 37700 22964 37706 22976
rect 37737 22967 37795 22973
rect 37737 22964 37749 22967
rect 37700 22936 37749 22964
rect 37700 22924 37706 22936
rect 37737 22933 37749 22936
rect 37783 22933 37795 22967
rect 38212 22964 38240 23004
rect 38286 22992 38292 23044
rect 38344 23032 38350 23044
rect 38381 23035 38439 23041
rect 38381 23032 38393 23035
rect 38344 23004 38393 23032
rect 38344 22992 38350 23004
rect 38381 23001 38393 23004
rect 38427 23001 38439 23035
rect 38381 22995 38439 23001
rect 39298 22964 39304 22976
rect 38212 22936 39304 22964
rect 37737 22927 37795 22933
rect 39298 22924 39304 22936
rect 39356 22964 39362 22976
rect 39408 22964 39436 23063
rect 39482 23060 39488 23112
rect 39540 23100 39546 23112
rect 40313 23103 40371 23109
rect 40313 23100 40325 23103
rect 39540 23072 40325 23100
rect 39540 23060 39546 23072
rect 40313 23069 40325 23072
rect 40359 23069 40371 23103
rect 40313 23063 40371 23069
rect 41874 23060 41880 23112
rect 41932 23100 41938 23112
rect 42702 23100 42708 23112
rect 41932 23072 42708 23100
rect 41932 23060 41938 23072
rect 42702 23060 42708 23072
rect 42760 23100 42766 23112
rect 42797 23103 42855 23109
rect 42797 23100 42809 23103
rect 42760 23072 42809 23100
rect 42760 23060 42766 23072
rect 42797 23069 42809 23072
rect 42843 23069 42855 23103
rect 42797 23063 42855 23069
rect 42981 23103 43039 23109
rect 42981 23069 42993 23103
rect 43027 23069 43039 23103
rect 42981 23063 43039 23069
rect 39758 22992 39764 23044
rect 39816 23032 39822 23044
rect 40037 23035 40095 23041
rect 40037 23032 40049 23035
rect 39816 23004 40049 23032
rect 39816 22992 39822 23004
rect 40037 23001 40049 23004
rect 40083 23001 40095 23035
rect 40037 22995 40095 23001
rect 42337 23035 42395 23041
rect 42337 23001 42349 23035
rect 42383 23032 42395 23035
rect 42426 23032 42432 23044
rect 42383 23004 42432 23032
rect 42383 23001 42395 23004
rect 42337 22995 42395 23001
rect 42426 22992 42432 23004
rect 42484 23032 42490 23044
rect 42996 23032 43024 23063
rect 43070 23032 43076 23044
rect 42484 23004 43076 23032
rect 42484 22992 42490 23004
rect 43070 22992 43076 23004
rect 43128 22992 43134 23044
rect 39356 22936 39436 22964
rect 39356 22924 39362 22936
rect 39666 22924 39672 22976
rect 39724 22964 39730 22976
rect 39942 22964 39948 22976
rect 39724 22936 39948 22964
rect 39724 22924 39730 22936
rect 39942 22924 39948 22936
rect 40000 22964 40006 22976
rect 40957 22967 41015 22973
rect 40957 22964 40969 22967
rect 40000 22936 40969 22964
rect 40000 22924 40006 22936
rect 40957 22933 40969 22936
rect 41003 22933 41015 22967
rect 40957 22927 41015 22933
rect 1104 22874 43884 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 43884 22874
rect 1104 22800 43884 22822
rect 15470 22720 15476 22772
rect 15528 22760 15534 22772
rect 16022 22760 16028 22772
rect 15528 22732 16028 22760
rect 15528 22720 15534 22732
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 17405 22763 17463 22769
rect 17405 22729 17417 22763
rect 17451 22760 17463 22763
rect 18966 22760 18972 22772
rect 17451 22732 18972 22760
rect 17451 22729 17463 22732
rect 17405 22723 17463 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 19334 22720 19340 22772
rect 19392 22720 19398 22772
rect 21266 22720 21272 22772
rect 21324 22720 21330 22772
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 25041 22763 25099 22769
rect 25041 22760 25053 22763
rect 24544 22732 25053 22760
rect 24544 22720 24550 22732
rect 25041 22729 25053 22732
rect 25087 22729 25099 22763
rect 25041 22723 25099 22729
rect 25148 22732 27752 22760
rect 15933 22695 15991 22701
rect 15933 22661 15945 22695
rect 15979 22692 15991 22695
rect 17586 22692 17592 22704
rect 15979 22664 17592 22692
rect 15979 22661 15991 22664
rect 15933 22655 15991 22661
rect 17586 22652 17592 22664
rect 17644 22652 17650 22704
rect 18414 22652 18420 22704
rect 18472 22692 18478 22704
rect 18472 22664 18828 22692
rect 18472 22652 18478 22664
rect 13538 22633 13544 22636
rect 13532 22624 13544 22633
rect 13499 22596 13544 22624
rect 13532 22587 13544 22596
rect 13538 22584 13544 22587
rect 13596 22584 13602 22636
rect 18046 22624 18052 22636
rect 16224 22596 18052 22624
rect 13262 22516 13268 22568
rect 13320 22516 13326 22568
rect 16224 22565 16252 22596
rect 18046 22584 18052 22596
rect 18104 22584 18110 22636
rect 18506 22584 18512 22636
rect 18564 22633 18570 22636
rect 18800 22633 18828 22664
rect 19978 22652 19984 22704
rect 20036 22692 20042 22704
rect 22741 22695 22799 22701
rect 20036 22664 22094 22692
rect 20036 22652 20042 22664
rect 18564 22624 18576 22633
rect 18785 22627 18843 22633
rect 18564 22596 18609 22624
rect 18564 22587 18576 22596
rect 18785 22593 18797 22627
rect 18831 22624 18843 22627
rect 20806 22624 20812 22636
rect 18831 22596 20812 22624
rect 18831 22593 18843 22596
rect 18785 22587 18843 22593
rect 18564 22584 18570 22587
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22525 16267 22559
rect 16209 22519 16267 22525
rect 14366 22448 14372 22500
rect 14424 22488 14430 22500
rect 14918 22488 14924 22500
rect 14424 22460 14924 22488
rect 14424 22448 14430 22460
rect 14918 22448 14924 22460
rect 14976 22488 14982 22500
rect 16853 22491 16911 22497
rect 16853 22488 16865 22491
rect 14976 22460 16865 22488
rect 14976 22448 14982 22460
rect 16853 22457 16865 22460
rect 16899 22457 16911 22491
rect 16853 22451 16911 22457
rect 20165 22491 20223 22497
rect 20165 22457 20177 22491
rect 20211 22488 20223 22491
rect 20898 22488 20904 22500
rect 20211 22460 20904 22488
rect 20211 22457 20223 22460
rect 20165 22451 20223 22457
rect 20898 22448 20904 22460
rect 20956 22448 20962 22500
rect 22066 22488 22094 22664
rect 22741 22661 22753 22695
rect 22787 22692 22799 22695
rect 23569 22695 23627 22701
rect 23569 22692 23581 22695
rect 22787 22664 23581 22692
rect 22787 22661 22799 22664
rect 22741 22655 22799 22661
rect 23569 22661 23581 22664
rect 23615 22692 23627 22695
rect 25148 22692 25176 22732
rect 27614 22692 27620 22704
rect 23615 22664 25176 22692
rect 25240 22664 27620 22692
rect 23615 22661 23627 22664
rect 23569 22655 23627 22661
rect 22646 22584 22652 22636
rect 22704 22584 22710 22636
rect 25240 22633 25268 22664
rect 27614 22652 27620 22664
rect 27672 22652 27678 22704
rect 27724 22692 27752 22732
rect 28350 22720 28356 22772
rect 28408 22720 28414 22772
rect 29362 22720 29368 22772
rect 29420 22720 29426 22772
rect 29917 22763 29975 22769
rect 29917 22729 29929 22763
rect 29963 22760 29975 22763
rect 30282 22760 30288 22772
rect 29963 22732 30288 22760
rect 29963 22729 29975 22732
rect 29917 22723 29975 22729
rect 30282 22720 30288 22732
rect 30340 22720 30346 22772
rect 30374 22720 30380 22772
rect 30432 22720 30438 22772
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 30837 22763 30895 22769
rect 30837 22760 30849 22763
rect 30524 22732 30849 22760
rect 30524 22720 30530 22732
rect 30837 22729 30849 22732
rect 30883 22729 30895 22763
rect 30837 22723 30895 22729
rect 32214 22720 32220 22772
rect 32272 22760 32278 22772
rect 32490 22760 32496 22772
rect 32272 22732 32496 22760
rect 32272 22720 32278 22732
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 32677 22763 32735 22769
rect 32677 22729 32689 22763
rect 32723 22760 32735 22763
rect 33410 22760 33416 22772
rect 32723 22732 33416 22760
rect 32723 22729 32735 22732
rect 32677 22723 32735 22729
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 34054 22760 34060 22772
rect 33704 22732 34060 22760
rect 30098 22692 30104 22704
rect 27724 22664 30104 22692
rect 30098 22652 30104 22664
rect 30156 22652 30162 22704
rect 31294 22692 31300 22704
rect 30208 22664 31300 22692
rect 25225 22627 25283 22633
rect 25225 22593 25237 22627
rect 25271 22593 25283 22627
rect 25225 22587 25283 22593
rect 25406 22584 25412 22636
rect 25464 22584 25470 22636
rect 27246 22584 27252 22636
rect 27304 22624 27310 22636
rect 28166 22624 28172 22636
rect 27304 22596 28172 22624
rect 27304 22584 27310 22596
rect 28166 22584 28172 22596
rect 28224 22624 28230 22636
rect 30208 22624 30236 22664
rect 31294 22652 31300 22664
rect 31352 22652 31358 22704
rect 32585 22695 32643 22701
rect 32585 22661 32597 22695
rect 32631 22692 32643 22695
rect 32950 22692 32956 22704
rect 32631 22664 32956 22692
rect 32631 22661 32643 22664
rect 32585 22655 32643 22661
rect 32950 22652 32956 22664
rect 33008 22692 33014 22704
rect 33321 22695 33379 22701
rect 33321 22692 33333 22695
rect 33008 22664 33333 22692
rect 33008 22652 33014 22664
rect 33321 22661 33333 22664
rect 33367 22661 33379 22695
rect 33321 22655 33379 22661
rect 28224 22596 30236 22624
rect 28224 22584 28230 22596
rect 30742 22584 30748 22636
rect 30800 22584 30806 22636
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33704 22633 33732 22732
rect 34054 22720 34060 22732
rect 34112 22760 34118 22772
rect 34330 22760 34336 22772
rect 34112 22732 34336 22760
rect 34112 22720 34118 22732
rect 34330 22720 34336 22732
rect 34388 22720 34394 22772
rect 34701 22763 34759 22769
rect 34701 22729 34713 22763
rect 34747 22760 34759 22763
rect 34790 22760 34796 22772
rect 34747 22732 34796 22760
rect 34747 22729 34759 22732
rect 34701 22723 34759 22729
rect 34790 22720 34796 22732
rect 34848 22720 34854 22772
rect 34882 22720 34888 22772
rect 34940 22760 34946 22772
rect 34940 22732 36768 22760
rect 34940 22720 34946 22732
rect 33778 22652 33784 22704
rect 33836 22692 33842 22704
rect 33962 22692 33968 22704
rect 33836 22664 33968 22692
rect 33836 22652 33842 22664
rect 33962 22652 33968 22664
rect 34020 22692 34026 22704
rect 36740 22692 36768 22732
rect 36814 22720 36820 22772
rect 36872 22720 36878 22772
rect 37918 22720 37924 22772
rect 37976 22760 37982 22772
rect 38378 22760 38384 22772
rect 37976 22732 38384 22760
rect 37976 22720 37982 22732
rect 38378 22720 38384 22732
rect 38436 22720 38442 22772
rect 38930 22720 38936 22772
rect 38988 22760 38994 22772
rect 39117 22763 39175 22769
rect 39117 22760 39129 22763
rect 38988 22732 39129 22760
rect 38988 22720 38994 22732
rect 39117 22729 39129 22732
rect 39163 22760 39175 22763
rect 39482 22760 39488 22772
rect 39163 22732 39488 22760
rect 39163 22729 39175 22732
rect 39117 22723 39175 22729
rect 39482 22720 39488 22732
rect 39540 22720 39546 22772
rect 42334 22720 42340 22772
rect 42392 22760 42398 22772
rect 43257 22763 43315 22769
rect 43257 22760 43269 22763
rect 42392 22732 43269 22760
rect 42392 22720 42398 22732
rect 43257 22729 43269 22732
rect 43303 22729 43315 22763
rect 43257 22723 43315 22729
rect 39666 22692 39672 22704
rect 34020 22664 34100 22692
rect 36740 22664 39672 22692
rect 34020 22652 34026 22664
rect 34072 22633 34100 22664
rect 39666 22652 39672 22664
rect 39724 22652 39730 22704
rect 41782 22652 41788 22704
rect 41840 22692 41846 22704
rect 42058 22692 42064 22704
rect 41840 22664 42064 22692
rect 41840 22652 41846 22664
rect 42058 22652 42064 22664
rect 42116 22692 42122 22704
rect 42613 22695 42671 22701
rect 42613 22692 42625 22695
rect 42116 22664 42625 22692
rect 42116 22652 42122 22664
rect 42613 22661 42625 22664
rect 42659 22661 42671 22695
rect 42613 22655 42671 22661
rect 33413 22627 33471 22633
rect 33413 22624 33425 22627
rect 33192 22596 33425 22624
rect 33192 22584 33198 22596
rect 33413 22593 33425 22596
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 33873 22627 33931 22633
rect 33873 22593 33885 22627
rect 33919 22593 33931 22627
rect 33873 22587 33931 22593
rect 34057 22627 34115 22633
rect 34057 22593 34069 22627
rect 34103 22593 34115 22627
rect 34057 22587 34115 22593
rect 22922 22516 22928 22568
rect 22980 22516 22986 22568
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25961 22559 26019 22565
rect 25961 22556 25973 22559
rect 24912 22528 25973 22556
rect 24912 22516 24918 22528
rect 25961 22525 25973 22528
rect 26007 22556 26019 22559
rect 26007 22528 30972 22556
rect 26007 22525 26019 22528
rect 25961 22519 26019 22525
rect 25682 22488 25688 22500
rect 22066 22460 25688 22488
rect 25682 22448 25688 22460
rect 25740 22488 25746 22500
rect 26326 22488 26332 22500
rect 25740 22460 26332 22488
rect 25740 22448 25746 22460
rect 26326 22448 26332 22460
rect 26384 22448 26390 22500
rect 27798 22448 27804 22500
rect 27856 22488 27862 22500
rect 28810 22488 28816 22500
rect 27856 22460 28816 22488
rect 27856 22448 27862 22460
rect 28810 22448 28816 22460
rect 28868 22448 28874 22500
rect 30944 22488 30972 22528
rect 31018 22516 31024 22568
rect 31076 22516 31082 22568
rect 30944 22460 31754 22488
rect 14458 22380 14464 22432
rect 14516 22420 14522 22432
rect 14645 22423 14703 22429
rect 14645 22420 14657 22423
rect 14516 22392 14657 22420
rect 14516 22380 14522 22392
rect 14645 22389 14657 22392
rect 14691 22389 14703 22423
rect 14645 22383 14703 22389
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15252 22392 15577 22420
rect 15252 22380 15258 22392
rect 15565 22389 15577 22392
rect 15611 22389 15623 22423
rect 15565 22383 15623 22389
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 22281 22423 22339 22429
rect 22281 22389 22293 22423
rect 22327 22420 22339 22423
rect 22370 22420 22376 22432
rect 22327 22392 22376 22420
rect 22327 22389 22339 22392
rect 22281 22383 22339 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 22646 22380 22652 22432
rect 22704 22420 22710 22432
rect 24121 22423 24179 22429
rect 24121 22420 24133 22423
rect 22704 22392 24133 22420
rect 22704 22380 22710 22392
rect 24121 22389 24133 22392
rect 24167 22420 24179 22423
rect 26605 22423 26663 22429
rect 26605 22420 26617 22423
rect 24167 22392 26617 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 26605 22389 26617 22392
rect 26651 22420 26663 22423
rect 26878 22420 26884 22432
rect 26651 22392 26884 22420
rect 26651 22389 26663 22392
rect 26605 22383 26663 22389
rect 26878 22380 26884 22392
rect 26936 22420 26942 22432
rect 30466 22420 30472 22432
rect 26936 22392 30472 22420
rect 26936 22380 26942 22392
rect 30466 22380 30472 22392
rect 30524 22380 30530 22432
rect 31570 22380 31576 22432
rect 31628 22380 31634 22432
rect 31726 22420 31754 22460
rect 32306 22448 32312 22500
rect 32364 22448 32370 22500
rect 32784 22460 33548 22488
rect 32784 22420 32812 22460
rect 31726 22392 32812 22420
rect 32858 22380 32864 22432
rect 32916 22380 32922 22432
rect 33520 22420 33548 22460
rect 33594 22448 33600 22500
rect 33652 22488 33658 22500
rect 33879 22488 33907 22587
rect 35618 22584 35624 22636
rect 35676 22584 35682 22636
rect 35894 22584 35900 22636
rect 35952 22584 35958 22636
rect 36078 22584 36084 22636
rect 36136 22584 36142 22636
rect 36630 22584 36636 22636
rect 36688 22584 36694 22636
rect 36814 22584 36820 22636
rect 36872 22584 36878 22636
rect 36998 22584 37004 22636
rect 37056 22624 37062 22636
rect 37461 22627 37519 22633
rect 37461 22624 37473 22627
rect 37056 22596 37473 22624
rect 37056 22584 37062 22596
rect 37461 22593 37473 22596
rect 37507 22593 37519 22627
rect 37461 22587 37519 22593
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37918 22624 37924 22636
rect 37608 22596 37924 22624
rect 37608 22584 37614 22596
rect 37918 22584 37924 22596
rect 37976 22584 37982 22636
rect 38194 22584 38200 22636
rect 38252 22624 38258 22636
rect 39025 22627 39083 22633
rect 39025 22624 39037 22627
rect 38252 22596 39037 22624
rect 38252 22584 38258 22596
rect 39025 22593 39037 22596
rect 39071 22593 39083 22627
rect 39025 22587 39083 22593
rect 39206 22584 39212 22636
rect 39264 22624 39270 22636
rect 39390 22624 39396 22636
rect 39264 22596 39396 22624
rect 39264 22584 39270 22596
rect 39390 22584 39396 22596
rect 39448 22584 39454 22636
rect 40862 22584 40868 22636
rect 40920 22584 40926 22636
rect 41877 22627 41935 22633
rect 41877 22593 41889 22627
rect 41923 22624 41935 22627
rect 42242 22624 42248 22636
rect 41923 22596 42248 22624
rect 41923 22593 41935 22596
rect 41877 22587 41935 22593
rect 42242 22584 42248 22596
rect 42300 22584 42306 22636
rect 43070 22584 43076 22636
rect 43128 22624 43134 22636
rect 43254 22624 43260 22636
rect 43128 22596 43260 22624
rect 43128 22584 43134 22596
rect 43254 22584 43260 22596
rect 43312 22584 43318 22636
rect 35802 22516 35808 22568
rect 35860 22556 35866 22568
rect 39669 22559 39727 22565
rect 39669 22556 39681 22559
rect 35860 22528 39681 22556
rect 35860 22516 35866 22528
rect 39669 22525 39681 22528
rect 39715 22525 39727 22559
rect 39669 22519 39727 22525
rect 42978 22516 42984 22568
rect 43036 22516 43042 22568
rect 38838 22488 38844 22500
rect 33652 22460 38844 22488
rect 33652 22448 33658 22460
rect 38838 22448 38844 22460
rect 38896 22448 38902 22500
rect 39298 22448 39304 22500
rect 39356 22488 39362 22500
rect 39482 22488 39488 22500
rect 39356 22460 39488 22488
rect 39356 22448 39362 22460
rect 39482 22448 39488 22460
rect 39540 22448 39546 22500
rect 40402 22488 40408 22500
rect 39960 22460 40408 22488
rect 34882 22420 34888 22432
rect 33520 22392 34888 22420
rect 34882 22380 34888 22392
rect 34940 22380 34946 22432
rect 34974 22380 34980 22432
rect 35032 22420 35038 22432
rect 35759 22423 35817 22429
rect 35759 22420 35771 22423
rect 35032 22392 35771 22420
rect 35032 22380 35038 22392
rect 35759 22389 35771 22392
rect 35805 22420 35817 22423
rect 35894 22420 35900 22432
rect 35805 22392 35900 22420
rect 35805 22389 35817 22392
rect 35759 22383 35817 22389
rect 35894 22380 35900 22392
rect 35952 22380 35958 22432
rect 35986 22380 35992 22432
rect 36044 22380 36050 22432
rect 36538 22380 36544 22432
rect 36596 22420 36602 22432
rect 37553 22423 37611 22429
rect 37553 22420 37565 22423
rect 36596 22392 37565 22420
rect 36596 22380 36602 22392
rect 37553 22389 37565 22392
rect 37599 22389 37611 22423
rect 37553 22383 37611 22389
rect 38197 22423 38255 22429
rect 38197 22389 38209 22423
rect 38243 22420 38255 22423
rect 39022 22420 39028 22432
rect 38243 22392 39028 22420
rect 38243 22389 38255 22392
rect 38197 22383 38255 22389
rect 39022 22380 39028 22392
rect 39080 22420 39086 22432
rect 39960 22420 39988 22460
rect 40402 22448 40408 22460
rect 40460 22448 40466 22500
rect 39080 22392 39988 22420
rect 39080 22380 39086 22392
rect 40034 22380 40040 22432
rect 40092 22420 40098 22432
rect 40221 22423 40279 22429
rect 40221 22420 40233 22423
rect 40092 22392 40233 22420
rect 40092 22380 40098 22392
rect 40221 22389 40233 22392
rect 40267 22389 40279 22423
rect 40221 22383 40279 22389
rect 41049 22423 41107 22429
rect 41049 22389 41061 22423
rect 41095 22420 41107 22423
rect 41782 22420 41788 22432
rect 41095 22392 41788 22420
rect 41095 22389 41107 22392
rect 41049 22383 41107 22389
rect 41782 22380 41788 22392
rect 41840 22380 41846 22432
rect 41969 22423 42027 22429
rect 41969 22389 41981 22423
rect 42015 22420 42027 22423
rect 42150 22420 42156 22432
rect 42015 22392 42156 22420
rect 42015 22389 42027 22392
rect 41969 22383 42027 22389
rect 42150 22380 42156 22392
rect 42208 22380 42214 22432
rect 42702 22380 42708 22432
rect 42760 22380 42766 22432
rect 1104 22330 43884 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 43884 22330
rect 1104 22256 43884 22278
rect 14274 22176 14280 22228
rect 14332 22176 14338 22228
rect 15470 22176 15476 22228
rect 15528 22176 15534 22228
rect 15838 22216 15844 22228
rect 15580 22188 15844 22216
rect 14366 22148 14372 22160
rect 13556 22120 14372 22148
rect 13556 22089 13584 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 15488 22148 15516 22176
rect 14660 22120 15516 22148
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 14660 22080 14688 22120
rect 13587 22052 13621 22080
rect 13740 22052 14688 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 13449 22015 13507 22021
rect 12391 21984 12756 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12526 21836 12532 21888
rect 12584 21836 12590 21888
rect 12728 21876 12756 21984
rect 13449 21981 13461 22015
rect 13495 22012 13507 22015
rect 13740 22012 13768 22052
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 14918 22040 14924 22092
rect 14976 22040 14982 22092
rect 15580 22089 15608 22188
rect 15838 22176 15844 22188
rect 15896 22216 15902 22228
rect 15896 22188 18736 22216
rect 15896 22176 15902 22188
rect 16945 22151 17003 22157
rect 16945 22117 16957 22151
rect 16991 22148 17003 22151
rect 17586 22148 17592 22160
rect 16991 22120 17592 22148
rect 16991 22117 17003 22120
rect 16945 22111 17003 22117
rect 17586 22108 17592 22120
rect 17644 22108 17650 22160
rect 18598 22108 18604 22160
rect 18656 22108 18662 22160
rect 18708 22148 18736 22188
rect 19334 22176 19340 22228
rect 19392 22216 19398 22228
rect 19705 22219 19763 22225
rect 19705 22216 19717 22219
rect 19392 22188 19717 22216
rect 19392 22176 19398 22188
rect 19705 22185 19717 22188
rect 19751 22185 19763 22219
rect 19705 22179 19763 22185
rect 22002 22176 22008 22228
rect 22060 22176 22066 22228
rect 24854 22176 24860 22228
rect 24912 22216 24918 22228
rect 24912 22188 28304 22216
rect 24912 22176 24918 22188
rect 22020 22148 22048 22176
rect 23750 22148 23756 22160
rect 18708 22120 20484 22148
rect 22020 22120 23756 22148
rect 15565 22083 15623 22089
rect 15565 22049 15577 22083
rect 15611 22049 15623 22083
rect 15565 22043 15623 22049
rect 18046 22040 18052 22092
rect 18104 22040 18110 22092
rect 18138 22040 18144 22092
rect 18196 22040 18202 22092
rect 20456 22089 20484 22120
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20487 22052 20521 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 21910 22080 21916 22092
rect 20864 22052 21916 22080
rect 20864 22040 20870 22052
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 13495 21984 13768 22012
rect 13495 21981 13507 21984
rect 13449 21975 13507 21981
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14516 21984 14657 22012
rect 14516 21972 14522 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 22012 18291 22015
rect 18966 22012 18972 22024
rect 18279 21984 18972 22012
rect 18279 21981 18291 21984
rect 18233 21975 18291 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 21269 22015 21327 22021
rect 21269 22012 21281 22015
rect 20772 21984 21281 22012
rect 20772 21972 20778 21984
rect 21269 21981 21281 21984
rect 21315 21981 21327 22015
rect 21269 21975 21327 21981
rect 15378 21904 15384 21956
rect 15436 21944 15442 21956
rect 15810 21947 15868 21953
rect 15810 21944 15822 21947
rect 15436 21916 15822 21944
rect 15436 21904 15442 21916
rect 15810 21913 15822 21916
rect 15856 21913 15868 21947
rect 15810 21907 15868 21913
rect 19889 21947 19947 21953
rect 19889 21913 19901 21947
rect 19935 21944 19947 21947
rect 20254 21944 20260 21956
rect 19935 21916 20260 21944
rect 19935 21913 19947 21916
rect 19889 21907 19947 21913
rect 20254 21904 20260 21916
rect 20312 21904 20318 21956
rect 21284 21944 21312 21975
rect 22094 21972 22100 22024
rect 22152 21972 22158 22024
rect 23584 22012 23612 22120
rect 23750 22108 23756 22120
rect 23808 22108 23814 22160
rect 28276 22148 28304 22188
rect 28902 22176 28908 22228
rect 28960 22216 28966 22228
rect 28960 22188 30696 22216
rect 28960 22176 28966 22188
rect 28994 22148 29000 22160
rect 28276 22120 29000 22148
rect 28994 22108 29000 22120
rect 29052 22108 29058 22160
rect 29730 22108 29736 22160
rect 29788 22108 29794 22160
rect 23661 22015 23719 22021
rect 23661 22012 23673 22015
rect 23584 21984 23673 22012
rect 23661 21981 23673 21984
rect 23707 22012 23719 22015
rect 24578 22012 24584 22024
rect 23707 21984 24584 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 26786 21972 26792 22024
rect 26844 22012 26850 22024
rect 26881 22015 26939 22021
rect 26881 22012 26893 22015
rect 26844 21984 26893 22012
rect 26844 21972 26850 21984
rect 26881 21981 26893 21984
rect 26927 22012 26939 22015
rect 27341 22015 27399 22021
rect 27341 22012 27353 22015
rect 26927 21984 27353 22012
rect 26927 21981 26939 21984
rect 26881 21975 26939 21981
rect 27341 21981 27353 21984
rect 27387 22012 27399 22015
rect 28534 22012 28540 22024
rect 27387 21984 28540 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 29886 22021 29914 22188
rect 30668 22148 30696 22188
rect 30742 22176 30748 22228
rect 30800 22216 30806 22228
rect 30837 22219 30895 22225
rect 30837 22216 30849 22219
rect 30800 22188 30849 22216
rect 30800 22176 30806 22188
rect 30837 22185 30849 22188
rect 30883 22185 30895 22219
rect 30837 22179 30895 22185
rect 34790 22176 34796 22228
rect 34848 22216 34854 22228
rect 35069 22219 35127 22225
rect 35069 22216 35081 22219
rect 34848 22188 35081 22216
rect 34848 22176 34854 22188
rect 35069 22185 35081 22188
rect 35115 22216 35127 22219
rect 35158 22216 35164 22228
rect 35115 22188 35164 22216
rect 35115 22185 35127 22188
rect 35069 22179 35127 22185
rect 35158 22176 35164 22188
rect 35216 22176 35222 22228
rect 35434 22176 35440 22228
rect 35492 22216 35498 22228
rect 37645 22219 37703 22225
rect 37645 22216 37657 22219
rect 35492 22188 37657 22216
rect 35492 22176 35498 22188
rect 37645 22185 37657 22188
rect 37691 22216 37703 22219
rect 39022 22216 39028 22228
rect 37691 22188 39028 22216
rect 37691 22185 37703 22188
rect 37645 22179 37703 22185
rect 39022 22176 39028 22188
rect 39080 22176 39086 22228
rect 39298 22176 39304 22228
rect 39356 22216 39362 22228
rect 42518 22216 42524 22228
rect 39356 22188 42524 22216
rect 39356 22176 39362 22188
rect 42518 22176 42524 22188
rect 42576 22176 42582 22228
rect 42978 22176 42984 22228
rect 43036 22216 43042 22228
rect 43211 22219 43269 22225
rect 43211 22216 43223 22219
rect 43036 22188 43223 22216
rect 43036 22176 43042 22188
rect 43211 22185 43223 22188
rect 43257 22185 43269 22219
rect 43211 22179 43269 22185
rect 31570 22148 31576 22160
rect 30668 22120 31576 22148
rect 31570 22108 31576 22120
rect 31628 22108 31634 22160
rect 32030 22108 32036 22160
rect 32088 22108 32094 22160
rect 35802 22108 35808 22160
rect 35860 22148 35866 22160
rect 35860 22120 36032 22148
rect 35860 22108 35866 22120
rect 30098 22040 30104 22092
rect 30156 22040 30162 22092
rect 33870 22040 33876 22092
rect 33928 22040 33934 22092
rect 35618 22040 35624 22092
rect 35676 22080 35682 22092
rect 36004 22080 36032 22120
rect 36446 22108 36452 22160
rect 36504 22148 36510 22160
rect 39942 22148 39948 22160
rect 36504 22120 39948 22148
rect 36504 22108 36510 22120
rect 35676 22052 36032 22080
rect 35676 22040 35682 22052
rect 36078 22040 36084 22092
rect 36136 22080 36142 22092
rect 36173 22083 36231 22089
rect 36173 22080 36185 22083
rect 36136 22052 36185 22080
rect 36136 22040 36142 22052
rect 36173 22049 36185 22052
rect 36219 22049 36231 22083
rect 36173 22043 36231 22049
rect 36538 22040 36544 22092
rect 36596 22040 36602 22092
rect 29871 22015 29929 22021
rect 29871 21981 29883 22015
rect 29917 21981 29929 22015
rect 30116 22012 30144 22040
rect 29871 21975 29929 21981
rect 30024 21984 30144 22012
rect 30285 22015 30343 22021
rect 22833 21947 22891 21953
rect 22833 21944 22845 21947
rect 21284 21916 22845 21944
rect 22833 21913 22845 21916
rect 22879 21944 22891 21947
rect 23842 21944 23848 21956
rect 22879 21916 23848 21944
rect 22879 21913 22891 21916
rect 22833 21907 22891 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 24848 21947 24906 21953
rect 24848 21913 24860 21947
rect 24894 21944 24906 21947
rect 25406 21944 25412 21956
rect 24894 21916 25412 21944
rect 24894 21913 24906 21916
rect 24848 21907 24906 21913
rect 25406 21904 25412 21916
rect 25464 21904 25470 21956
rect 27608 21947 27666 21953
rect 27608 21913 27620 21947
rect 27654 21944 27666 21947
rect 28074 21944 28080 21956
rect 27654 21916 28080 21944
rect 27654 21913 27666 21916
rect 27608 21907 27666 21913
rect 28074 21904 28080 21916
rect 28132 21904 28138 21956
rect 28902 21904 28908 21956
rect 28960 21944 28966 21956
rect 30024 21953 30052 21984
rect 30285 21981 30297 22015
rect 30331 21981 30343 22015
rect 30285 21975 30343 21981
rect 30009 21947 30067 21953
rect 28960 21904 28994 21944
rect 30009 21913 30021 21947
rect 30055 21913 30067 21947
rect 30009 21907 30067 21913
rect 30101 21947 30159 21953
rect 30101 21913 30113 21947
rect 30147 21944 30159 21947
rect 30190 21944 30196 21956
rect 30147 21916 30196 21944
rect 30147 21913 30159 21916
rect 30101 21907 30159 21913
rect 30190 21904 30196 21916
rect 30248 21904 30254 21956
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 12728 21848 13001 21876
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 12989 21839 13047 21845
rect 13357 21879 13415 21885
rect 13357 21845 13369 21879
rect 13403 21876 13415 21879
rect 14734 21876 14740 21888
rect 13403 21848 14740 21876
rect 13403 21845 13415 21848
rect 13357 21839 13415 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 19484 21848 19533 21876
rect 19484 21836 19490 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 19521 21839 19579 21845
rect 19689 21879 19747 21885
rect 19689 21845 19701 21879
rect 19735 21876 19747 21879
rect 19978 21876 19984 21888
rect 19735 21848 19984 21876
rect 19735 21845 19747 21848
rect 19689 21839 19747 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 25682 21876 25688 21888
rect 23072 21848 25688 21876
rect 23072 21836 23078 21848
rect 25682 21836 25688 21848
rect 25740 21876 25746 21888
rect 25961 21879 26019 21885
rect 25961 21876 25973 21879
rect 25740 21848 25973 21876
rect 25740 21836 25746 21848
rect 25961 21845 25973 21848
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 28718 21836 28724 21888
rect 28776 21836 28782 21888
rect 28966 21876 28994 21904
rect 30300 21876 30328 21975
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 31110 22012 31116 22024
rect 30984 21984 31116 22012
rect 30984 21972 30990 21984
rect 31110 21972 31116 21984
rect 31168 21972 31174 22024
rect 31757 22015 31815 22021
rect 31757 21981 31769 22015
rect 31803 22012 31815 22015
rect 32030 22012 32036 22024
rect 31803 21984 32036 22012
rect 31803 21981 31815 21984
rect 31757 21975 31815 21981
rect 32030 21972 32036 21984
rect 32088 21972 32094 22024
rect 32490 21972 32496 22024
rect 32548 21972 32554 22024
rect 32950 21972 32956 22024
rect 33008 21972 33014 22024
rect 33410 21972 33416 22024
rect 33468 21972 33474 22024
rect 36354 21972 36360 22024
rect 36412 21972 36418 22024
rect 36630 21972 36636 22024
rect 36688 21972 36694 22024
rect 36740 22021 36768 22120
rect 39942 22108 39948 22120
rect 40000 22108 40006 22160
rect 38194 22040 38200 22092
rect 38252 22080 38258 22092
rect 38252 22052 38792 22080
rect 38252 22040 38258 22052
rect 36725 22015 36783 22021
rect 36725 21981 36737 22015
rect 36771 21981 36783 22015
rect 36725 21975 36783 21981
rect 36909 22015 36967 22021
rect 36909 21981 36921 22015
rect 36955 22012 36967 22015
rect 37182 22012 37188 22024
rect 36955 21984 37188 22012
rect 36955 21981 36967 21984
rect 36909 21975 36967 21981
rect 37182 21972 37188 21984
rect 37240 21972 37246 22024
rect 37458 21972 37464 22024
rect 37516 22012 37522 22024
rect 37645 22015 37703 22021
rect 37645 22012 37657 22015
rect 37516 21984 37657 22012
rect 37516 21972 37522 21984
rect 37645 21981 37657 21984
rect 37691 21981 37703 22015
rect 37645 21975 37703 21981
rect 37829 22015 37887 22021
rect 37829 21981 37841 22015
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 37921 22015 37979 22021
rect 37921 21981 37933 22015
rect 37967 22012 37979 22015
rect 38010 22012 38016 22024
rect 37967 21984 38016 22012
rect 37967 21981 37979 21984
rect 37921 21975 37979 21981
rect 34977 21947 35035 21953
rect 34977 21913 34989 21947
rect 35023 21913 35035 21947
rect 34977 21907 35035 21913
rect 28966 21848 30328 21876
rect 31386 21836 31392 21888
rect 31444 21876 31450 21888
rect 31662 21876 31668 21888
rect 31444 21848 31668 21876
rect 31444 21836 31450 21848
rect 31662 21836 31668 21848
rect 31720 21836 31726 21888
rect 34330 21836 34336 21888
rect 34388 21876 34394 21888
rect 34992 21876 35020 21907
rect 36078 21904 36084 21956
rect 36136 21944 36142 21956
rect 37734 21944 37740 21956
rect 36136 21916 37740 21944
rect 36136 21904 36142 21916
rect 37734 21904 37740 21916
rect 37792 21944 37798 21956
rect 37844 21944 37872 21975
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 38562 21972 38568 22024
rect 38620 21972 38626 22024
rect 38764 22021 38792 22052
rect 39114 22040 39120 22092
rect 39172 22080 39178 22092
rect 39172 22052 40080 22080
rect 39172 22040 39178 22052
rect 38749 22015 38807 22021
rect 38749 21981 38761 22015
rect 38795 21981 38807 22015
rect 38749 21975 38807 21981
rect 38838 21972 38844 22024
rect 38896 22012 38902 22024
rect 40052 22021 40080 22052
rect 40310 22040 40316 22092
rect 40368 22080 40374 22092
rect 41417 22083 41475 22089
rect 41417 22080 41429 22083
rect 40368 22052 41429 22080
rect 40368 22040 40374 22052
rect 41417 22049 41429 22052
rect 41463 22049 41475 22083
rect 41417 22043 41475 22049
rect 41782 22040 41788 22092
rect 41840 22040 41846 22092
rect 40037 22015 40095 22021
rect 38896 21984 39436 22012
rect 38896 21972 38902 21984
rect 38657 21947 38715 21953
rect 37792 21916 37872 21944
rect 37917 21916 38240 21944
rect 37792 21904 37798 21916
rect 37917 21876 37945 21916
rect 34388 21848 37945 21876
rect 34388 21836 34394 21848
rect 38102 21836 38108 21888
rect 38160 21836 38166 21888
rect 38212 21876 38240 21916
rect 38657 21913 38669 21947
rect 38703 21944 38715 21947
rect 39114 21944 39120 21956
rect 38703 21916 39120 21944
rect 38703 21913 38715 21916
rect 38657 21907 38715 21913
rect 39114 21904 39120 21916
rect 39172 21904 39178 21956
rect 39408 21944 39436 21984
rect 40037 21981 40049 22015
rect 40083 21981 40095 22015
rect 40037 21975 40095 21981
rect 40218 21972 40224 22024
rect 40276 21972 40282 22024
rect 40865 22015 40923 22021
rect 40865 21981 40877 22015
rect 40911 21981 40923 22015
rect 40865 21975 40923 21981
rect 40880 21944 40908 21975
rect 39408 21916 40908 21944
rect 42150 21904 42156 21956
rect 42208 21904 42214 21956
rect 39298 21876 39304 21888
rect 38212 21848 39304 21876
rect 39298 21836 39304 21848
rect 39356 21836 39362 21888
rect 39666 21836 39672 21888
rect 39724 21876 39730 21888
rect 40129 21879 40187 21885
rect 40129 21876 40141 21879
rect 39724 21848 40141 21876
rect 39724 21836 39730 21848
rect 40129 21845 40141 21848
rect 40175 21845 40187 21879
rect 40129 21839 40187 21845
rect 40678 21836 40684 21888
rect 40736 21836 40742 21888
rect 1104 21786 43884 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 43884 21786
rect 1104 21712 43884 21734
rect 14734 21632 14740 21684
rect 14792 21632 14798 21684
rect 15197 21675 15255 21681
rect 15197 21641 15209 21675
rect 15243 21672 15255 21675
rect 15286 21672 15292 21684
rect 15243 21644 15292 21672
rect 15243 21641 15255 21644
rect 15197 21635 15255 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 20809 21675 20867 21681
rect 20809 21641 20821 21675
rect 20855 21672 20867 21675
rect 20990 21672 20996 21684
rect 20855 21644 20996 21672
rect 20855 21641 20867 21644
rect 20809 21635 20867 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 22066 21644 22508 21672
rect 13262 21564 13268 21616
rect 13320 21604 13326 21616
rect 15838 21604 15844 21616
rect 13320 21576 15844 21604
rect 13320 21564 13326 21576
rect 13372 21545 13400 21576
rect 15838 21564 15844 21576
rect 15896 21564 15902 21616
rect 19426 21564 19432 21616
rect 19484 21604 19490 21616
rect 19613 21607 19671 21613
rect 19613 21604 19625 21607
rect 19484 21576 19625 21604
rect 19484 21564 19490 21576
rect 19613 21573 19625 21576
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 22066 21604 22094 21644
rect 22278 21613 22284 21616
rect 20956 21576 22094 21604
rect 20956 21564 20962 21576
rect 22272 21567 22284 21613
rect 22278 21564 22284 21567
rect 22336 21564 22342 21616
rect 22480 21604 22508 21644
rect 23842 21632 23848 21684
rect 23900 21632 23906 21684
rect 25498 21632 25504 21684
rect 25556 21672 25562 21684
rect 25685 21675 25743 21681
rect 25685 21672 25697 21675
rect 25556 21644 25697 21672
rect 25556 21632 25562 21644
rect 25685 21641 25697 21644
rect 25731 21641 25743 21675
rect 25685 21635 25743 21641
rect 25777 21675 25835 21681
rect 25777 21641 25789 21675
rect 25823 21672 25835 21675
rect 27157 21675 27215 21681
rect 27157 21672 27169 21675
rect 25823 21644 27169 21672
rect 25823 21641 25835 21644
rect 25777 21635 25835 21641
rect 27157 21641 27169 21644
rect 27203 21641 27215 21675
rect 27157 21635 27215 21641
rect 28074 21632 28080 21684
rect 28132 21672 28138 21684
rect 28902 21672 28908 21684
rect 28132 21644 28908 21672
rect 28132 21632 28138 21644
rect 28902 21632 28908 21644
rect 28960 21632 28966 21684
rect 29822 21632 29828 21684
rect 29880 21672 29886 21684
rect 29917 21675 29975 21681
rect 29917 21672 29929 21675
rect 29880 21644 29929 21672
rect 29880 21632 29886 21644
rect 29917 21641 29929 21644
rect 29963 21672 29975 21675
rect 30098 21672 30104 21684
rect 29963 21644 30104 21672
rect 29963 21641 29975 21644
rect 29917 21635 29975 21641
rect 30098 21632 30104 21644
rect 30156 21632 30162 21684
rect 34606 21672 34612 21684
rect 30760 21644 34612 21672
rect 28804 21607 28862 21613
rect 22480 21576 26648 21604
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13613 21539 13671 21545
rect 13613 21536 13625 21539
rect 13357 21499 13415 21505
rect 13464 21508 13625 21536
rect 12526 21428 12532 21480
rect 12584 21468 12590 21480
rect 13464 21468 13492 21508
rect 13613 21505 13625 21508
rect 13659 21505 13671 21539
rect 13613 21499 13671 21505
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 14792 21508 15393 21536
rect 14792 21496 14798 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 15746 21536 15752 21548
rect 15620 21508 15752 21536
rect 15620 21496 15626 21508
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 16298 21496 16304 21548
rect 16356 21496 16362 21548
rect 17126 21496 17132 21548
rect 17184 21496 17190 21548
rect 17862 21496 17868 21548
rect 17920 21496 17926 21548
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21536 18199 21539
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18187 21508 18705 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 12584 21440 13492 21468
rect 17972 21468 18000 21499
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 26620 21545 26648 21576
rect 28804 21573 28816 21607
rect 28850 21604 28862 21607
rect 29730 21604 29736 21616
rect 28850 21576 29736 21604
rect 28850 21573 28862 21576
rect 28804 21567 28862 21573
rect 29730 21564 29736 21576
rect 29788 21564 29794 21616
rect 30760 21613 30788 21644
rect 34606 21632 34612 21644
rect 34664 21632 34670 21684
rect 35989 21675 36047 21681
rect 35989 21641 36001 21675
rect 36035 21672 36047 21675
rect 36078 21672 36084 21684
rect 36035 21644 36084 21672
rect 36035 21641 36047 21644
rect 35989 21635 36047 21641
rect 36078 21632 36084 21644
rect 36136 21632 36142 21684
rect 38749 21675 38807 21681
rect 37844 21644 38700 21672
rect 30745 21607 30803 21613
rect 30745 21573 30757 21607
rect 30791 21573 30803 21607
rect 32398 21604 32404 21616
rect 30745 21567 30803 21573
rect 30852 21576 32404 21604
rect 24857 21539 24915 21545
rect 20036 21508 24808 21536
rect 20036 21496 20042 21508
rect 19996 21468 20024 21496
rect 17972 21440 20024 21468
rect 12584 21428 12590 21440
rect 21082 21428 21088 21480
rect 21140 21428 21146 21480
rect 22002 21428 22008 21480
rect 22060 21428 22066 21480
rect 18230 21360 18236 21412
rect 18288 21400 18294 21412
rect 20441 21403 20499 21409
rect 20441 21400 20453 21403
rect 18288 21372 20453 21400
rect 18288 21360 18294 21372
rect 20441 21369 20453 21372
rect 20487 21369 20499 21403
rect 20441 21363 20499 21369
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 17313 21335 17371 21341
rect 17313 21301 17325 21335
rect 17359 21332 17371 21335
rect 17494 21332 17500 21344
rect 17359 21304 17500 21332
rect 17359 21301 17371 21304
rect 17313 21295 17371 21301
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 18966 21332 18972 21344
rect 18104 21304 18972 21332
rect 18104 21292 18110 21304
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 19889 21335 19947 21341
rect 19889 21301 19901 21335
rect 19935 21332 19947 21335
rect 20346 21332 20352 21344
rect 19935 21304 20352 21332
rect 19935 21301 19947 21304
rect 19889 21295 19947 21301
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 23382 21292 23388 21344
rect 23440 21292 23446 21344
rect 24670 21292 24676 21344
rect 24728 21292 24734 21344
rect 24780 21332 24808 21508
rect 24857 21505 24869 21539
rect 24903 21536 24915 21539
rect 26605 21539 26663 21545
rect 24903 21508 25360 21536
rect 24903 21505 24915 21508
rect 24857 21499 24915 21505
rect 25332 21409 25360 21508
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26878 21536 26884 21548
rect 26651 21508 26884 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 26878 21496 26884 21508
rect 26936 21536 26942 21548
rect 27062 21536 27068 21548
rect 26936 21508 27068 21536
rect 26936 21496 26942 21508
rect 27062 21496 27068 21508
rect 27120 21536 27126 21548
rect 27525 21539 27583 21545
rect 27525 21536 27537 21539
rect 27120 21508 27537 21536
rect 27120 21496 27126 21508
rect 27525 21505 27537 21508
rect 27571 21505 27583 21539
rect 29362 21536 29368 21548
rect 27525 21499 27583 21505
rect 27816 21508 29368 21536
rect 25961 21471 26019 21477
rect 25961 21437 25973 21471
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 25317 21403 25375 21409
rect 25317 21369 25329 21403
rect 25363 21369 25375 21403
rect 25976 21400 26004 21431
rect 27614 21428 27620 21480
rect 27672 21428 27678 21480
rect 27816 21477 27844 21508
rect 29362 21496 29368 21508
rect 29420 21496 29426 21548
rect 30558 21496 30564 21548
rect 30616 21496 30622 21548
rect 30852 21545 30880 21576
rect 32398 21564 32404 21576
rect 32456 21564 32462 21616
rect 32692 21576 33548 21604
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21505 30895 21539
rect 30837 21499 30895 21505
rect 31018 21496 31024 21548
rect 31076 21536 31082 21548
rect 32692 21545 32720 21576
rect 31297 21539 31355 21545
rect 31297 21536 31309 21539
rect 31076 21508 31309 21536
rect 31076 21496 31082 21508
rect 31297 21505 31309 21508
rect 31343 21505 31355 21539
rect 31297 21499 31355 21505
rect 32677 21539 32735 21545
rect 32677 21505 32689 21539
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 32858 21496 32864 21548
rect 32916 21496 32922 21548
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21437 27859 21471
rect 27801 21431 27859 21437
rect 28534 21428 28540 21480
rect 28592 21428 28598 21480
rect 32953 21471 33011 21477
rect 32953 21468 32965 21471
rect 32692 21440 32965 21468
rect 32692 21412 32720 21440
rect 32953 21437 32965 21440
rect 32999 21437 33011 21471
rect 32953 21431 33011 21437
rect 33134 21428 33140 21480
rect 33192 21428 33198 21480
rect 33520 21468 33548 21576
rect 35710 21564 35716 21616
rect 35768 21564 35774 21616
rect 36906 21564 36912 21616
rect 36964 21604 36970 21616
rect 37461 21607 37519 21613
rect 37461 21604 37473 21607
rect 36964 21576 37473 21604
rect 36964 21564 36970 21576
rect 37461 21573 37473 21576
rect 37507 21573 37519 21607
rect 37461 21567 37519 21573
rect 33594 21496 33600 21548
rect 33652 21536 33658 21548
rect 33781 21539 33839 21545
rect 33652 21508 33732 21536
rect 33652 21496 33658 21508
rect 33704 21468 33732 21508
rect 33781 21505 33793 21539
rect 33827 21536 33839 21539
rect 33962 21536 33968 21548
rect 33827 21508 33968 21536
rect 33827 21505 33839 21508
rect 33781 21499 33839 21505
rect 33962 21496 33968 21508
rect 34020 21496 34026 21548
rect 34057 21539 34115 21545
rect 34057 21505 34069 21539
rect 34103 21536 34115 21539
rect 34790 21536 34796 21548
rect 34103 21508 34796 21536
rect 34103 21505 34115 21508
rect 34057 21499 34115 21505
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 35158 21496 35164 21548
rect 35216 21536 35222 21548
rect 35434 21536 35440 21548
rect 35216 21508 35440 21536
rect 35216 21496 35222 21508
rect 35434 21496 35440 21508
rect 35492 21496 35498 21548
rect 35621 21539 35679 21545
rect 35621 21505 35633 21539
rect 35667 21505 35679 21539
rect 35621 21499 35679 21505
rect 33873 21471 33931 21477
rect 33873 21468 33885 21471
rect 33520 21440 33640 21468
rect 33704 21440 33885 21468
rect 28166 21400 28172 21412
rect 25976 21372 28172 21400
rect 25317 21363 25375 21369
rect 28166 21360 28172 21372
rect 28224 21360 28230 21412
rect 30834 21360 30840 21412
rect 30892 21400 30898 21412
rect 31481 21403 31539 21409
rect 31481 21400 31493 21403
rect 30892 21372 31493 21400
rect 30892 21360 30898 21372
rect 31481 21369 31493 21372
rect 31527 21369 31539 21403
rect 31481 21363 31539 21369
rect 31570 21360 31576 21412
rect 31628 21400 31634 21412
rect 32401 21403 32459 21409
rect 32401 21400 32413 21403
rect 31628 21372 32413 21400
rect 31628 21360 31634 21372
rect 32401 21369 32413 21372
rect 32447 21369 32459 21403
rect 32401 21363 32459 21369
rect 32674 21360 32680 21412
rect 32732 21360 32738 21412
rect 32769 21403 32827 21409
rect 32769 21369 32781 21403
rect 32815 21400 32827 21403
rect 33502 21400 33508 21412
rect 32815 21372 33508 21400
rect 32815 21369 32827 21372
rect 32769 21363 32827 21369
rect 33502 21360 33508 21372
rect 33560 21360 33566 21412
rect 33612 21400 33640 21440
rect 33873 21437 33885 21440
rect 33919 21437 33931 21471
rect 35636 21468 35664 21499
rect 35802 21496 35808 21548
rect 35860 21496 35866 21548
rect 35986 21496 35992 21548
rect 36044 21536 36050 21548
rect 37737 21539 37795 21545
rect 37737 21536 37749 21539
rect 36044 21508 37749 21536
rect 36044 21496 36050 21508
rect 37737 21505 37749 21508
rect 37783 21505 37795 21539
rect 37737 21499 37795 21505
rect 35710 21468 35716 21480
rect 35636 21440 35716 21468
rect 33873 21431 33931 21437
rect 35710 21428 35716 21440
rect 35768 21428 35774 21480
rect 37366 21428 37372 21480
rect 37424 21468 37430 21480
rect 37553 21471 37611 21477
rect 37553 21468 37565 21471
rect 37424 21440 37565 21468
rect 37424 21428 37430 21440
rect 37553 21437 37565 21440
rect 37599 21437 37611 21471
rect 37553 21431 37611 21437
rect 33965 21403 34023 21409
rect 33965 21400 33977 21403
rect 33612 21372 33977 21400
rect 33965 21369 33977 21372
rect 34011 21400 34023 21403
rect 34054 21400 34060 21412
rect 34011 21372 34060 21400
rect 34011 21369 34023 21372
rect 33965 21363 34023 21369
rect 34054 21360 34060 21372
rect 34112 21360 34118 21412
rect 37844 21400 37872 21644
rect 38672 21604 38700 21644
rect 38749 21641 38761 21675
rect 38795 21672 38807 21675
rect 38838 21672 38844 21684
rect 38795 21644 38844 21672
rect 38795 21641 38807 21644
rect 38749 21635 38807 21641
rect 38838 21632 38844 21644
rect 38896 21632 38902 21684
rect 39853 21675 39911 21681
rect 39853 21641 39865 21675
rect 39899 21672 39911 21675
rect 40862 21672 40868 21684
rect 39899 21644 40868 21672
rect 39899 21641 39911 21644
rect 39853 21635 39911 21641
rect 40862 21632 40868 21644
rect 40920 21632 40926 21684
rect 42058 21632 42064 21684
rect 42116 21632 42122 21684
rect 43346 21632 43352 21684
rect 43404 21632 43410 21684
rect 40034 21604 40040 21616
rect 38672 21576 40040 21604
rect 40034 21564 40040 21576
rect 40092 21604 40098 21616
rect 40494 21604 40500 21616
rect 40092 21576 40500 21604
rect 40092 21564 40098 21576
rect 40494 21564 40500 21576
rect 40552 21564 40558 21616
rect 40589 21607 40647 21613
rect 40589 21573 40601 21607
rect 40635 21604 40647 21607
rect 40678 21604 40684 21616
rect 40635 21576 40684 21604
rect 40635 21573 40647 21576
rect 40589 21567 40647 21573
rect 40678 21564 40684 21576
rect 40736 21564 40742 21616
rect 42705 21607 42763 21613
rect 42705 21604 42717 21607
rect 41814 21576 42717 21604
rect 42705 21573 42717 21576
rect 42751 21573 42763 21607
rect 42705 21567 42763 21573
rect 38102 21496 38108 21548
rect 38160 21536 38166 21548
rect 38381 21539 38439 21545
rect 38381 21536 38393 21539
rect 38160 21508 38393 21536
rect 38160 21496 38166 21508
rect 38381 21505 38393 21508
rect 38427 21505 38439 21539
rect 38381 21499 38439 21505
rect 38746 21496 38752 21548
rect 38804 21536 38810 21548
rect 39209 21539 39267 21545
rect 39209 21536 39221 21539
rect 38804 21508 39221 21536
rect 38804 21496 38810 21508
rect 39209 21505 39221 21508
rect 39255 21505 39267 21539
rect 39209 21499 39267 21505
rect 39574 21496 39580 21548
rect 39632 21536 39638 21548
rect 39669 21539 39727 21545
rect 39669 21536 39681 21539
rect 39632 21508 39681 21536
rect 39632 21496 39638 21508
rect 39669 21505 39681 21508
rect 39715 21505 39727 21539
rect 39669 21499 39727 21505
rect 40310 21496 40316 21548
rect 40368 21496 40374 21548
rect 42242 21496 42248 21548
rect 42300 21536 42306 21548
rect 42797 21539 42855 21545
rect 42797 21536 42809 21539
rect 42300 21508 42809 21536
rect 42300 21496 42306 21508
rect 42797 21505 42809 21508
rect 42843 21505 42855 21539
rect 42797 21499 42855 21505
rect 38470 21428 38476 21480
rect 38528 21428 38534 21480
rect 39485 21471 39543 21477
rect 39485 21437 39497 21471
rect 39531 21437 39543 21471
rect 39485 21431 39543 21437
rect 37016 21372 37872 21400
rect 37921 21403 37979 21409
rect 37016 21344 37044 21372
rect 37921 21369 37933 21403
rect 37967 21400 37979 21403
rect 39500 21400 39528 21431
rect 37967 21372 39528 21400
rect 37967 21369 37979 21372
rect 37921 21363 37979 21369
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 24780 21304 30665 21332
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 30653 21295 30711 21301
rect 33042 21292 33048 21344
rect 33100 21332 33106 21344
rect 33597 21335 33655 21341
rect 33597 21332 33609 21335
rect 33100 21304 33609 21332
rect 33100 21292 33106 21304
rect 33597 21301 33609 21304
rect 33643 21301 33655 21335
rect 33597 21295 33655 21301
rect 34793 21335 34851 21341
rect 34793 21301 34805 21335
rect 34839 21332 34851 21335
rect 35526 21332 35532 21344
rect 34839 21304 35532 21332
rect 34839 21301 34851 21304
rect 34793 21295 34851 21301
rect 35526 21292 35532 21304
rect 35584 21292 35590 21344
rect 35618 21292 35624 21344
rect 35676 21332 35682 21344
rect 35894 21332 35900 21344
rect 35676 21304 35900 21332
rect 35676 21292 35682 21304
rect 35894 21292 35900 21304
rect 35952 21332 35958 21344
rect 36541 21335 36599 21341
rect 36541 21332 36553 21335
rect 35952 21304 36553 21332
rect 35952 21292 35958 21304
rect 36541 21301 36553 21304
rect 36587 21332 36599 21335
rect 36998 21332 37004 21344
rect 36587 21304 37004 21332
rect 36587 21301 36599 21304
rect 36541 21295 36599 21301
rect 36998 21292 37004 21304
rect 37056 21292 37062 21344
rect 37458 21292 37464 21344
rect 37516 21292 37522 21344
rect 38565 21335 38623 21341
rect 38565 21301 38577 21335
rect 38611 21332 38623 21335
rect 39206 21332 39212 21344
rect 38611 21304 39212 21332
rect 38611 21301 38623 21304
rect 38565 21295 38623 21301
rect 39206 21292 39212 21304
rect 39264 21292 39270 21344
rect 39666 21292 39672 21344
rect 39724 21292 39730 21344
rect 1104 21242 43884 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 43884 21242
rect 1104 21168 43884 21190
rect 15378 21088 15384 21140
rect 15436 21088 15442 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17773 21131 17831 21137
rect 17773 21128 17785 21131
rect 17184 21100 17785 21128
rect 17184 21088 17190 21100
rect 17773 21097 17785 21100
rect 17819 21097 17831 21131
rect 17773 21091 17831 21097
rect 22094 21088 22100 21140
rect 22152 21088 22158 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 24854 21128 24860 21140
rect 22336 21100 24860 21128
rect 22336 21088 22342 21100
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 25958 21128 25964 21140
rect 25556 21100 25964 21128
rect 25556 21088 25562 21100
rect 25958 21088 25964 21100
rect 26016 21088 26022 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 26421 21131 26479 21137
rect 26421 21128 26433 21131
rect 26384 21100 26433 21128
rect 26384 21088 26390 21100
rect 26421 21097 26433 21100
rect 26467 21097 26479 21131
rect 26421 21091 26479 21097
rect 26436 21060 26464 21091
rect 27614 21088 27620 21140
rect 27672 21128 27678 21140
rect 27709 21131 27767 21137
rect 27709 21128 27721 21131
rect 27672 21100 27721 21128
rect 27672 21088 27678 21100
rect 27709 21097 27721 21100
rect 27755 21097 27767 21131
rect 27709 21091 27767 21097
rect 28166 21088 28172 21140
rect 28224 21088 28230 21140
rect 28534 21088 28540 21140
rect 28592 21128 28598 21140
rect 29089 21131 29147 21137
rect 29089 21128 29101 21131
rect 28592 21100 29101 21128
rect 28592 21088 28598 21100
rect 29089 21097 29101 21100
rect 29135 21097 29147 21131
rect 32493 21131 32551 21137
rect 32493 21128 32505 21131
rect 29089 21091 29147 21097
rect 29196 21100 32505 21128
rect 21100 21032 22094 21060
rect 18230 20952 18236 21004
rect 18288 20952 18294 21004
rect 18322 20952 18328 21004
rect 18380 20992 18386 21004
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 18380 20964 18429 20992
rect 18380 20952 18386 20964
rect 18417 20961 18429 20964
rect 18463 20992 18475 20995
rect 18463 20964 19104 20992
rect 18463 20961 18475 20964
rect 18417 20955 18475 20961
rect 19076 20936 19104 20964
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 15838 20884 15844 20936
rect 15896 20884 15902 20936
rect 16114 20933 16120 20936
rect 16108 20924 16120 20933
rect 16075 20896 16120 20924
rect 16108 20887 16120 20896
rect 16114 20884 16120 20887
rect 16172 20884 16178 20936
rect 19058 20884 19064 20936
rect 19116 20924 19122 20936
rect 21100 20933 21128 21032
rect 22066 20992 22094 21032
rect 22296 21032 23704 21060
rect 26436 21032 27292 21060
rect 22296 20992 22324 21032
rect 22649 20995 22707 21001
rect 22649 20992 22661 20995
rect 22066 20964 22324 20992
rect 22388 20964 22661 20992
rect 21085 20927 21143 20933
rect 19116 20896 21036 20924
rect 19116 20884 19122 20896
rect 15102 20816 15108 20868
rect 15160 20856 15166 20868
rect 19889 20859 19947 20865
rect 19889 20856 19901 20859
rect 15160 20828 19901 20856
rect 15160 20816 15166 20828
rect 19889 20825 19901 20828
rect 19935 20825 19947 20859
rect 19889 20819 19947 20825
rect 20257 20859 20315 20865
rect 20257 20825 20269 20859
rect 20303 20856 20315 20859
rect 20438 20856 20444 20868
rect 20303 20828 20444 20856
rect 20303 20825 20315 20828
rect 20257 20819 20315 20825
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13872 20760 14289 20788
rect 13872 20748 13878 20760
rect 14277 20757 14289 20760
rect 14323 20788 14335 20791
rect 14366 20788 14372 20800
rect 14323 20760 14372 20788
rect 14323 20757 14335 20760
rect 14277 20751 14335 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 17221 20791 17279 20797
rect 17221 20788 17233 20791
rect 16632 20760 17233 20788
rect 16632 20748 16638 20760
rect 17221 20757 17233 20760
rect 17267 20788 17279 20791
rect 17770 20788 17776 20800
rect 17267 20760 17776 20788
rect 17267 20757 17279 20760
rect 17221 20751 17279 20757
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 18138 20748 18144 20800
rect 18196 20748 18202 20800
rect 20898 20748 20904 20800
rect 20956 20748 20962 20800
rect 21008 20788 21036 20896
rect 21085 20893 21097 20927
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 21269 20927 21327 20933
rect 21269 20893 21281 20927
rect 21315 20924 21327 20927
rect 22278 20924 22284 20936
rect 21315 20896 22284 20924
rect 21315 20893 21327 20896
rect 21269 20887 21327 20893
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22388 20788 22416 20964
rect 22649 20961 22661 20964
rect 22695 20961 22707 20995
rect 22649 20955 22707 20961
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 22738 20924 22744 20936
rect 22511 20896 22744 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 22738 20884 22744 20896
rect 22796 20924 22802 20936
rect 23382 20924 23388 20936
rect 22796 20896 23388 20924
rect 22796 20884 22802 20896
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 23474 20884 23480 20936
rect 23532 20884 23538 20936
rect 23566 20884 23572 20936
rect 23624 20884 23630 20936
rect 22554 20816 22560 20868
rect 22612 20816 22618 20868
rect 21008 20760 22416 20788
rect 23676 20788 23704 21032
rect 24578 20952 24584 21004
rect 24636 20952 24642 21004
rect 27264 21001 27292 21032
rect 27157 20995 27215 21001
rect 27157 20961 27169 20995
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 27249 20995 27307 21001
rect 27249 20961 27261 20995
rect 27295 20961 27307 20995
rect 27249 20955 27307 20961
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20992 28595 20995
rect 29086 20992 29092 21004
rect 28583 20964 29092 20992
rect 28583 20961 28595 20964
rect 28537 20955 28595 20961
rect 23753 20927 23811 20933
rect 23753 20893 23765 20927
rect 23799 20924 23811 20927
rect 24302 20924 24308 20936
rect 23799 20896 24308 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24670 20884 24676 20936
rect 24728 20924 24734 20936
rect 24837 20927 24895 20933
rect 24837 20924 24849 20927
rect 24728 20896 24849 20924
rect 24728 20884 24734 20896
rect 24837 20893 24849 20896
rect 24883 20893 24895 20927
rect 27172 20924 27200 20955
rect 29086 20952 29092 20964
rect 29144 20952 29150 21004
rect 27614 20924 27620 20936
rect 27172 20896 27620 20924
rect 24837 20887 24895 20893
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 28350 20884 28356 20936
rect 28408 20884 28414 20936
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20924 28687 20927
rect 28810 20924 28816 20936
rect 28675 20896 28816 20924
rect 28675 20893 28687 20896
rect 28629 20887 28687 20893
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 23937 20859 23995 20865
rect 23937 20825 23949 20859
rect 23983 20856 23995 20859
rect 27154 20856 27160 20868
rect 23983 20828 27160 20856
rect 23983 20825 23995 20828
rect 23937 20819 23995 20825
rect 27154 20816 27160 20828
rect 27212 20816 27218 20868
rect 29196 20856 29224 21100
rect 32493 21097 32505 21100
rect 32539 21097 32551 21131
rect 32493 21091 32551 21097
rect 33134 21088 33140 21140
rect 33192 21128 33198 21140
rect 33597 21131 33655 21137
rect 33597 21128 33609 21131
rect 33192 21100 33609 21128
rect 33192 21088 33198 21100
rect 33597 21097 33609 21100
rect 33643 21128 33655 21131
rect 34330 21128 34336 21140
rect 33643 21100 34336 21128
rect 33643 21097 33655 21100
rect 33597 21091 33655 21097
rect 34330 21088 34336 21100
rect 34388 21088 34394 21140
rect 35253 21131 35311 21137
rect 35253 21097 35265 21131
rect 35299 21097 35311 21131
rect 35253 21091 35311 21097
rect 35621 21131 35679 21137
rect 35621 21097 35633 21131
rect 35667 21128 35679 21131
rect 35802 21128 35808 21140
rect 35667 21100 35808 21128
rect 35667 21097 35679 21100
rect 35621 21091 35679 21097
rect 31478 21020 31484 21072
rect 31536 21060 31542 21072
rect 35268 21060 35296 21091
rect 35802 21088 35808 21100
rect 35860 21088 35866 21140
rect 35894 21088 35900 21140
rect 35952 21128 35958 21140
rect 36173 21131 36231 21137
rect 36173 21128 36185 21131
rect 35952 21100 36185 21128
rect 35952 21088 35958 21100
rect 36173 21097 36185 21100
rect 36219 21128 36231 21131
rect 36219 21100 36492 21128
rect 36219 21097 36231 21100
rect 36173 21091 36231 21097
rect 36354 21060 36360 21072
rect 31536 21032 36360 21060
rect 31536 21020 31542 21032
rect 36354 21020 36360 21032
rect 36412 21020 36418 21072
rect 36464 21060 36492 21100
rect 36722 21088 36728 21140
rect 36780 21088 36786 21140
rect 37458 21088 37464 21140
rect 37516 21128 37522 21140
rect 37553 21131 37611 21137
rect 37553 21128 37565 21131
rect 37516 21100 37565 21128
rect 37516 21088 37522 21100
rect 37553 21097 37565 21100
rect 37599 21097 37611 21131
rect 39850 21128 39856 21140
rect 37553 21091 37611 21097
rect 37660 21100 39856 21128
rect 37660 21060 37688 21100
rect 39850 21088 39856 21100
rect 39908 21088 39914 21140
rect 40034 21088 40040 21140
rect 40092 21128 40098 21140
rect 40129 21131 40187 21137
rect 40129 21128 40141 21131
rect 40092 21100 40141 21128
rect 40092 21088 40098 21100
rect 40129 21097 40141 21100
rect 40175 21097 40187 21131
rect 40129 21091 40187 21097
rect 40218 21088 40224 21140
rect 40276 21128 40282 21140
rect 40681 21131 40739 21137
rect 40681 21128 40693 21131
rect 40276 21100 40693 21128
rect 40276 21088 40282 21100
rect 40681 21097 40693 21100
rect 40727 21097 40739 21131
rect 40681 21091 40739 21097
rect 37826 21060 37832 21072
rect 36464 21032 37688 21060
rect 37752 21032 37832 21060
rect 33134 20992 33140 21004
rect 32692 20964 33140 20992
rect 31481 20927 31539 20933
rect 31481 20893 31493 20927
rect 31527 20924 31539 20927
rect 31754 20924 31760 20936
rect 31527 20896 31760 20924
rect 31527 20893 31539 20896
rect 31481 20887 31539 20893
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 32214 20884 32220 20936
rect 32272 20924 32278 20936
rect 32692 20933 32720 20964
rect 33134 20952 33140 20964
rect 33192 20952 33198 21004
rect 35618 20992 35624 21004
rect 35268 20964 35624 20992
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32272 20896 32689 20924
rect 32272 20884 32278 20896
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 32769 20927 32827 20933
rect 32769 20893 32781 20927
rect 32815 20924 32827 20927
rect 32858 20924 32864 20936
rect 32815 20896 32864 20924
rect 32815 20893 32827 20896
rect 32769 20887 32827 20893
rect 32858 20884 32864 20896
rect 32916 20884 32922 20936
rect 32950 20884 32956 20936
rect 33008 20884 33014 20936
rect 33042 20884 33048 20936
rect 33100 20884 33106 20936
rect 35268 20933 35296 20964
rect 35618 20952 35624 20964
rect 35676 20952 35682 21004
rect 35986 20952 35992 21004
rect 36044 20992 36050 21004
rect 37752 21001 37780 21032
rect 37826 21020 37832 21032
rect 37884 21020 37890 21072
rect 38013 21063 38071 21069
rect 38013 21029 38025 21063
rect 38059 21029 38071 21063
rect 38013 21023 38071 21029
rect 36817 20995 36875 21001
rect 36817 20992 36829 20995
rect 36044 20964 36829 20992
rect 36044 20952 36050 20964
rect 36817 20961 36829 20964
rect 36863 20961 36875 20995
rect 36817 20955 36875 20961
rect 37737 20995 37795 21001
rect 37737 20961 37749 20995
rect 37783 20961 37795 20995
rect 38028 20992 38056 21023
rect 40494 21020 40500 21072
rect 40552 21060 40558 21072
rect 41141 21063 41199 21069
rect 41141 21060 41153 21063
rect 40552 21032 41153 21060
rect 40552 21020 40558 21032
rect 41141 21029 41153 21032
rect 41187 21029 41199 21063
rect 41141 21023 41199 21029
rect 38470 20992 38476 21004
rect 38028 20964 38476 20992
rect 37737 20955 37795 20961
rect 38470 20952 38476 20964
rect 38528 20992 38534 21004
rect 38933 20995 38991 21001
rect 38933 20992 38945 20995
rect 38528 20964 38945 20992
rect 38528 20952 38534 20964
rect 38933 20961 38945 20964
rect 38979 20961 38991 20995
rect 38933 20955 38991 20961
rect 39022 20952 39028 21004
rect 39080 20952 39086 21004
rect 35253 20927 35311 20933
rect 35253 20893 35265 20927
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 35437 20927 35495 20933
rect 35437 20893 35449 20927
rect 35483 20924 35495 20927
rect 35526 20924 35532 20936
rect 35483 20896 35532 20924
rect 35483 20893 35495 20896
rect 35437 20887 35495 20893
rect 35526 20884 35532 20896
rect 35584 20884 35590 20936
rect 36722 20884 36728 20936
rect 36780 20884 36786 20936
rect 37829 20927 37887 20933
rect 37829 20893 37841 20927
rect 37875 20924 37887 20927
rect 37918 20924 37924 20936
rect 37875 20896 37924 20924
rect 37875 20893 37887 20896
rect 37829 20887 37887 20893
rect 37918 20884 37924 20896
rect 37976 20884 37982 20936
rect 38746 20884 38752 20936
rect 38804 20924 38810 20936
rect 38841 20927 38899 20933
rect 38841 20924 38853 20927
rect 38804 20896 38853 20924
rect 38804 20884 38810 20896
rect 38841 20893 38853 20896
rect 38887 20893 38899 20927
rect 39206 20924 39212 20936
rect 38841 20887 38899 20893
rect 38948 20896 39212 20924
rect 27264 20828 29224 20856
rect 24762 20788 24768 20800
rect 23676 20760 24768 20788
rect 24762 20748 24768 20760
rect 24820 20788 24826 20800
rect 27264 20788 27292 20828
rect 30374 20816 30380 20868
rect 30432 20856 30438 20868
rect 31214 20859 31272 20865
rect 31214 20856 31226 20859
rect 30432 20828 31226 20856
rect 30432 20816 30438 20828
rect 31214 20825 31226 20828
rect 31260 20825 31272 20859
rect 35894 20856 35900 20868
rect 31214 20819 31272 20825
rect 32784 20828 35900 20856
rect 32784 20800 32812 20828
rect 35894 20816 35900 20828
rect 35952 20816 35958 20868
rect 37550 20816 37556 20868
rect 37608 20816 37614 20868
rect 37734 20816 37740 20868
rect 37792 20856 37798 20868
rect 38948 20856 38976 20896
rect 39206 20884 39212 20896
rect 39264 20884 39270 20936
rect 40126 20884 40132 20936
rect 40184 20924 40190 20936
rect 40313 20927 40371 20933
rect 40313 20924 40325 20927
rect 40184 20896 40325 20924
rect 40184 20884 40190 20896
rect 40313 20893 40325 20896
rect 40359 20893 40371 20927
rect 40313 20887 40371 20893
rect 40494 20884 40500 20936
rect 40552 20884 40558 20936
rect 40037 20859 40095 20865
rect 40037 20856 40049 20859
rect 37792 20828 38976 20856
rect 39224 20828 40049 20856
rect 37792 20816 37798 20828
rect 24820 20760 27292 20788
rect 27341 20791 27399 20797
rect 24820 20748 24826 20760
rect 27341 20757 27353 20791
rect 27387 20788 27399 20791
rect 29086 20788 29092 20800
rect 27387 20760 29092 20788
rect 27387 20757 27399 20760
rect 27341 20751 27399 20757
rect 29086 20748 29092 20760
rect 29144 20748 29150 20800
rect 30101 20791 30159 20797
rect 30101 20757 30113 20791
rect 30147 20788 30159 20791
rect 31018 20788 31024 20800
rect 30147 20760 31024 20788
rect 30147 20757 30159 20760
rect 30101 20751 30159 20757
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 32766 20748 32772 20800
rect 32824 20748 32830 20800
rect 35434 20748 35440 20800
rect 35492 20788 35498 20800
rect 35802 20788 35808 20800
rect 35492 20760 35808 20788
rect 35492 20748 35498 20760
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 37093 20791 37151 20797
rect 37093 20757 37105 20791
rect 37139 20788 37151 20791
rect 38010 20788 38016 20800
rect 37139 20760 38016 20788
rect 37139 20757 37151 20760
rect 37093 20751 37151 20757
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 39022 20748 39028 20800
rect 39080 20788 39086 20800
rect 39224 20797 39252 20828
rect 40037 20825 40049 20828
rect 40083 20825 40095 20859
rect 40037 20819 40095 20825
rect 40402 20816 40408 20868
rect 40460 20856 40466 20868
rect 40460 20828 41276 20856
rect 40460 20816 40466 20828
rect 39209 20791 39267 20797
rect 39209 20788 39221 20791
rect 39080 20760 39221 20788
rect 39080 20748 39086 20760
rect 39209 20757 39221 20760
rect 39255 20757 39267 20791
rect 41248 20788 41276 20828
rect 41322 20816 41328 20868
rect 41380 20856 41386 20868
rect 42889 20859 42947 20865
rect 42889 20856 42901 20859
rect 41380 20828 42901 20856
rect 41380 20816 41386 20828
rect 42889 20825 42901 20828
rect 42935 20825 42947 20859
rect 42889 20819 42947 20825
rect 43257 20859 43315 20865
rect 43257 20825 43269 20859
rect 43303 20856 43315 20859
rect 43346 20856 43352 20868
rect 43303 20828 43352 20856
rect 43303 20825 43315 20828
rect 43257 20819 43315 20825
rect 43346 20816 43352 20828
rect 43404 20856 43410 20868
rect 43990 20856 43996 20868
rect 43404 20828 43996 20856
rect 43404 20816 43410 20828
rect 43990 20816 43996 20828
rect 44048 20816 44054 20868
rect 41693 20791 41751 20797
rect 41693 20788 41705 20791
rect 41248 20760 41705 20788
rect 39209 20751 39267 20757
rect 41693 20757 41705 20760
rect 41739 20757 41751 20791
rect 41693 20751 41751 20757
rect 42242 20748 42248 20800
rect 42300 20748 42306 20800
rect 1104 20698 43884 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 43884 20698
rect 1104 20624 43884 20646
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17218 20584 17224 20596
rect 17175 20556 17224 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 12986 20408 12992 20460
rect 13044 20408 13050 20460
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20448 13691 20451
rect 14292 20448 14320 20547
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20273 20587 20331 20593
rect 20273 20584 20285 20587
rect 20036 20556 20285 20584
rect 20036 20544 20042 20556
rect 20273 20553 20285 20556
rect 20319 20553 20331 20587
rect 20273 20547 20331 20553
rect 20438 20544 20444 20596
rect 20496 20544 20502 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 22738 20584 22744 20596
rect 22695 20556 22744 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 25406 20544 25412 20596
rect 25464 20544 25470 20596
rect 27430 20584 27436 20596
rect 25608 20556 27436 20584
rect 14737 20519 14795 20525
rect 14737 20485 14749 20519
rect 14783 20516 14795 20519
rect 18230 20516 18236 20528
rect 14783 20488 18236 20516
rect 14783 20485 14795 20488
rect 14737 20479 14795 20485
rect 13679 20420 14320 20448
rect 13679 20417 13691 20420
rect 13633 20411 13691 20417
rect 14642 20408 14648 20460
rect 14700 20408 14706 20460
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14752 20380 14780 20479
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 20073 20519 20131 20525
rect 20073 20485 20085 20519
rect 20119 20516 20131 20519
rect 20714 20516 20720 20528
rect 20119 20488 20720 20516
rect 20119 20485 20131 20488
rect 20073 20479 20131 20485
rect 20714 20476 20720 20488
rect 20772 20516 20778 20528
rect 20898 20516 20904 20528
rect 20772 20488 20904 20516
rect 20772 20476 20778 20488
rect 20898 20476 20904 20488
rect 20956 20476 20962 20528
rect 23658 20516 23664 20528
rect 23492 20488 23664 20516
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 13504 20352 14780 20380
rect 14921 20383 14979 20389
rect 13504 20340 13510 20352
rect 14921 20349 14933 20383
rect 14967 20380 14979 20383
rect 15102 20380 15108 20392
rect 14967 20352 15108 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 15488 20380 15516 20411
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15620 20420 15669 20448
rect 15620 20408 15626 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 15988 20420 16865 20448
rect 15988 20408 15994 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17678 20408 17684 20460
rect 17736 20408 17742 20460
rect 17770 20408 17776 20460
rect 17828 20448 17834 20460
rect 18141 20451 18199 20457
rect 18141 20448 18153 20451
rect 17828 20420 18153 20448
rect 17828 20408 17834 20420
rect 18141 20417 18153 20420
rect 18187 20417 18199 20451
rect 18141 20411 18199 20417
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 19116 20420 19165 20448
rect 19116 20408 19122 20420
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 19484 20420 19533 20448
rect 19484 20408 19490 20420
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 21082 20408 21088 20460
rect 21140 20408 21146 20460
rect 23492 20457 23520 20488
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20417 23535 20451
rect 23750 20448 23756 20460
rect 23477 20411 23535 20417
rect 23584 20420 23756 20448
rect 15746 20380 15752 20392
rect 15488 20352 15752 20380
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 17865 20383 17923 20389
rect 17865 20349 17877 20383
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 15470 20272 15476 20324
rect 15528 20312 15534 20324
rect 15654 20312 15660 20324
rect 15528 20284 15660 20312
rect 15528 20272 15534 20284
rect 15654 20272 15660 20284
rect 15712 20312 15718 20324
rect 17880 20312 17908 20343
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 18012 20352 18061 20380
rect 18012 20340 18018 20352
rect 18049 20349 18061 20352
rect 18095 20349 18107 20383
rect 18049 20343 18107 20349
rect 21634 20340 21640 20392
rect 21692 20380 21698 20392
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 21692 20352 22753 20380
rect 21692 20340 21698 20352
rect 22741 20349 22753 20352
rect 22787 20349 22799 20383
rect 22741 20343 22799 20349
rect 22925 20383 22983 20389
rect 22925 20349 22937 20383
rect 22971 20380 22983 20383
rect 23584 20380 23612 20420
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 25608 20457 25636 20556
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 27522 20544 27528 20596
rect 27580 20584 27586 20596
rect 27709 20587 27767 20593
rect 27709 20584 27721 20587
rect 27580 20556 27721 20584
rect 27580 20544 27586 20556
rect 27709 20553 27721 20556
rect 27755 20553 27767 20587
rect 27709 20547 27767 20553
rect 28169 20587 28227 20593
rect 28169 20553 28181 20587
rect 28215 20584 28227 20587
rect 28350 20584 28356 20596
rect 28215 20556 28356 20584
rect 28215 20553 28227 20556
rect 28169 20547 28227 20553
rect 28350 20544 28356 20556
rect 28408 20544 28414 20596
rect 28644 20556 29224 20584
rect 25682 20476 25688 20528
rect 25740 20476 25746 20528
rect 27154 20476 27160 20528
rect 27212 20516 27218 20528
rect 28644 20525 28672 20556
rect 27249 20519 27307 20525
rect 27249 20516 27261 20519
rect 27212 20488 27261 20516
rect 27212 20476 27218 20488
rect 27249 20485 27261 20488
rect 27295 20485 27307 20519
rect 28629 20519 28687 20525
rect 28629 20516 28641 20519
rect 27249 20479 27307 20485
rect 27448 20488 28641 20516
rect 27448 20460 27476 20488
rect 28629 20485 28641 20488
rect 28675 20485 28687 20519
rect 28629 20479 28687 20485
rect 29086 20476 29092 20528
rect 29144 20476 29150 20528
rect 29196 20516 29224 20556
rect 30558 20544 30564 20596
rect 30616 20544 30622 20596
rect 31757 20587 31815 20593
rect 31757 20553 31769 20587
rect 31803 20584 31815 20587
rect 32214 20584 32220 20596
rect 31803 20556 32220 20584
rect 31803 20553 31815 20556
rect 31757 20547 31815 20553
rect 32214 20544 32220 20556
rect 32272 20544 32278 20596
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 34977 20587 35035 20593
rect 34977 20584 34989 20587
rect 34848 20556 34989 20584
rect 34848 20544 34854 20556
rect 34977 20553 34989 20556
rect 35023 20553 35035 20587
rect 34977 20547 35035 20553
rect 35989 20587 36047 20593
rect 35989 20553 36001 20587
rect 36035 20584 36047 20587
rect 37458 20584 37464 20596
rect 36035 20556 37464 20584
rect 36035 20553 36047 20556
rect 35989 20547 36047 20553
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 39301 20587 39359 20593
rect 39301 20553 39313 20587
rect 39347 20584 39359 20587
rect 40126 20584 40132 20596
rect 39347 20556 40132 20584
rect 39347 20553 39359 20556
rect 39301 20547 39359 20553
rect 40126 20544 40132 20556
rect 40184 20544 40190 20596
rect 40310 20544 40316 20596
rect 40368 20544 40374 20596
rect 41969 20587 42027 20593
rect 41969 20553 41981 20587
rect 42015 20584 42027 20587
rect 42702 20584 42708 20596
rect 42015 20556 42708 20584
rect 42015 20553 42027 20556
rect 41969 20547 42027 20553
rect 42702 20544 42708 20556
rect 42760 20544 42766 20596
rect 29196 20488 30880 20516
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 22971 20352 23612 20380
rect 23661 20383 23719 20389
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 23661 20349 23673 20383
rect 23707 20349 23719 20383
rect 25792 20380 25820 20411
rect 25958 20408 25964 20460
rect 26016 20408 26022 20460
rect 27430 20408 27436 20460
rect 27488 20408 27494 20460
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20448 27583 20451
rect 27614 20448 27620 20460
rect 27571 20420 27620 20448
rect 27571 20417 27583 20420
rect 27525 20411 27583 20417
rect 27614 20408 27620 20420
rect 27672 20448 27678 20460
rect 28353 20451 28411 20457
rect 28353 20448 28365 20451
rect 27672 20420 28365 20448
rect 27672 20408 27678 20420
rect 28353 20417 28365 20420
rect 28399 20448 28411 20451
rect 28399 20420 28847 20448
rect 28399 20417 28411 20420
rect 28353 20411 28411 20417
rect 27890 20380 27896 20392
rect 25792 20352 27896 20380
rect 23661 20343 23719 20349
rect 18138 20312 18144 20324
rect 15712 20284 17816 20312
rect 17880 20284 18144 20312
rect 15712 20272 15718 20284
rect 13170 20204 13176 20256
rect 13228 20204 13234 20256
rect 13814 20204 13820 20256
rect 13872 20204 13878 20256
rect 15286 20204 15292 20256
rect 15344 20244 15350 20256
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15344 20216 15853 20244
rect 15344 20204 15350 20216
rect 15841 20213 15853 20216
rect 15887 20213 15899 20247
rect 17788 20244 17816 20284
rect 18138 20272 18144 20284
rect 18196 20312 18202 20324
rect 18782 20312 18788 20324
rect 18196 20284 18788 20312
rect 18196 20272 18202 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19334 20312 19340 20324
rect 19168 20284 19340 20312
rect 18322 20244 18328 20256
rect 17788 20216 18328 20244
rect 15841 20207 15899 20213
rect 18322 20204 18328 20216
rect 18380 20244 18386 20256
rect 19168 20244 19196 20284
rect 19334 20272 19340 20284
rect 19392 20312 19398 20324
rect 23566 20312 23572 20324
rect 19392 20284 23572 20312
rect 19392 20272 19398 20284
rect 20272 20253 20300 20284
rect 23566 20272 23572 20284
rect 23624 20312 23630 20324
rect 23676 20312 23704 20343
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 27982 20340 27988 20392
rect 28040 20380 28046 20392
rect 28445 20383 28503 20389
rect 28445 20380 28457 20383
rect 28040 20352 28457 20380
rect 28040 20340 28046 20352
rect 28445 20349 28457 20352
rect 28491 20349 28503 20383
rect 28819 20380 28847 20420
rect 28902 20408 28908 20460
rect 28960 20448 28966 20460
rect 29181 20451 29239 20457
rect 29181 20448 29193 20451
rect 28960 20420 29193 20448
rect 28960 20408 28966 20420
rect 29181 20417 29193 20420
rect 29227 20417 29239 20451
rect 29181 20411 29239 20417
rect 30742 20380 30748 20392
rect 28819 20352 30748 20380
rect 28445 20343 28503 20349
rect 30742 20340 30748 20352
rect 30800 20340 30806 20392
rect 30852 20389 30880 20488
rect 31662 20476 31668 20528
rect 31720 20516 31726 20528
rect 40328 20516 40356 20544
rect 41874 20516 41880 20528
rect 31720 20488 32720 20516
rect 31720 20476 31726 20488
rect 31110 20408 31116 20460
rect 31168 20408 31174 20460
rect 32306 20408 32312 20460
rect 32364 20408 32370 20460
rect 32398 20408 32404 20460
rect 32456 20448 32462 20460
rect 32493 20451 32551 20457
rect 32493 20448 32505 20451
rect 32456 20420 32505 20448
rect 32456 20408 32462 20420
rect 32493 20417 32505 20420
rect 32539 20417 32551 20451
rect 32493 20411 32551 20417
rect 32582 20408 32588 20460
rect 32640 20408 32646 20460
rect 32692 20457 32720 20488
rect 33612 20488 40356 20516
rect 41722 20488 41880 20516
rect 32677 20451 32735 20457
rect 32677 20417 32689 20451
rect 32723 20448 32735 20451
rect 32766 20448 32772 20460
rect 32723 20420 32772 20448
rect 32723 20417 32735 20420
rect 32677 20411 32735 20417
rect 32766 20408 32772 20420
rect 32824 20408 32830 20460
rect 33042 20408 33048 20460
rect 33100 20448 33106 20460
rect 33612 20457 33640 20488
rect 33870 20457 33876 20460
rect 33597 20451 33655 20457
rect 33597 20448 33609 20451
rect 33100 20420 33609 20448
rect 33100 20408 33106 20420
rect 33597 20417 33609 20420
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 33864 20411 33876 20457
rect 33870 20408 33876 20411
rect 33928 20408 33934 20460
rect 35342 20408 35348 20460
rect 35400 20448 35406 20460
rect 35437 20451 35495 20457
rect 35437 20448 35449 20451
rect 35400 20420 35449 20448
rect 35400 20408 35406 20420
rect 35437 20417 35449 20420
rect 35483 20417 35495 20451
rect 35437 20411 35495 20417
rect 36906 20408 36912 20460
rect 36964 20408 36970 20460
rect 37642 20408 37648 20460
rect 37700 20408 37706 20460
rect 37829 20451 37887 20457
rect 37829 20417 37841 20451
rect 37875 20448 37887 20451
rect 38010 20448 38016 20460
rect 37875 20420 38016 20448
rect 37875 20417 37887 20420
rect 37829 20411 37887 20417
rect 38010 20408 38016 20420
rect 38068 20408 38074 20460
rect 38841 20451 38899 20457
rect 38841 20417 38853 20451
rect 38887 20448 38899 20451
rect 39117 20451 39175 20457
rect 38887 20420 39068 20448
rect 38887 20417 38899 20420
rect 38841 20411 38899 20417
rect 30837 20383 30895 20389
rect 30837 20349 30849 20383
rect 30883 20380 30895 20383
rect 33502 20380 33508 20392
rect 30883 20352 33508 20380
rect 30883 20349 30895 20352
rect 30837 20343 30895 20349
rect 33502 20340 33508 20352
rect 33560 20340 33566 20392
rect 34606 20340 34612 20392
rect 34664 20380 34670 20392
rect 35713 20383 35771 20389
rect 35713 20380 35725 20383
rect 34664 20352 35725 20380
rect 34664 20340 34670 20352
rect 35713 20349 35725 20352
rect 35759 20349 35771 20383
rect 35713 20343 35771 20349
rect 36170 20340 36176 20392
rect 36228 20380 36234 20392
rect 36633 20383 36691 20389
rect 36633 20380 36645 20383
rect 36228 20352 36645 20380
rect 36228 20340 36234 20352
rect 36633 20349 36645 20352
rect 36679 20349 36691 20383
rect 36633 20343 36691 20349
rect 38930 20340 38936 20392
rect 38988 20340 38994 20392
rect 39040 20380 39068 20420
rect 39117 20417 39129 20451
rect 39163 20448 39175 20451
rect 39206 20448 39212 20460
rect 39163 20420 39212 20448
rect 39163 20417 39175 20420
rect 39117 20411 39175 20417
rect 39206 20408 39212 20420
rect 39264 20408 39270 20460
rect 40236 20457 40264 20488
rect 41874 20476 41880 20488
rect 41932 20476 41938 20528
rect 40221 20451 40279 20457
rect 40221 20417 40233 20451
rect 40267 20417 40279 20451
rect 40221 20411 40279 20417
rect 42242 20408 42248 20460
rect 42300 20448 42306 20460
rect 42981 20451 43039 20457
rect 42981 20448 42993 20451
rect 42300 20420 42993 20448
rect 42300 20408 42306 20420
rect 42981 20417 42993 20420
rect 43027 20417 43039 20451
rect 42981 20411 43039 20417
rect 39040 20352 39160 20380
rect 39132 20324 39160 20352
rect 40494 20340 40500 20392
rect 40552 20340 40558 20392
rect 23624 20284 23704 20312
rect 23624 20272 23630 20284
rect 28810 20272 28816 20324
rect 28868 20312 28874 20324
rect 32398 20312 32404 20324
rect 28868 20284 32404 20312
rect 28868 20272 28874 20284
rect 32398 20272 32404 20284
rect 32456 20272 32462 20324
rect 36725 20315 36783 20321
rect 32692 20284 33640 20312
rect 18380 20216 19196 20244
rect 20257 20247 20315 20253
rect 18380 20204 18386 20216
rect 20257 20213 20269 20247
rect 20303 20213 20315 20247
rect 20257 20207 20315 20213
rect 20898 20204 20904 20256
rect 20956 20204 20962 20256
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 22462 20244 22468 20256
rect 22327 20216 22468 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 27338 20204 27344 20256
rect 27396 20204 27402 20256
rect 28350 20204 28356 20256
rect 28408 20244 28414 20256
rect 28902 20244 28908 20256
rect 28408 20216 28908 20244
rect 28408 20204 28414 20216
rect 28902 20204 28908 20216
rect 28960 20204 28966 20256
rect 30098 20204 30104 20256
rect 30156 20204 30162 20256
rect 31018 20204 31024 20256
rect 31076 20204 31082 20256
rect 31386 20204 31392 20256
rect 31444 20244 31450 20256
rect 32692 20244 32720 20284
rect 31444 20216 32720 20244
rect 31444 20204 31450 20216
rect 32766 20204 32772 20256
rect 32824 20244 32830 20256
rect 32861 20247 32919 20253
rect 32861 20244 32873 20247
rect 32824 20216 32873 20244
rect 32824 20204 32830 20216
rect 32861 20213 32873 20216
rect 32907 20213 32919 20247
rect 33612 20244 33640 20284
rect 36725 20281 36737 20315
rect 36771 20312 36783 20315
rect 37366 20312 37372 20324
rect 36771 20284 37372 20312
rect 36771 20281 36783 20284
rect 36725 20275 36783 20281
rect 37366 20272 37372 20284
rect 37424 20312 37430 20324
rect 37424 20284 38884 20312
rect 37424 20272 37430 20284
rect 34606 20244 34612 20256
rect 33612 20216 34612 20244
rect 32861 20207 32919 20213
rect 34606 20204 34612 20216
rect 34664 20204 34670 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 35529 20247 35587 20253
rect 35529 20244 35541 20247
rect 34756 20216 35541 20244
rect 34756 20204 34762 20216
rect 35529 20213 35541 20216
rect 35575 20244 35587 20247
rect 35618 20244 35624 20256
rect 35575 20216 35624 20244
rect 35575 20213 35587 20216
rect 35529 20207 35587 20213
rect 35618 20204 35624 20216
rect 35676 20204 35682 20256
rect 36817 20247 36875 20253
rect 36817 20213 36829 20247
rect 36863 20244 36875 20247
rect 37458 20244 37464 20256
rect 36863 20216 37464 20244
rect 36863 20213 36875 20216
rect 36817 20207 36875 20213
rect 37458 20204 37464 20216
rect 37516 20204 37522 20256
rect 37642 20204 37648 20256
rect 37700 20204 37706 20256
rect 38010 20204 38016 20256
rect 38068 20204 38074 20256
rect 38856 20253 38884 20284
rect 39114 20272 39120 20324
rect 39172 20272 39178 20324
rect 38841 20247 38899 20253
rect 38841 20213 38853 20247
rect 38887 20213 38899 20247
rect 38841 20207 38899 20213
rect 42886 20204 42892 20256
rect 42944 20204 42950 20256
rect 1104 20154 43884 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 43884 20154
rect 1104 20080 43884 20102
rect 12986 20000 12992 20052
rect 13044 20000 13050 20052
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 15654 20040 15660 20052
rect 14700 20012 15660 20040
rect 14700 20000 14706 20012
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16209 20043 16267 20049
rect 16209 20009 16221 20043
rect 16255 20040 16267 20043
rect 16298 20040 16304 20052
rect 16255 20012 16304 20040
rect 16255 20009 16267 20012
rect 16209 20003 16267 20009
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 18782 20000 18788 20052
rect 18840 20000 18846 20052
rect 19426 20000 19432 20052
rect 19484 20000 19490 20052
rect 21634 20000 21640 20052
rect 21692 20000 21698 20052
rect 22097 20043 22155 20049
rect 22097 20009 22109 20043
rect 22143 20040 22155 20043
rect 22186 20040 22192 20052
rect 22143 20012 22192 20040
rect 22143 20009 22155 20012
rect 22097 20003 22155 20009
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 23934 20040 23940 20052
rect 23716 20012 23940 20040
rect 23716 20000 23722 20012
rect 23934 20000 23940 20012
rect 23992 20040 23998 20052
rect 23992 20012 28212 20040
rect 23992 20000 23998 20012
rect 12529 19975 12587 19981
rect 12529 19941 12541 19975
rect 12575 19972 12587 19975
rect 23676 19972 23704 20000
rect 12575 19944 13676 19972
rect 12575 19941 12587 19944
rect 12529 19935 12587 19941
rect 13648 19916 13676 19944
rect 22756 19944 23704 19972
rect 13446 19864 13452 19916
rect 13504 19864 13510 19916
rect 13630 19864 13636 19916
rect 13688 19864 13694 19916
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19904 16911 19907
rect 16942 19904 16948 19916
rect 16899 19876 16948 19904
rect 16899 19873 16911 19876
rect 16853 19867 16911 19873
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 19978 19904 19984 19916
rect 19628 19876 19984 19904
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 13412 19808 14289 19836
rect 13412 19796 13418 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 14323 19808 15792 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 13372 19740 13768 19768
rect 13372 19709 13400 19740
rect 13357 19703 13415 19709
rect 13357 19669 13369 19703
rect 13403 19669 13415 19703
rect 13740 19700 13768 19740
rect 13814 19728 13820 19780
rect 13872 19768 13878 19780
rect 14522 19771 14580 19777
rect 14522 19768 14534 19771
rect 13872 19740 14534 19768
rect 13872 19728 13878 19740
rect 14522 19737 14534 19740
rect 14568 19737 14580 19771
rect 15764 19768 15792 19808
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 15896 19808 17417 19836
rect 15896 19796 15902 19808
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 19628 19845 19656 19876
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 22756 19913 22784 19944
rect 24302 19932 24308 19984
rect 24360 19972 24366 19984
rect 26142 19972 26148 19984
rect 24360 19944 26148 19972
rect 24360 19932 24366 19944
rect 26142 19932 26148 19944
rect 26200 19932 26206 19984
rect 28184 19972 28212 20012
rect 28258 20000 28264 20052
rect 28316 20000 28322 20052
rect 28718 20000 28724 20052
rect 28776 20000 28782 20052
rect 29825 20043 29883 20049
rect 29825 20009 29837 20043
rect 29871 20040 29883 20043
rect 30098 20040 30104 20052
rect 29871 20012 30104 20040
rect 29871 20009 29883 20012
rect 29825 20003 29883 20009
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 30374 20000 30380 20052
rect 30432 20000 30438 20052
rect 32122 20000 32128 20052
rect 32180 20040 32186 20052
rect 33137 20043 33195 20049
rect 33137 20040 33149 20043
rect 32180 20012 33149 20040
rect 32180 20000 32186 20012
rect 33137 20009 33149 20012
rect 33183 20009 33195 20043
rect 33137 20003 33195 20009
rect 33870 20000 33876 20052
rect 33928 20000 33934 20052
rect 34882 20000 34888 20052
rect 34940 20040 34946 20052
rect 36449 20043 36507 20049
rect 34940 20012 35572 20040
rect 34940 20000 34946 20012
rect 31570 19972 31576 19984
rect 28184 19944 31576 19972
rect 31570 19932 31576 19944
rect 31628 19932 31634 19984
rect 34606 19932 34612 19984
rect 34664 19972 34670 19984
rect 35544 19972 35572 20012
rect 36449 20009 36461 20043
rect 36495 20040 36507 20043
rect 36722 20040 36728 20052
rect 36495 20012 36728 20040
rect 36495 20009 36507 20012
rect 36449 20003 36507 20009
rect 36722 20000 36728 20012
rect 36780 20000 36786 20052
rect 38105 20043 38163 20049
rect 38105 20009 38117 20043
rect 38151 20040 38163 20043
rect 38562 20040 38568 20052
rect 38151 20012 38568 20040
rect 38151 20009 38163 20012
rect 38105 20003 38163 20009
rect 38562 20000 38568 20012
rect 38620 20000 38626 20052
rect 40221 20043 40279 20049
rect 40221 20009 40233 20043
rect 40267 20040 40279 20043
rect 40494 20040 40500 20052
rect 40267 20012 40500 20040
rect 40267 20009 40279 20012
rect 40221 20003 40279 20009
rect 40494 20000 40500 20012
rect 40552 20000 40558 20052
rect 43254 20000 43260 20052
rect 43312 20000 43318 20052
rect 37642 19972 37648 19984
rect 34664 19944 35480 19972
rect 35544 19944 37648 19972
rect 34664 19932 34670 19944
rect 22741 19907 22799 19913
rect 22741 19873 22753 19907
rect 22787 19873 22799 19907
rect 22741 19867 22799 19873
rect 23566 19864 23572 19916
rect 23624 19864 23630 19916
rect 24854 19904 24860 19916
rect 24596 19876 24860 19904
rect 17661 19839 17719 19845
rect 17661 19836 17673 19839
rect 17552 19808 17673 19836
rect 17552 19796 17558 19808
rect 17661 19805 17673 19808
rect 17707 19805 17719 19839
rect 17661 19799 17719 19805
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 22002 19836 22008 19848
rect 20303 19808 22008 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 16850 19768 16856 19780
rect 15764 19740 16856 19768
rect 14522 19731 14580 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 19720 19768 19748 19799
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 22462 19796 22468 19848
rect 22520 19796 22526 19848
rect 23290 19796 23296 19848
rect 23348 19796 23354 19848
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19836 23443 19839
rect 23750 19836 23756 19848
rect 23431 19808 23756 19836
rect 23431 19805 23443 19808
rect 23385 19799 23443 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 24486 19796 24492 19848
rect 24544 19836 24550 19848
rect 24596 19845 24624 19876
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 28000 19904 28212 19912
rect 28810 19904 28816 19916
rect 27724 19884 28816 19904
rect 27724 19876 28028 19884
rect 28184 19876 28816 19884
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24544 19808 24593 19836
rect 24544 19796 24550 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 27249 19839 27307 19845
rect 27249 19805 27261 19839
rect 27295 19836 27307 19839
rect 27430 19836 27436 19848
rect 27295 19808 27436 19836
rect 27295 19805 27307 19808
rect 27249 19799 27307 19805
rect 27430 19796 27436 19808
rect 27488 19796 27494 19848
rect 27724 19845 27752 19876
rect 28810 19864 28816 19876
rect 28868 19864 28874 19916
rect 28902 19864 28908 19916
rect 28960 19904 28966 19916
rect 31110 19904 31116 19916
rect 28960 19876 31116 19904
rect 28960 19864 28966 19876
rect 31110 19864 31116 19876
rect 31168 19864 31174 19916
rect 34790 19864 34796 19916
rect 34848 19904 34854 19916
rect 35452 19913 35480 19944
rect 37642 19932 37648 19944
rect 37700 19932 37706 19984
rect 37737 19975 37795 19981
rect 37737 19941 37749 19975
rect 37783 19972 37795 19975
rect 37826 19972 37832 19984
rect 37783 19944 37832 19972
rect 37783 19941 37795 19944
rect 37737 19935 37795 19941
rect 37826 19932 37832 19944
rect 37884 19932 37890 19984
rect 40402 19932 40408 19984
rect 40460 19972 40466 19984
rect 40681 19975 40739 19981
rect 40681 19972 40693 19975
rect 40460 19944 40693 19972
rect 40460 19932 40466 19944
rect 40681 19941 40693 19944
rect 40727 19941 40739 19975
rect 40681 19935 40739 19941
rect 35437 19907 35495 19913
rect 34848 19876 35296 19904
rect 34848 19864 34854 19876
rect 27709 19839 27767 19845
rect 27709 19805 27721 19839
rect 27755 19805 27767 19839
rect 27709 19799 27767 19805
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 17920 19740 19748 19768
rect 20524 19771 20582 19777
rect 17920 19728 17926 19740
rect 20524 19737 20536 19771
rect 20570 19768 20582 19771
rect 20898 19768 20904 19780
rect 20570 19740 20904 19768
rect 20570 19737 20582 19740
rect 20524 19731 20582 19737
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 23768 19768 23796 19796
rect 24673 19771 24731 19777
rect 24673 19768 24685 19771
rect 23768 19740 24685 19768
rect 24673 19737 24685 19740
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 27893 19771 27951 19777
rect 27893 19737 27905 19771
rect 27939 19737 27951 19771
rect 27893 19731 27951 19737
rect 15562 19700 15568 19712
rect 13740 19672 15568 19700
rect 13357 19663 13415 19669
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16574 19660 16580 19712
rect 16632 19660 16638 19712
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 18230 19700 18236 19712
rect 16715 19672 18236 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 22554 19660 22560 19712
rect 22612 19660 22618 19712
rect 23569 19703 23627 19709
rect 23569 19669 23581 19703
rect 23615 19700 23627 19703
rect 23658 19700 23664 19712
rect 23615 19672 23664 19700
rect 23615 19669 23627 19672
rect 23569 19663 23627 19669
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 27065 19703 27123 19709
rect 27065 19669 27077 19703
rect 27111 19700 27123 19703
rect 27246 19700 27252 19712
rect 27111 19672 27252 19700
rect 27111 19669 27123 19672
rect 27065 19663 27123 19669
rect 27246 19660 27252 19672
rect 27304 19660 27310 19712
rect 27908 19700 27936 19731
rect 27982 19728 27988 19780
rect 28040 19728 28046 19780
rect 28092 19768 28120 19799
rect 29178 19796 29184 19848
rect 29236 19836 29242 19848
rect 30561 19839 30619 19845
rect 30561 19836 30573 19839
rect 29236 19808 30573 19836
rect 29236 19796 29242 19808
rect 30561 19805 30573 19808
rect 30607 19805 30619 19839
rect 30561 19799 30619 19805
rect 30653 19839 30711 19845
rect 30653 19805 30665 19839
rect 30699 19836 30711 19839
rect 30834 19836 30840 19848
rect 30699 19808 30840 19836
rect 30699 19805 30711 19808
rect 30653 19799 30711 19805
rect 30834 19796 30840 19808
rect 30892 19796 30898 19848
rect 30929 19839 30987 19845
rect 30929 19805 30941 19839
rect 30975 19836 30987 19839
rect 31018 19836 31024 19848
rect 30975 19808 31024 19836
rect 30975 19805 30987 19808
rect 30929 19799 30987 19805
rect 31018 19796 31024 19808
rect 31076 19796 31082 19848
rect 31754 19796 31760 19848
rect 31812 19836 31818 19848
rect 33042 19836 33048 19848
rect 31812 19808 33048 19836
rect 31812 19796 31818 19808
rect 33042 19796 33048 19808
rect 33100 19796 33106 19848
rect 35268 19845 35296 19876
rect 35437 19873 35449 19907
rect 35483 19873 35495 19907
rect 35437 19867 35495 19873
rect 38010 19864 38016 19916
rect 38068 19904 38074 19916
rect 38068 19876 40080 19904
rect 38068 19864 38074 19876
rect 34057 19839 34115 19845
rect 34057 19805 34069 19839
rect 34103 19836 34115 19839
rect 35253 19839 35311 19845
rect 34103 19808 34928 19836
rect 34103 19805 34115 19808
rect 34057 19799 34115 19805
rect 28166 19768 28172 19780
rect 28092 19740 28172 19768
rect 28166 19728 28172 19740
rect 28224 19728 28230 19780
rect 29362 19768 29368 19780
rect 28276 19740 29368 19768
rect 28276 19700 28304 19740
rect 29362 19728 29368 19740
rect 29420 19728 29426 19780
rect 30745 19771 30803 19777
rect 30745 19737 30757 19771
rect 30791 19768 30803 19771
rect 30791 19740 31754 19768
rect 30791 19737 30803 19740
rect 30745 19731 30803 19737
rect 27908 19672 28304 19700
rect 31726 19700 31754 19740
rect 31846 19728 31852 19780
rect 31904 19768 31910 19780
rect 32002 19771 32060 19777
rect 32002 19768 32014 19771
rect 31904 19740 32014 19768
rect 31904 19728 31910 19740
rect 32002 19737 32014 19740
rect 32048 19737 32060 19771
rect 34698 19768 34704 19780
rect 32002 19731 32060 19737
rect 33060 19740 34704 19768
rect 33060 19700 33088 19740
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 34900 19709 34928 19808
rect 35253 19805 35265 19839
rect 35299 19805 35311 19839
rect 35253 19799 35311 19805
rect 36446 19796 36452 19848
rect 36504 19796 36510 19848
rect 36538 19796 36544 19848
rect 36596 19836 36602 19848
rect 36633 19839 36691 19845
rect 36633 19836 36645 19839
rect 36596 19808 36645 19836
rect 36596 19796 36602 19808
rect 36633 19805 36645 19808
rect 36679 19836 36691 19839
rect 37182 19836 37188 19848
rect 36679 19808 37188 19836
rect 36679 19805 36691 19808
rect 36633 19799 36691 19805
rect 37182 19796 37188 19808
rect 37240 19796 37246 19848
rect 37274 19796 37280 19848
rect 37332 19836 37338 19848
rect 37645 19839 37703 19845
rect 37645 19836 37657 19839
rect 37332 19808 37657 19836
rect 37332 19796 37338 19808
rect 37645 19805 37657 19808
rect 37691 19805 37703 19839
rect 37645 19799 37703 19805
rect 37734 19796 37740 19848
rect 37792 19836 37798 19848
rect 37829 19839 37887 19845
rect 37829 19836 37841 19839
rect 37792 19808 37841 19836
rect 37792 19796 37798 19808
rect 37829 19805 37841 19808
rect 37875 19805 37887 19839
rect 37829 19799 37887 19805
rect 37921 19839 37979 19845
rect 37921 19805 37933 19839
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 36906 19728 36912 19780
rect 36964 19768 36970 19780
rect 37366 19768 37372 19780
rect 36964 19740 37372 19768
rect 36964 19728 36970 19740
rect 37366 19728 37372 19740
rect 37424 19768 37430 19780
rect 37936 19768 37964 19799
rect 38654 19796 38660 19848
rect 38712 19836 38718 19848
rect 38841 19839 38899 19845
rect 38841 19836 38853 19839
rect 38712 19808 38853 19836
rect 38712 19796 38718 19808
rect 38841 19805 38853 19808
rect 38887 19805 38899 19839
rect 38841 19799 38899 19805
rect 38933 19839 38991 19845
rect 38933 19805 38945 19839
rect 38979 19805 38991 19839
rect 38933 19799 38991 19805
rect 37424 19740 37964 19768
rect 37424 19728 37430 19740
rect 38562 19728 38568 19780
rect 38620 19768 38626 19780
rect 38948 19768 38976 19799
rect 39022 19796 39028 19848
rect 39080 19796 39086 19848
rect 40052 19845 40080 19876
rect 40310 19864 40316 19916
rect 40368 19904 40374 19916
rect 41509 19907 41567 19913
rect 41509 19904 41521 19907
rect 40368 19876 41521 19904
rect 40368 19864 40374 19876
rect 41509 19873 41521 19876
rect 41555 19873 41567 19907
rect 41509 19867 41567 19873
rect 40037 19839 40095 19845
rect 40037 19805 40049 19839
rect 40083 19805 40095 19839
rect 40037 19799 40095 19805
rect 42886 19796 42892 19848
rect 42944 19796 42950 19848
rect 38620 19740 38976 19768
rect 39209 19771 39267 19777
rect 38620 19728 38626 19740
rect 39209 19737 39221 19771
rect 39255 19768 39267 19771
rect 41785 19771 41843 19777
rect 41785 19768 41797 19771
rect 39255 19740 41797 19768
rect 39255 19737 39267 19740
rect 39209 19731 39267 19737
rect 41785 19737 41797 19740
rect 41831 19737 41843 19771
rect 41785 19731 41843 19737
rect 31726 19672 33088 19700
rect 34885 19703 34943 19709
rect 34885 19669 34897 19703
rect 34931 19669 34943 19703
rect 34885 19663 34943 19669
rect 35345 19703 35403 19709
rect 35345 19669 35357 19703
rect 35391 19700 35403 19703
rect 35434 19700 35440 19712
rect 35391 19672 35440 19700
rect 35391 19669 35403 19672
rect 35345 19663 35403 19669
rect 35434 19660 35440 19672
rect 35492 19660 35498 19712
rect 39298 19660 39304 19712
rect 39356 19700 39362 19712
rect 39942 19700 39948 19712
rect 39356 19672 39948 19700
rect 39356 19660 39362 19672
rect 39942 19660 39948 19672
rect 40000 19660 40006 19712
rect 1104 19610 43884 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 43884 19610
rect 1104 19536 43884 19558
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 15562 19496 15568 19508
rect 14783 19468 15568 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 15930 19456 15936 19508
rect 15988 19456 15994 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18012 19468 18337 19496
rect 18012 19456 18018 19468
rect 18325 19465 18337 19468
rect 18371 19496 18383 19499
rect 18598 19496 18604 19508
rect 18371 19468 18604 19496
rect 18371 19465 18383 19468
rect 18325 19459 18383 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 19978 19496 19984 19508
rect 19843 19468 19984 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 22281 19499 22339 19505
rect 22281 19496 22293 19499
rect 20128 19468 22293 19496
rect 20128 19456 20134 19468
rect 22281 19465 22293 19468
rect 22327 19465 22339 19499
rect 22281 19459 22339 19465
rect 22738 19456 22744 19508
rect 22796 19456 22802 19508
rect 23658 19456 23664 19508
rect 23716 19456 23722 19508
rect 24118 19456 24124 19508
rect 24176 19456 24182 19508
rect 26237 19499 26295 19505
rect 26237 19465 26249 19499
rect 26283 19496 26295 19499
rect 26510 19496 26516 19508
rect 26283 19468 26516 19496
rect 26283 19465 26295 19468
rect 26237 19459 26295 19465
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 27157 19499 27215 19505
rect 27157 19465 27169 19499
rect 27203 19496 27215 19499
rect 27982 19496 27988 19508
rect 27203 19468 27988 19496
rect 27203 19465 27215 19468
rect 27157 19459 27215 19465
rect 27982 19456 27988 19468
rect 28040 19456 28046 19508
rect 28350 19456 28356 19508
rect 28408 19456 28414 19508
rect 28902 19456 28908 19508
rect 28960 19496 28966 19508
rect 31662 19496 31668 19508
rect 28960 19468 30144 19496
rect 28960 19456 28966 19468
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13602 19431 13660 19437
rect 13602 19428 13614 19431
rect 13228 19400 13614 19428
rect 13228 19388 13234 19400
rect 13602 19397 13614 19400
rect 13648 19397 13660 19431
rect 13602 19391 13660 19397
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 15436 19400 15608 19428
rect 15436 19388 15442 19400
rect 13354 19320 13360 19372
rect 13412 19320 13418 19372
rect 15286 19320 15292 19372
rect 15344 19320 15350 19372
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 15580 19369 15608 19400
rect 15746 19388 15752 19440
rect 15804 19428 15810 19440
rect 20714 19428 20720 19440
rect 15804 19400 20720 19428
rect 15804 19388 15810 19400
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19329 15623 19363
rect 15565 19323 15623 19329
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17880 19369 17908 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 21174 19388 21180 19440
rect 21232 19428 21238 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 21232 19400 22385 19428
rect 21232 19388 21238 19400
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 28258 19428 28264 19440
rect 28316 19437 28322 19440
rect 28228 19400 28264 19428
rect 22373 19391 22431 19397
rect 28258 19388 28264 19400
rect 28316 19391 28328 19437
rect 28368 19428 28396 19456
rect 30116 19440 30144 19468
rect 31404 19468 31668 19496
rect 29273 19431 29331 19437
rect 29273 19428 29285 19431
rect 28368 19400 29285 19428
rect 29273 19397 29285 19400
rect 29319 19397 29331 19431
rect 29273 19391 29331 19397
rect 28316 19388 28322 19391
rect 29362 19388 29368 19440
rect 29420 19388 29426 19440
rect 30098 19388 30104 19440
rect 30156 19428 30162 19440
rect 31404 19437 31432 19468
rect 31662 19456 31668 19468
rect 31720 19456 31726 19508
rect 31757 19499 31815 19505
rect 31757 19465 31769 19499
rect 31803 19496 31815 19499
rect 31846 19496 31852 19508
rect 31803 19468 31852 19496
rect 31803 19465 31815 19468
rect 31757 19459 31815 19465
rect 31846 19456 31852 19468
rect 31904 19456 31910 19508
rect 33962 19456 33968 19508
rect 34020 19496 34026 19508
rect 35161 19499 35219 19505
rect 35161 19496 35173 19499
rect 34020 19468 35173 19496
rect 34020 19456 34026 19468
rect 35161 19465 35173 19468
rect 35207 19496 35219 19499
rect 35802 19496 35808 19508
rect 35207 19468 35808 19496
rect 35207 19465 35219 19468
rect 35161 19459 35219 19465
rect 35802 19456 35808 19468
rect 35860 19456 35866 19508
rect 35989 19499 36047 19505
rect 35989 19465 36001 19499
rect 36035 19496 36047 19499
rect 36906 19496 36912 19508
rect 36035 19468 36912 19496
rect 36035 19465 36047 19468
rect 35989 19459 36047 19465
rect 30745 19431 30803 19437
rect 30745 19428 30757 19431
rect 30156 19400 30757 19428
rect 30156 19388 30162 19400
rect 30745 19397 30757 19400
rect 30791 19428 30803 19431
rect 31389 19431 31447 19437
rect 30791 19400 31340 19428
rect 30791 19397 30803 19400
rect 30745 19391 30803 19397
rect 17865 19363 17923 19369
rect 17000 19332 17816 19360
rect 17000 19320 17006 19332
rect 17788 19292 17816 19332
rect 17865 19329 17877 19363
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 18322 19320 18328 19372
rect 18380 19320 18386 19372
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19978 19360 19984 19372
rect 19751 19332 19984 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22002 19360 22008 19372
rect 21499 19332 22008 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 23753 19363 23811 19369
rect 23753 19360 23765 19363
rect 22336 19332 23765 19360
rect 22336 19320 22342 19332
rect 23753 19329 23765 19332
rect 23799 19329 23811 19363
rect 23753 19323 23811 19329
rect 24857 19363 24915 19369
rect 24857 19329 24869 19363
rect 24903 19329 24915 19363
rect 24857 19323 24915 19329
rect 25124 19363 25182 19369
rect 25124 19329 25136 19363
rect 25170 19360 25182 19363
rect 27798 19360 27804 19372
rect 25170 19332 27804 19360
rect 25170 19329 25182 19332
rect 25124 19323 25182 19329
rect 18966 19292 18972 19304
rect 17788 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19292 19030 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19024 19264 19901 19292
rect 19024 19252 19030 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 19904 19224 19932 19255
rect 20714 19252 20720 19304
rect 20772 19252 20778 19304
rect 22189 19295 22247 19301
rect 22189 19261 22201 19295
rect 22235 19292 22247 19295
rect 23569 19295 23627 19301
rect 23569 19292 23581 19295
rect 22235 19264 23581 19292
rect 22235 19261 22247 19264
rect 22189 19255 22247 19261
rect 23569 19261 23581 19264
rect 23615 19292 23627 19295
rect 23934 19292 23940 19304
rect 23615 19264 23940 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24578 19252 24584 19304
rect 24636 19292 24642 19304
rect 24872 19292 24900 19323
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 29178 19320 29184 19372
rect 29236 19320 29242 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 30374 19360 30380 19372
rect 29595 19332 30380 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 30374 19320 30380 19332
rect 30432 19360 30438 19372
rect 31205 19363 31263 19369
rect 31205 19360 31217 19363
rect 30432 19332 31217 19360
rect 30432 19320 30438 19332
rect 31205 19329 31217 19332
rect 31251 19329 31263 19363
rect 31312 19360 31340 19400
rect 31389 19397 31401 19431
rect 31435 19397 31447 19431
rect 31389 19391 31447 19397
rect 31481 19431 31539 19437
rect 31481 19397 31493 19431
rect 31527 19428 31539 19431
rect 31527 19400 31754 19428
rect 31527 19397 31539 19400
rect 31481 19391 31539 19397
rect 31570 19360 31576 19372
rect 31312 19332 31576 19360
rect 31205 19323 31263 19329
rect 31570 19320 31576 19332
rect 31628 19320 31634 19372
rect 31726 19360 31754 19400
rect 33502 19388 33508 19440
rect 33560 19428 33566 19440
rect 36004 19428 36032 19459
rect 36906 19456 36912 19468
rect 36964 19456 36970 19508
rect 37829 19499 37887 19505
rect 37829 19465 37841 19499
rect 37875 19496 37887 19499
rect 38286 19496 38292 19508
rect 37875 19468 38292 19496
rect 37875 19465 37887 19468
rect 37829 19459 37887 19465
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 39114 19496 39120 19508
rect 38488 19468 39120 19496
rect 33560 19400 36032 19428
rect 33560 19388 33566 19400
rect 37090 19388 37096 19440
rect 37148 19428 37154 19440
rect 38488 19428 38516 19468
rect 39114 19456 39120 19468
rect 39172 19456 39178 19508
rect 39294 19499 39352 19505
rect 39294 19465 39306 19499
rect 39340 19496 39352 19499
rect 40126 19496 40132 19508
rect 39340 19468 40132 19496
rect 39340 19465 39352 19468
rect 39294 19459 39352 19465
rect 40126 19456 40132 19468
rect 40184 19456 40190 19508
rect 41874 19456 41880 19508
rect 41932 19456 41938 19508
rect 37148 19400 38516 19428
rect 37148 19388 37154 19400
rect 32122 19360 32128 19372
rect 31726 19332 32128 19360
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 32401 19363 32459 19369
rect 32401 19329 32413 19363
rect 32447 19329 32459 19363
rect 32401 19323 32459 19329
rect 24636 19264 24900 19292
rect 24636 19252 24642 19264
rect 28534 19252 28540 19304
rect 28592 19252 28598 19304
rect 28994 19252 29000 19304
rect 29052 19292 29058 19304
rect 30006 19292 30012 19304
rect 29052 19264 30012 19292
rect 29052 19252 29058 19264
rect 30006 19252 30012 19264
rect 30064 19292 30070 19304
rect 30101 19295 30159 19301
rect 30101 19292 30113 19295
rect 30064 19264 30113 19292
rect 30064 19252 30070 19264
rect 30101 19261 30113 19264
rect 30147 19292 30159 19295
rect 32416 19292 32444 19323
rect 33042 19320 33048 19372
rect 33100 19360 33106 19372
rect 34054 19369 34060 19372
rect 33229 19363 33287 19369
rect 33229 19360 33241 19363
rect 33100 19332 33241 19360
rect 33100 19320 33106 19332
rect 33229 19329 33241 19332
rect 33275 19360 33287 19363
rect 33781 19363 33839 19369
rect 33781 19360 33793 19363
rect 33275 19332 33793 19360
rect 33275 19329 33287 19332
rect 33229 19323 33287 19329
rect 33781 19329 33793 19332
rect 33827 19329 33839 19363
rect 33781 19323 33839 19329
rect 34048 19323 34060 19369
rect 34054 19320 34060 19323
rect 34112 19320 34118 19372
rect 35805 19363 35863 19369
rect 35805 19329 35817 19363
rect 35851 19360 35863 19363
rect 35986 19360 35992 19372
rect 35851 19332 35992 19360
rect 35851 19329 35863 19332
rect 35805 19323 35863 19329
rect 35986 19320 35992 19332
rect 36044 19360 36050 19372
rect 37461 19363 37519 19369
rect 36044 19332 37228 19360
rect 36044 19320 36050 19332
rect 37200 19304 37228 19332
rect 37461 19329 37473 19363
rect 37507 19360 37519 19363
rect 37734 19360 37740 19372
rect 37507 19332 37740 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 37734 19320 37740 19332
rect 37792 19320 37798 19372
rect 38488 19369 38516 19400
rect 38562 19388 38568 19440
rect 38620 19428 38626 19440
rect 39666 19428 39672 19440
rect 38620 19400 39672 19428
rect 38620 19388 38626 19400
rect 39666 19388 39672 19400
rect 39724 19388 39730 19440
rect 39942 19388 39948 19440
rect 40000 19388 40006 19440
rect 38473 19363 38531 19369
rect 38473 19329 38485 19363
rect 38519 19329 38531 19363
rect 38473 19323 38531 19329
rect 38657 19363 38715 19369
rect 38657 19329 38669 19363
rect 38703 19360 38715 19363
rect 39022 19360 39028 19372
rect 38703 19332 39028 19360
rect 38703 19329 38715 19332
rect 38657 19323 38715 19329
rect 39022 19320 39028 19332
rect 39080 19320 39086 19372
rect 39117 19363 39175 19369
rect 39117 19329 39129 19363
rect 39163 19329 39175 19363
rect 39117 19323 39175 19329
rect 30147 19264 32444 19292
rect 30147 19261 30159 19264
rect 30101 19255 30159 19261
rect 35894 19252 35900 19304
rect 35952 19292 35958 19304
rect 36541 19295 36599 19301
rect 36541 19292 36553 19295
rect 35952 19264 36553 19292
rect 35952 19252 35958 19264
rect 36541 19261 36553 19264
rect 36587 19261 36599 19295
rect 36541 19255 36599 19261
rect 37182 19252 37188 19304
rect 37240 19292 37246 19304
rect 37553 19295 37611 19301
rect 37553 19292 37565 19295
rect 37240 19264 37565 19292
rect 37240 19252 37246 19264
rect 37553 19261 37565 19264
rect 37599 19261 37611 19295
rect 37553 19255 37611 19261
rect 38930 19252 38936 19304
rect 38988 19292 38994 19304
rect 39132 19292 39160 19323
rect 39206 19320 39212 19372
rect 39264 19320 39270 19372
rect 39298 19320 39304 19372
rect 39356 19360 39362 19372
rect 39393 19363 39451 19369
rect 39393 19360 39405 19363
rect 39356 19332 39405 19360
rect 39356 19320 39362 19332
rect 39393 19329 39405 19332
rect 39439 19329 39451 19363
rect 39393 19323 39451 19329
rect 39841 19363 39899 19369
rect 39841 19329 39853 19363
rect 39887 19329 39899 19363
rect 39841 19323 39899 19329
rect 38988 19264 39160 19292
rect 38988 19252 38994 19264
rect 39666 19252 39672 19304
rect 39724 19292 39730 19304
rect 39868 19292 39896 19323
rect 39724 19264 39896 19292
rect 39960 19292 39988 19388
rect 40037 19363 40095 19369
rect 40037 19329 40049 19363
rect 40083 19360 40095 19363
rect 40126 19360 40132 19372
rect 40083 19332 40132 19360
rect 40083 19329 40095 19332
rect 40037 19323 40095 19329
rect 40126 19320 40132 19332
rect 40184 19320 40190 19372
rect 40678 19320 40684 19372
rect 40736 19320 40742 19372
rect 40770 19320 40776 19372
rect 40828 19320 40834 19372
rect 40957 19363 41015 19369
rect 40957 19329 40969 19363
rect 41003 19360 41015 19363
rect 41046 19360 41052 19372
rect 41003 19332 41052 19360
rect 41003 19329 41015 19332
rect 40957 19323 41015 19329
rect 41046 19320 41052 19332
rect 41104 19360 41110 19372
rect 41969 19363 42027 19369
rect 41969 19360 41981 19363
rect 41104 19332 41981 19360
rect 41104 19320 41110 19332
rect 41969 19329 41981 19332
rect 42015 19360 42027 19363
rect 42242 19360 42248 19372
rect 42015 19332 42248 19360
rect 42015 19329 42027 19332
rect 41969 19323 42027 19329
rect 42242 19320 42248 19332
rect 42300 19320 42306 19372
rect 40310 19292 40316 19304
rect 39960 19264 40316 19292
rect 39724 19252 39730 19264
rect 40310 19252 40316 19264
rect 40368 19292 40374 19304
rect 42613 19295 42671 19301
rect 42613 19292 42625 19295
rect 40368 19264 42625 19292
rect 40368 19252 40374 19264
rect 42613 19261 42625 19264
rect 42659 19292 42671 19295
rect 43165 19295 43223 19301
rect 43165 19292 43177 19295
rect 42659 19264 43177 19292
rect 42659 19261 42671 19264
rect 42613 19255 42671 19261
rect 43165 19261 43177 19264
rect 43211 19261 43223 19295
rect 43165 19255 43223 19261
rect 21266 19224 21272 19236
rect 19904 19196 21272 19224
rect 21266 19184 21272 19196
rect 21324 19184 21330 19236
rect 31754 19184 31760 19236
rect 31812 19224 31818 19236
rect 32306 19224 32312 19236
rect 31812 19196 32312 19224
rect 31812 19184 31818 19196
rect 32306 19184 32312 19196
rect 32364 19184 32370 19236
rect 38657 19227 38715 19233
rect 38657 19193 38669 19227
rect 38703 19224 38715 19227
rect 39758 19224 39764 19236
rect 38703 19196 39764 19224
rect 38703 19193 38715 19196
rect 38657 19187 38715 19193
rect 39758 19184 39764 19196
rect 39816 19184 39822 19236
rect 40034 19184 40040 19236
rect 40092 19184 40098 19236
rect 19334 19116 19340 19168
rect 19392 19116 19398 19168
rect 28997 19159 29055 19165
rect 28997 19125 29009 19159
rect 29043 19156 29055 19159
rect 29086 19156 29092 19168
rect 29043 19128 29092 19156
rect 29043 19125 29055 19128
rect 28997 19119 29055 19125
rect 29086 19116 29092 19128
rect 29144 19116 29150 19168
rect 37642 19116 37648 19168
rect 37700 19116 37706 19168
rect 40954 19116 40960 19168
rect 41012 19116 41018 19168
rect 1104 19066 43884 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 43884 19066
rect 1104 18992 43884 19014
rect 15194 18912 15200 18964
rect 15252 18912 15258 18964
rect 21082 18912 21088 18964
rect 21140 18952 21146 18964
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 21140 18924 21281 18952
rect 21140 18912 21146 18924
rect 21269 18921 21281 18924
rect 21315 18921 21327 18955
rect 21269 18915 21327 18921
rect 22557 18955 22615 18961
rect 22557 18921 22569 18955
rect 22603 18952 22615 18955
rect 23842 18952 23848 18964
rect 22603 18924 23848 18952
rect 22603 18921 22615 18924
rect 22557 18915 22615 18921
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 18012 18788 18337 18816
rect 18012 18776 18018 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 21821 18819 21879 18825
rect 21821 18816 21833 18819
rect 21324 18788 21833 18816
rect 21324 18776 21330 18788
rect 21821 18785 21833 18788
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17034 18748 17040 18760
rect 16899 18720 17040 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 15378 18640 15384 18692
rect 15436 18680 15442 18692
rect 17604 18680 17632 18711
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 19150 18708 19156 18760
rect 19208 18748 19214 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19208 18720 19441 18748
rect 19208 18708 19214 18720
rect 19429 18717 19441 18720
rect 19475 18748 19487 18751
rect 20714 18748 20720 18760
rect 19475 18720 20720 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21634 18708 21640 18760
rect 21692 18708 21698 18760
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 22646 18748 22652 18760
rect 21775 18720 22652 18748
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 23124 18757 23152 18924
rect 23842 18912 23848 18924
rect 23900 18952 23906 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 23900 18924 24593 18952
rect 23900 18912 23906 18924
rect 24581 18921 24593 18924
rect 24627 18952 24639 18955
rect 28994 18952 29000 18964
rect 24627 18924 29000 18952
rect 24627 18921 24639 18924
rect 24581 18915 24639 18921
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 31113 18955 31171 18961
rect 31113 18952 31125 18955
rect 29104 18924 31125 18952
rect 28077 18887 28135 18893
rect 28077 18853 28089 18887
rect 28123 18884 28135 18887
rect 28350 18884 28356 18896
rect 28123 18856 28356 18884
rect 28123 18853 28135 18856
rect 28077 18847 28135 18853
rect 28350 18844 28356 18856
rect 28408 18844 28414 18896
rect 29104 18884 29132 18924
rect 31113 18921 31125 18924
rect 31159 18952 31171 18955
rect 31202 18952 31208 18964
rect 31159 18924 31208 18952
rect 31159 18921 31171 18924
rect 31113 18915 31171 18921
rect 31202 18912 31208 18924
rect 31260 18912 31266 18964
rect 34054 18912 34060 18964
rect 34112 18952 34118 18964
rect 34241 18955 34299 18961
rect 34241 18952 34253 18955
rect 34112 18924 34253 18952
rect 34112 18912 34118 18924
rect 34241 18921 34253 18924
rect 34287 18921 34299 18955
rect 34241 18915 34299 18921
rect 34977 18955 35035 18961
rect 34977 18921 34989 18955
rect 35023 18952 35035 18955
rect 35526 18952 35532 18964
rect 35023 18924 35532 18952
rect 35023 18921 35035 18924
rect 34977 18915 35035 18921
rect 35526 18912 35532 18924
rect 35584 18912 35590 18964
rect 35618 18912 35624 18964
rect 35676 18912 35682 18964
rect 36446 18912 36452 18964
rect 36504 18952 36510 18964
rect 36541 18955 36599 18961
rect 36541 18952 36553 18955
rect 36504 18924 36553 18952
rect 36504 18912 36510 18924
rect 36541 18921 36553 18924
rect 36587 18921 36599 18955
rect 36541 18915 36599 18921
rect 36906 18912 36912 18964
rect 36964 18912 36970 18964
rect 37550 18912 37556 18964
rect 37608 18912 37614 18964
rect 37918 18912 37924 18964
rect 37976 18952 37982 18964
rect 38013 18955 38071 18961
rect 38013 18952 38025 18955
rect 37976 18924 38025 18952
rect 37976 18912 37982 18924
rect 38013 18921 38025 18924
rect 38059 18921 38071 18955
rect 38013 18915 38071 18921
rect 39298 18912 39304 18964
rect 39356 18912 39362 18964
rect 40221 18955 40279 18961
rect 40221 18921 40233 18955
rect 40267 18952 40279 18955
rect 40678 18952 40684 18964
rect 40267 18924 40684 18952
rect 40267 18921 40279 18924
rect 40221 18915 40279 18921
rect 40678 18912 40684 18924
rect 40736 18912 40742 18964
rect 40770 18912 40776 18964
rect 40828 18952 40834 18964
rect 41782 18952 41788 18964
rect 40828 18924 41788 18952
rect 40828 18912 40834 18924
rect 41782 18912 41788 18924
rect 41840 18952 41846 18964
rect 43073 18955 43131 18961
rect 43073 18952 43085 18955
rect 41840 18924 43085 18952
rect 41840 18912 41846 18924
rect 43073 18921 43085 18924
rect 43119 18921 43131 18955
rect 43073 18915 43131 18921
rect 28920 18856 29132 18884
rect 28810 18816 28816 18828
rect 28644 18788 28816 18816
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18717 23167 18751
rect 23109 18711 23167 18717
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18748 23995 18751
rect 24578 18748 24584 18760
rect 23983 18720 24584 18748
rect 23983 18717 23995 18720
rect 23937 18711 23995 18717
rect 19242 18680 19248 18692
rect 15436 18652 19248 18680
rect 15436 18640 15442 18652
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 19674 18683 19732 18689
rect 19674 18680 19686 18683
rect 19444 18652 19686 18680
rect 19444 18624 19472 18652
rect 19674 18649 19686 18652
rect 19720 18649 19732 18683
rect 19674 18643 19732 18649
rect 22002 18640 22008 18692
rect 22060 18680 22066 18692
rect 23124 18680 23152 18711
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 28644 18757 28672 18788
rect 28810 18776 28816 18788
rect 28868 18776 28874 18828
rect 28920 18757 28948 18856
rect 37366 18844 37372 18896
rect 37424 18884 37430 18896
rect 38838 18884 38844 18896
rect 37424 18856 38844 18884
rect 37424 18844 37430 18856
rect 38838 18844 38844 18856
rect 38896 18884 38902 18896
rect 39666 18884 39672 18896
rect 38896 18856 39672 18884
rect 38896 18844 38902 18856
rect 39666 18844 39672 18856
rect 39724 18844 39730 18896
rect 32968 18788 40172 18816
rect 32968 18760 32996 18788
rect 26964 18751 27022 18757
rect 26964 18717 26976 18751
rect 27010 18748 27022 18751
rect 28629 18751 28687 18757
rect 27010 18720 28028 18748
rect 27010 18717 27022 18720
rect 26964 18711 27022 18717
rect 22060 18652 23152 18680
rect 22060 18640 22066 18652
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18612 17095 18615
rect 17126 18612 17132 18624
rect 17083 18584 17132 18612
rect 17083 18581 17095 18584
rect 17037 18575 17095 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 19426 18572 19432 18624
rect 19484 18572 19490 18624
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20809 18615 20867 18621
rect 20809 18612 20821 18615
rect 20036 18584 20821 18612
rect 20036 18572 20042 18584
rect 20809 18581 20821 18584
rect 20855 18581 20867 18615
rect 28000 18612 28028 18720
rect 28629 18717 28641 18751
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 28905 18751 28963 18757
rect 28905 18717 28917 18751
rect 28951 18717 28963 18751
rect 28905 18711 28963 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29178 18748 29184 18760
rect 29043 18720 29184 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29178 18708 29184 18720
rect 29236 18748 29242 18760
rect 29454 18748 29460 18760
rect 29236 18720 29460 18748
rect 29236 18708 29242 18720
rect 29454 18708 29460 18720
rect 29512 18708 29518 18760
rect 29546 18708 29552 18760
rect 29604 18748 29610 18760
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 29604 18720 29745 18748
rect 29604 18708 29610 18720
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 32766 18708 32772 18760
rect 32824 18757 32830 18760
rect 32824 18748 32836 18757
rect 32824 18720 32869 18748
rect 32824 18711 32836 18720
rect 32824 18708 32830 18711
rect 32950 18708 32956 18760
rect 33008 18708 33014 18760
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18748 33103 18751
rect 33594 18748 33600 18760
rect 33091 18720 33600 18748
rect 33091 18717 33103 18720
rect 33045 18711 33103 18717
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 33689 18751 33747 18757
rect 33689 18717 33701 18751
rect 33735 18748 33747 18751
rect 33735 18720 33824 18748
rect 33735 18717 33747 18720
rect 33689 18711 33747 18717
rect 28350 18640 28356 18692
rect 28408 18680 28414 18692
rect 28813 18683 28871 18689
rect 28813 18680 28825 18683
rect 28408 18652 28825 18680
rect 28408 18640 28414 18652
rect 28813 18649 28825 18652
rect 28859 18649 28871 18683
rect 29978 18683 30036 18689
rect 29978 18680 29990 18683
rect 28813 18643 28871 18649
rect 29196 18652 29990 18680
rect 29086 18612 29092 18624
rect 28000 18584 29092 18612
rect 20809 18575 20867 18581
rect 29086 18572 29092 18584
rect 29144 18572 29150 18624
rect 29196 18621 29224 18652
rect 29978 18649 29990 18652
rect 30024 18649 30036 18683
rect 29978 18643 30036 18649
rect 31018 18640 31024 18692
rect 31076 18680 31082 18692
rect 33796 18680 33824 18720
rect 33962 18708 33968 18760
rect 34020 18708 34026 18760
rect 34072 18757 34100 18788
rect 40144 18760 40172 18788
rect 40218 18776 40224 18828
rect 40276 18816 40282 18828
rect 41601 18819 41659 18825
rect 41601 18816 41613 18819
rect 40276 18788 41613 18816
rect 40276 18776 40282 18788
rect 41601 18785 41613 18788
rect 41647 18785 41659 18819
rect 41601 18779 41659 18785
rect 34057 18751 34115 18757
rect 34057 18717 34069 18751
rect 34103 18717 34115 18751
rect 34057 18711 34115 18717
rect 35437 18751 35495 18757
rect 35437 18717 35449 18751
rect 35483 18717 35495 18751
rect 35437 18711 35495 18717
rect 31076 18652 33824 18680
rect 31076 18640 31082 18652
rect 29181 18615 29239 18621
rect 29181 18581 29193 18615
rect 29227 18581 29239 18615
rect 29181 18575 29239 18581
rect 31665 18615 31723 18621
rect 31665 18581 31677 18615
rect 31711 18612 31723 18615
rect 32582 18612 32588 18624
rect 31711 18584 32588 18612
rect 31711 18581 31723 18584
rect 31665 18575 31723 18581
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 33796 18612 33824 18652
rect 33873 18683 33931 18689
rect 33873 18649 33885 18683
rect 33919 18680 33931 18683
rect 34790 18680 34796 18692
rect 33919 18652 34796 18680
rect 33919 18649 33931 18652
rect 33873 18643 33931 18649
rect 34790 18640 34796 18652
rect 34848 18640 34854 18692
rect 35452 18680 35480 18711
rect 35618 18708 35624 18760
rect 35676 18708 35682 18760
rect 36817 18751 36875 18757
rect 36817 18717 36829 18751
rect 36863 18717 36875 18751
rect 36817 18711 36875 18717
rect 36909 18751 36967 18757
rect 36909 18717 36921 18751
rect 36955 18748 36967 18751
rect 37090 18748 37096 18760
rect 36955 18720 37096 18748
rect 36955 18717 36967 18720
rect 36909 18711 36967 18717
rect 35986 18680 35992 18692
rect 35452 18652 35992 18680
rect 35986 18640 35992 18652
rect 36044 18640 36050 18692
rect 36832 18680 36860 18711
rect 37090 18708 37096 18720
rect 37148 18708 37154 18760
rect 37366 18708 37372 18760
rect 37424 18708 37430 18760
rect 37550 18708 37556 18760
rect 37608 18748 37614 18760
rect 37918 18748 37924 18760
rect 37608 18720 37924 18748
rect 37608 18708 37614 18720
rect 37918 18708 37924 18720
rect 37976 18708 37982 18760
rect 40126 18708 40132 18760
rect 40184 18708 40190 18760
rect 40313 18751 40371 18757
rect 40313 18717 40325 18751
rect 40359 18748 40371 18751
rect 41690 18748 41696 18760
rect 40359 18720 41696 18748
rect 40359 18717 40371 18720
rect 40313 18711 40371 18717
rect 41690 18708 41696 18720
rect 41748 18708 41754 18760
rect 42610 18708 42616 18760
rect 42668 18708 42674 18760
rect 37734 18680 37740 18692
rect 36832 18652 37740 18680
rect 37734 18640 37740 18652
rect 37792 18640 37798 18692
rect 38654 18640 38660 18692
rect 38712 18680 38718 18692
rect 38749 18683 38807 18689
rect 38749 18680 38761 18683
rect 38712 18652 38761 18680
rect 38712 18640 38718 18652
rect 38749 18649 38761 18652
rect 38795 18680 38807 18683
rect 39942 18680 39948 18692
rect 38795 18652 39948 18680
rect 38795 18649 38807 18652
rect 38749 18643 38807 18649
rect 39942 18640 39948 18652
rect 40000 18640 40006 18692
rect 40770 18640 40776 18692
rect 40828 18640 40834 18692
rect 40957 18683 41015 18689
rect 40957 18649 40969 18683
rect 41003 18680 41015 18683
rect 41046 18680 41052 18692
rect 41003 18652 41052 18680
rect 41003 18649 41015 18652
rect 40957 18643 41015 18649
rect 41046 18640 41052 18652
rect 41104 18640 41110 18692
rect 34698 18612 34704 18624
rect 33796 18584 34704 18612
rect 34698 18572 34704 18584
rect 34756 18572 34762 18624
rect 36354 18572 36360 18624
rect 36412 18612 36418 18624
rect 38930 18612 38936 18624
rect 36412 18584 38936 18612
rect 36412 18572 36418 18584
rect 38930 18572 38936 18584
rect 38988 18572 38994 18624
rect 39022 18572 39028 18624
rect 39080 18572 39086 18624
rect 39114 18572 39120 18624
rect 39172 18572 39178 18624
rect 41138 18572 41144 18624
rect 41196 18572 41202 18624
rect 42242 18572 42248 18624
rect 42300 18612 42306 18624
rect 42429 18615 42487 18621
rect 42429 18612 42441 18615
rect 42300 18584 42441 18612
rect 42300 18572 42306 18584
rect 42429 18581 42441 18584
rect 42475 18581 42487 18615
rect 42429 18575 42487 18581
rect 1104 18522 43884 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 43884 18522
rect 1104 18448 43884 18470
rect 15286 18408 15292 18420
rect 14660 18380 15292 18408
rect 14660 18349 14688 18380
rect 15286 18368 15292 18380
rect 15344 18408 15350 18420
rect 15746 18408 15752 18420
rect 15344 18380 15752 18408
rect 15344 18368 15350 18380
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 19889 18411 19947 18417
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 19978 18408 19984 18420
rect 19935 18380 19984 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 22373 18411 22431 18417
rect 22373 18377 22385 18411
rect 22419 18408 22431 18411
rect 22554 18408 22560 18420
rect 22419 18380 22560 18408
rect 22419 18377 22431 18380
rect 22373 18371 22431 18377
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 25038 18368 25044 18420
rect 25096 18408 25102 18420
rect 27614 18408 27620 18420
rect 25096 18380 27620 18408
rect 25096 18368 25102 18380
rect 27614 18368 27620 18380
rect 27672 18368 27678 18420
rect 32306 18368 32312 18420
rect 32364 18408 32370 18420
rect 32401 18411 32459 18417
rect 32401 18408 32413 18411
rect 32364 18380 32413 18408
rect 32364 18368 32370 18380
rect 32401 18377 32413 18380
rect 32447 18377 32459 18411
rect 32401 18371 32459 18377
rect 34606 18368 34612 18420
rect 34664 18408 34670 18420
rect 35069 18411 35127 18417
rect 35069 18408 35081 18411
rect 34664 18380 35081 18408
rect 34664 18368 34670 18380
rect 35069 18377 35081 18380
rect 35115 18377 35127 18411
rect 35069 18371 35127 18377
rect 36173 18411 36231 18417
rect 36173 18377 36185 18411
rect 36219 18408 36231 18411
rect 36446 18408 36452 18420
rect 36219 18380 36452 18408
rect 36219 18377 36231 18380
rect 36173 18371 36231 18377
rect 36446 18368 36452 18380
rect 36504 18368 36510 18420
rect 37458 18368 37464 18420
rect 37516 18408 37522 18420
rect 37737 18411 37795 18417
rect 37737 18408 37749 18411
rect 37516 18380 37749 18408
rect 37516 18368 37522 18380
rect 37737 18377 37749 18380
rect 37783 18408 37795 18411
rect 38010 18408 38016 18420
rect 37783 18380 38016 18408
rect 37783 18377 37795 18380
rect 37737 18371 37795 18377
rect 38010 18368 38016 18380
rect 38068 18368 38074 18420
rect 38197 18411 38255 18417
rect 38197 18377 38209 18411
rect 38243 18408 38255 18411
rect 39022 18408 39028 18420
rect 38243 18380 39028 18408
rect 38243 18377 38255 18380
rect 38197 18371 38255 18377
rect 39022 18368 39028 18380
rect 39080 18368 39086 18420
rect 39206 18368 39212 18420
rect 39264 18408 39270 18420
rect 40037 18411 40095 18417
rect 40037 18408 40049 18411
rect 39264 18380 40049 18408
rect 39264 18368 39270 18380
rect 40037 18377 40049 18380
rect 40083 18377 40095 18411
rect 40037 18371 40095 18377
rect 42610 18368 42616 18420
rect 42668 18368 42674 18420
rect 14645 18343 14703 18349
rect 14645 18309 14657 18343
rect 14691 18309 14703 18343
rect 14645 18303 14703 18309
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 20254 18340 20260 18352
rect 15436 18312 15792 18340
rect 15436 18300 15442 18312
rect 15764 18284 15792 18312
rect 19904 18312 20260 18340
rect 19904 18284 19932 18312
rect 20254 18300 20260 18312
rect 20312 18340 20318 18352
rect 23474 18340 23480 18352
rect 20312 18312 23480 18340
rect 20312 18300 20318 18312
rect 23474 18300 23480 18312
rect 23532 18340 23538 18352
rect 23845 18343 23903 18349
rect 23845 18340 23857 18343
rect 23532 18312 23857 18340
rect 23532 18300 23538 18312
rect 23845 18309 23857 18312
rect 23891 18309 23903 18343
rect 23845 18303 23903 18309
rect 28994 18300 29000 18352
rect 29052 18340 29058 18352
rect 30742 18340 30748 18352
rect 29052 18312 30748 18340
rect 29052 18300 29058 18312
rect 30742 18300 30748 18312
rect 30800 18340 30806 18352
rect 31478 18340 31484 18352
rect 30800 18312 31484 18340
rect 30800 18300 30806 18312
rect 31478 18300 31484 18312
rect 31536 18340 31542 18352
rect 33042 18340 33048 18352
rect 31536 18312 33048 18340
rect 31536 18300 31542 18312
rect 33042 18300 33048 18312
rect 33100 18300 33106 18352
rect 35618 18300 35624 18352
rect 35676 18340 35682 18352
rect 37918 18349 37924 18352
rect 37829 18343 37887 18349
rect 37829 18340 37841 18343
rect 35676 18312 37841 18340
rect 35676 18300 35682 18312
rect 37829 18309 37841 18312
rect 37875 18309 37887 18343
rect 37829 18303 37887 18309
rect 37915 18303 37924 18349
rect 37976 18340 37982 18352
rect 39853 18343 39911 18349
rect 39853 18340 39865 18343
rect 37976 18312 38015 18340
rect 38672 18312 39865 18340
rect 37918 18300 37924 18303
rect 37976 18300 37982 18312
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15562 18272 15568 18284
rect 15519 18244 15568 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15562 18232 15568 18244
rect 15620 18232 15626 18284
rect 15654 18232 15660 18284
rect 15712 18232 15718 18284
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 17405 18275 17463 18281
rect 17405 18272 17417 18275
rect 15841 18235 15899 18241
rect 16132 18244 17417 18272
rect 14918 18164 14924 18216
rect 14976 18204 14982 18216
rect 15856 18204 15884 18235
rect 16132 18213 16160 18244
rect 17405 18241 17417 18244
rect 17451 18241 17463 18275
rect 17405 18235 17463 18241
rect 17862 18232 17868 18284
rect 17920 18232 17926 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18012 18244 18245 18272
rect 18012 18232 18018 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18598 18232 18604 18284
rect 18656 18232 18662 18284
rect 18690 18232 18696 18284
rect 18748 18232 18754 18284
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19300 18244 19809 18272
rect 19300 18232 19306 18244
rect 19797 18241 19809 18244
rect 19843 18272 19855 18275
rect 19886 18272 19892 18284
rect 19843 18244 19892 18272
rect 19843 18241 19855 18244
rect 19797 18235 19855 18241
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20073 18275 20131 18281
rect 20073 18241 20085 18275
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 20806 18272 20812 18284
rect 20763 18244 20812 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 14976 18176 15884 18204
rect 16117 18207 16175 18213
rect 14976 18164 14982 18176
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 18138 18164 18144 18216
rect 18196 18164 18202 18216
rect 20088 18204 20116 18235
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 20898 18232 20904 18284
rect 20956 18232 20962 18284
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21082 18272 21088 18284
rect 21039 18244 21088 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 22738 18232 22744 18284
rect 22796 18232 22802 18284
rect 23569 18275 23627 18281
rect 23569 18241 23581 18275
rect 23615 18272 23627 18275
rect 23750 18272 23756 18284
rect 23615 18244 23756 18272
rect 23615 18241 23627 18244
rect 23569 18235 23627 18241
rect 20088 18176 21036 18204
rect 21008 18148 21036 18176
rect 22830 18164 22836 18216
rect 22888 18164 22894 18216
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23584 18204 23612 18235
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 26165 18275 26223 18281
rect 26165 18241 26177 18275
rect 26211 18272 26223 18275
rect 27430 18272 27436 18284
rect 26211 18244 27436 18272
rect 26211 18241 26223 18244
rect 26165 18235 26223 18241
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 29914 18281 29920 18284
rect 29908 18235 29920 18281
rect 29914 18232 29920 18235
rect 29972 18232 29978 18284
rect 32309 18275 32367 18281
rect 32309 18241 32321 18275
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 32493 18275 32551 18281
rect 32493 18241 32505 18275
rect 32539 18272 32551 18275
rect 32582 18272 32588 18284
rect 32539 18244 32588 18272
rect 32539 18241 32551 18244
rect 32493 18235 32551 18241
rect 22980 18176 23612 18204
rect 26421 18207 26479 18213
rect 22980 18164 22986 18176
rect 26421 18173 26433 18207
rect 26467 18204 26479 18207
rect 26694 18204 26700 18216
rect 26467 18176 26700 18204
rect 26467 18173 26479 18176
rect 26421 18167 26479 18173
rect 26694 18164 26700 18176
rect 26752 18204 26758 18216
rect 27154 18204 27160 18216
rect 26752 18176 27160 18204
rect 26752 18164 26758 18176
rect 27154 18164 27160 18176
rect 27212 18204 27218 18216
rect 28169 18207 28227 18213
rect 28169 18204 28181 18207
rect 27212 18176 28181 18204
rect 27212 18164 27218 18176
rect 28169 18173 28181 18176
rect 28215 18204 28227 18207
rect 28534 18204 28540 18216
rect 28215 18176 28540 18204
rect 28215 18173 28227 18176
rect 28169 18167 28227 18173
rect 28534 18164 28540 18176
rect 28592 18164 28598 18216
rect 29546 18164 29552 18216
rect 29604 18204 29610 18216
rect 29641 18207 29699 18213
rect 29641 18204 29653 18207
rect 29604 18176 29653 18204
rect 29604 18164 29610 18176
rect 29641 18173 29653 18176
rect 29687 18173 29699 18207
rect 29641 18167 29699 18173
rect 31938 18164 31944 18216
rect 31996 18204 32002 18216
rect 32324 18204 32352 18235
rect 32582 18232 32588 18244
rect 32640 18232 32646 18284
rect 34422 18232 34428 18284
rect 34480 18232 34486 18284
rect 34609 18275 34667 18281
rect 34609 18241 34621 18275
rect 34655 18272 34667 18275
rect 34698 18272 34704 18284
rect 34655 18244 34704 18272
rect 34655 18241 34667 18244
rect 34609 18235 34667 18241
rect 34698 18232 34704 18244
rect 34756 18232 34762 18284
rect 37461 18275 37519 18281
rect 37461 18241 37473 18275
rect 37507 18272 37519 18275
rect 37734 18272 37740 18284
rect 37507 18244 37740 18272
rect 37507 18241 37519 18244
rect 37461 18235 37519 18241
rect 37734 18232 37740 18244
rect 37792 18272 37798 18284
rect 38672 18281 38700 18312
rect 39853 18309 39865 18312
rect 39899 18309 39911 18343
rect 39853 18303 39911 18309
rect 40856 18343 40914 18349
rect 40856 18309 40868 18343
rect 40902 18340 40914 18343
rect 40954 18340 40960 18352
rect 40902 18312 40960 18340
rect 40902 18309 40914 18312
rect 40856 18303 40914 18309
rect 40954 18300 40960 18312
rect 41012 18300 41018 18352
rect 38657 18275 38715 18281
rect 38657 18272 38669 18275
rect 37792 18244 38669 18272
rect 37792 18232 37798 18244
rect 38657 18241 38669 18244
rect 38703 18241 38715 18275
rect 38657 18235 38715 18241
rect 38749 18275 38807 18281
rect 38749 18241 38761 18275
rect 38795 18272 38807 18275
rect 38838 18272 38844 18284
rect 38795 18244 38844 18272
rect 38795 18241 38807 18244
rect 38749 18235 38807 18241
rect 38838 18232 38844 18244
rect 38896 18232 38902 18284
rect 38933 18275 38991 18281
rect 38933 18241 38945 18275
rect 38979 18241 38991 18275
rect 38933 18235 38991 18241
rect 39025 18275 39083 18281
rect 39025 18241 39037 18275
rect 39071 18272 39083 18275
rect 39206 18272 39212 18284
rect 39071 18244 39212 18272
rect 39071 18241 39083 18244
rect 39025 18235 39083 18241
rect 32950 18204 32956 18216
rect 31996 18176 32956 18204
rect 31996 18164 32002 18176
rect 32950 18164 32956 18176
rect 33008 18164 33014 18216
rect 33594 18164 33600 18216
rect 33652 18204 33658 18216
rect 33781 18207 33839 18213
rect 33781 18204 33793 18207
rect 33652 18176 33793 18204
rect 33652 18164 33658 18176
rect 33781 18173 33793 18176
rect 33827 18204 33839 18207
rect 33827 18176 37412 18204
rect 33827 18173 33839 18176
rect 33781 18167 33839 18173
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20119 18108 20944 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15470 18068 15476 18080
rect 15059 18040 15476 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 20530 18028 20536 18080
rect 20588 18028 20594 18080
rect 20916 18068 20944 18108
rect 20990 18096 20996 18148
rect 21048 18096 21054 18148
rect 32490 18096 32496 18148
rect 32548 18136 32554 18148
rect 34422 18136 34428 18148
rect 32548 18108 34428 18136
rect 32548 18096 32554 18108
rect 34422 18096 34428 18108
rect 34480 18096 34486 18148
rect 35710 18096 35716 18148
rect 35768 18136 35774 18148
rect 35805 18139 35863 18145
rect 35805 18136 35817 18139
rect 35768 18108 35817 18136
rect 35768 18096 35774 18108
rect 35805 18105 35817 18108
rect 35851 18105 35863 18139
rect 35805 18099 35863 18105
rect 36354 18096 36360 18148
rect 36412 18096 36418 18148
rect 37384 18136 37412 18176
rect 37550 18164 37556 18216
rect 37608 18204 37614 18216
rect 38948 18204 38976 18235
rect 39206 18232 39212 18244
rect 39264 18272 39270 18284
rect 39669 18275 39727 18281
rect 39669 18272 39681 18275
rect 39264 18244 39681 18272
rect 39264 18232 39270 18244
rect 39669 18241 39681 18244
rect 39715 18241 39727 18275
rect 39669 18235 39727 18241
rect 42981 18275 43039 18281
rect 42981 18241 42993 18275
rect 43027 18272 43039 18275
rect 43530 18272 43536 18284
rect 43027 18244 43536 18272
rect 43027 18241 43039 18244
rect 42981 18235 43039 18241
rect 43530 18232 43536 18244
rect 43588 18232 43594 18284
rect 39298 18204 39304 18216
rect 37608 18176 39304 18204
rect 37608 18164 37614 18176
rect 39298 18164 39304 18176
rect 39356 18164 39362 18216
rect 40589 18207 40647 18213
rect 40589 18173 40601 18207
rect 40635 18173 40647 18207
rect 40589 18167 40647 18173
rect 40604 18136 40632 18167
rect 43070 18164 43076 18216
rect 43128 18164 43134 18216
rect 43165 18207 43223 18213
rect 43165 18173 43177 18207
rect 43211 18173 43223 18207
rect 43165 18167 43223 18173
rect 37384 18108 40632 18136
rect 21174 18068 21180 18080
rect 20916 18040 21180 18068
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 27617 18071 27675 18077
rect 27617 18037 27629 18071
rect 27663 18068 27675 18071
rect 28166 18068 28172 18080
rect 27663 18040 28172 18068
rect 27663 18037 27675 18040
rect 27617 18031 27675 18037
rect 28166 18028 28172 18040
rect 28224 18068 28230 18080
rect 28902 18068 28908 18080
rect 28224 18040 28908 18068
rect 28224 18028 28230 18040
rect 28902 18028 28908 18040
rect 28960 18028 28966 18080
rect 30650 18028 30656 18080
rect 30708 18068 30714 18080
rect 30926 18068 30932 18080
rect 30708 18040 30932 18068
rect 30708 18028 30714 18040
rect 30926 18028 30932 18040
rect 30984 18068 30990 18080
rect 31021 18071 31079 18077
rect 31021 18068 31033 18071
rect 30984 18040 31033 18068
rect 30984 18028 30990 18040
rect 31021 18037 31033 18040
rect 31067 18037 31079 18071
rect 31021 18031 31079 18037
rect 34514 18028 34520 18080
rect 34572 18028 34578 18080
rect 36170 18028 36176 18080
rect 36228 18028 36234 18080
rect 36909 18071 36967 18077
rect 36909 18037 36921 18071
rect 36955 18068 36967 18071
rect 37182 18068 37188 18080
rect 36955 18040 37188 18068
rect 36955 18037 36967 18040
rect 36909 18031 36967 18037
rect 37182 18028 37188 18040
rect 37240 18028 37246 18080
rect 37550 18028 37556 18080
rect 37608 18028 37614 18080
rect 38746 18028 38752 18080
rect 38804 18068 38810 18080
rect 39209 18071 39267 18077
rect 39209 18068 39221 18071
rect 38804 18040 39221 18068
rect 38804 18028 38810 18040
rect 39209 18037 39221 18040
rect 39255 18037 39267 18071
rect 40604 18068 40632 18108
rect 42978 18096 42984 18148
rect 43036 18136 43042 18148
rect 43180 18136 43208 18167
rect 43036 18108 43208 18136
rect 43036 18096 43042 18108
rect 41322 18068 41328 18080
rect 40604 18040 41328 18068
rect 39209 18031 39267 18037
rect 41322 18028 41328 18040
rect 41380 18028 41386 18080
rect 41690 18028 41696 18080
rect 41748 18068 41754 18080
rect 41969 18071 42027 18077
rect 41969 18068 41981 18071
rect 41748 18040 41981 18068
rect 41748 18028 41754 18040
rect 41969 18037 41981 18040
rect 42015 18037 42027 18071
rect 41969 18031 42027 18037
rect 1104 17978 43884 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 43884 17978
rect 1104 17904 43884 17926
rect 19886 17824 19892 17876
rect 19944 17824 19950 17876
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20070 17864 20076 17876
rect 20027 17836 20076 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20898 17824 20904 17876
rect 20956 17864 20962 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 20956 17836 21097 17864
rect 20956 17824 20962 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 21085 17827 21143 17833
rect 21100 17796 21128 17827
rect 22278 17824 22284 17876
rect 22336 17824 22342 17876
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 22940 17796 22968 17827
rect 23566 17824 23572 17876
rect 23624 17824 23630 17876
rect 24762 17864 24768 17876
rect 24596 17836 24768 17864
rect 23934 17796 23940 17808
rect 21100 17768 23940 17796
rect 23934 17756 23940 17768
rect 23992 17796 23998 17808
rect 24486 17796 24492 17808
rect 23992 17768 24492 17796
rect 23992 17756 23998 17768
rect 24486 17756 24492 17768
rect 24544 17756 24550 17808
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 13725 17731 13783 17737
rect 13725 17728 13737 17731
rect 13688 17700 13737 17728
rect 13688 17688 13694 17700
rect 13725 17697 13737 17700
rect 13771 17728 13783 17731
rect 14921 17731 14979 17737
rect 14921 17728 14933 17731
rect 13771 17700 14933 17728
rect 13771 17697 13783 17700
rect 13725 17691 13783 17697
rect 14921 17697 14933 17700
rect 14967 17728 14979 17731
rect 15010 17728 15016 17740
rect 14967 17700 15016 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 17310 17688 17316 17740
rect 17368 17688 17374 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20530 17728 20536 17740
rect 20119 17700 20536 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 24596 17728 24624 17836
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 25314 17824 25320 17876
rect 25372 17864 25378 17876
rect 25774 17864 25780 17876
rect 25372 17836 25780 17864
rect 25372 17824 25378 17836
rect 25774 17824 25780 17836
rect 25832 17864 25838 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 25832 17836 25973 17864
rect 25832 17824 25838 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 27430 17824 27436 17876
rect 27488 17824 27494 17876
rect 27890 17824 27896 17876
rect 27948 17864 27954 17876
rect 28445 17867 28503 17873
rect 28445 17864 28457 17867
rect 27948 17836 28457 17864
rect 27948 17824 27954 17836
rect 28445 17833 28457 17836
rect 28491 17833 28503 17867
rect 28445 17827 28503 17833
rect 28629 17867 28687 17873
rect 28629 17833 28641 17867
rect 28675 17864 28687 17867
rect 28810 17864 28816 17876
rect 28675 17836 28816 17864
rect 28675 17833 28687 17836
rect 28629 17827 28687 17833
rect 28810 17824 28816 17836
rect 28868 17824 28874 17876
rect 29825 17867 29883 17873
rect 29825 17833 29837 17867
rect 29871 17864 29883 17867
rect 29914 17864 29920 17876
rect 29871 17836 29920 17864
rect 29871 17833 29883 17836
rect 29825 17827 29883 17833
rect 29914 17824 29920 17836
rect 29972 17824 29978 17876
rect 31478 17824 31484 17876
rect 31536 17824 31542 17876
rect 33042 17824 33048 17876
rect 33100 17864 33106 17876
rect 33505 17867 33563 17873
rect 33505 17864 33517 17867
rect 33100 17836 33517 17864
rect 33100 17824 33106 17836
rect 33505 17833 33517 17836
rect 33551 17833 33563 17867
rect 33505 17827 33563 17833
rect 34333 17867 34391 17873
rect 34333 17833 34345 17867
rect 34379 17864 34391 17867
rect 34606 17864 34612 17876
rect 34379 17836 34612 17864
rect 34379 17833 34391 17836
rect 34333 17827 34391 17833
rect 34606 17824 34612 17836
rect 34664 17864 34670 17876
rect 35069 17867 35127 17873
rect 35069 17864 35081 17867
rect 34664 17836 35081 17864
rect 34664 17824 34670 17836
rect 35069 17833 35081 17836
rect 35115 17833 35127 17867
rect 35069 17827 35127 17833
rect 35802 17824 35808 17876
rect 35860 17824 35866 17876
rect 36262 17824 36268 17876
rect 36320 17864 36326 17876
rect 37642 17864 37648 17876
rect 36320 17836 37648 17864
rect 36320 17824 36326 17836
rect 37642 17824 37648 17836
rect 37700 17864 37706 17876
rect 37918 17864 37924 17876
rect 37700 17836 37924 17864
rect 37700 17824 37706 17836
rect 37918 17824 37924 17836
rect 37976 17824 37982 17876
rect 38933 17867 38991 17873
rect 38933 17833 38945 17867
rect 38979 17864 38991 17867
rect 39022 17864 39028 17876
rect 38979 17836 39028 17864
rect 38979 17833 38991 17836
rect 38933 17827 38991 17833
rect 39022 17824 39028 17836
rect 39080 17824 39086 17876
rect 40126 17824 40132 17876
rect 40184 17824 40190 17876
rect 41325 17867 41383 17873
rect 41325 17833 41337 17867
rect 41371 17864 41383 17867
rect 42978 17864 42984 17876
rect 41371 17836 42984 17864
rect 41371 17833 41383 17836
rect 41325 17827 41383 17833
rect 42978 17824 42984 17836
rect 43036 17824 43042 17876
rect 43070 17824 43076 17876
rect 43128 17864 43134 17876
rect 43349 17867 43407 17873
rect 43349 17864 43361 17867
rect 43128 17836 43361 17864
rect 43128 17824 43134 17836
rect 43349 17833 43361 17836
rect 43395 17833 43407 17867
rect 43349 17827 43407 17833
rect 27614 17756 27620 17808
rect 27672 17756 27678 17808
rect 29454 17756 29460 17808
rect 29512 17796 29518 17808
rect 31938 17796 31944 17808
rect 29512 17768 31944 17796
rect 29512 17756 29518 17768
rect 21376 17700 24624 17728
rect 27632 17728 27660 17756
rect 27632 17700 27752 17728
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 15746 17620 15752 17672
rect 15804 17620 15810 17672
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17218 17660 17224 17672
rect 17175 17632 17224 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 16117 17595 16175 17601
rect 16117 17561 16129 17595
rect 16163 17592 16175 17595
rect 16592 17592 16620 17623
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17954 17660 17960 17672
rect 17543 17632 17960 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18598 17660 18604 17672
rect 18463 17632 18604 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 16163 17564 16620 17592
rect 19812 17592 19840 17623
rect 19978 17592 19984 17604
rect 19812 17564 19984 17592
rect 16163 17561 16175 17564
rect 16117 17555 16175 17561
rect 19978 17552 19984 17564
rect 20036 17552 20042 17604
rect 20530 17552 20536 17604
rect 20588 17592 20594 17604
rect 21269 17595 21327 17601
rect 21269 17592 21281 17595
rect 20588 17564 21281 17592
rect 20588 17552 20594 17564
rect 21269 17561 21281 17564
rect 21315 17561 21327 17595
rect 21269 17555 21327 17561
rect 14274 17484 14280 17536
rect 14332 17484 14338 17536
rect 14642 17484 14648 17536
rect 14700 17484 14706 17536
rect 14734 17484 14740 17536
rect 14792 17484 14798 17536
rect 20898 17484 20904 17536
rect 20956 17484 20962 17536
rect 21082 17533 21088 17536
rect 21069 17527 21088 17533
rect 21069 17493 21081 17527
rect 21140 17524 21146 17536
rect 21376 17524 21404 17700
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22922 17660 22928 17672
rect 22051 17632 22928 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 22281 17595 22339 17601
rect 22281 17561 22293 17595
rect 22327 17592 22339 17595
rect 22327 17564 22784 17592
rect 22327 17561 22339 17564
rect 22281 17555 22339 17561
rect 21140 17496 21404 17524
rect 21069 17487 21088 17493
rect 21082 17484 21088 17487
rect 21140 17484 21146 17496
rect 21450 17484 21456 17536
rect 21508 17524 21514 17536
rect 22756 17533 22784 17564
rect 22097 17527 22155 17533
rect 22097 17524 22109 17527
rect 21508 17496 22109 17524
rect 21508 17484 21514 17496
rect 22097 17493 22109 17496
rect 22143 17493 22155 17527
rect 22097 17487 22155 17493
rect 22741 17527 22799 17533
rect 22741 17493 22753 17527
rect 22787 17493 22799 17527
rect 22741 17487 22799 17493
rect 22909 17527 22967 17533
rect 22909 17493 22921 17527
rect 22955 17524 22967 17527
rect 23032 17524 23060 17700
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 23934 17620 23940 17672
rect 23992 17620 23998 17672
rect 24044 17669 24072 17700
rect 24029 17663 24087 17669
rect 24029 17629 24041 17663
rect 24075 17660 24087 17663
rect 24075 17632 24109 17660
rect 24075 17629 24087 17632
rect 24029 17623 24087 17629
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 27724 17669 27752 17700
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17629 27675 17663
rect 27617 17623 27675 17629
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17629 27767 17663
rect 27709 17623 27767 17629
rect 23109 17595 23167 17601
rect 23109 17561 23121 17595
rect 23155 17592 23167 17595
rect 23382 17592 23388 17604
rect 23155 17564 23388 17592
rect 23155 17561 23167 17564
rect 23109 17555 23167 17561
rect 23382 17552 23388 17564
rect 23440 17552 23446 17604
rect 24848 17595 24906 17601
rect 24848 17561 24860 17595
rect 24894 17592 24906 17595
rect 25038 17592 25044 17604
rect 24894 17564 25044 17592
rect 24894 17561 24906 17564
rect 24848 17555 24906 17561
rect 25038 17552 25044 17564
rect 25096 17552 25102 17604
rect 27632 17592 27660 17623
rect 27982 17620 27988 17672
rect 28040 17620 28046 17672
rect 28350 17620 28356 17672
rect 28408 17660 28414 17672
rect 30024 17669 30052 17768
rect 30650 17728 30656 17740
rect 30116 17700 30656 17728
rect 30116 17669 30144 17700
rect 30650 17688 30656 17700
rect 30708 17688 30714 17740
rect 30009 17663 30067 17669
rect 28408 17632 28948 17660
rect 28408 17620 28414 17632
rect 27632 17564 27752 17592
rect 22955 17496 23060 17524
rect 27724 17524 27752 17564
rect 27798 17552 27804 17604
rect 27856 17552 27862 17604
rect 28813 17595 28871 17601
rect 28813 17561 28825 17595
rect 28859 17561 28871 17595
rect 28920 17592 28948 17632
rect 30009 17629 30021 17663
rect 30055 17629 30067 17663
rect 30009 17623 30067 17629
rect 30101 17663 30159 17669
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 30374 17620 30380 17672
rect 30432 17620 30438 17672
rect 30852 17669 30880 17768
rect 31938 17756 31944 17768
rect 31996 17756 32002 17808
rect 32125 17799 32183 17805
rect 32125 17765 32137 17799
rect 32171 17796 32183 17799
rect 38197 17799 38255 17805
rect 32171 17768 38148 17796
rect 32171 17765 32183 17768
rect 32125 17759 32183 17765
rect 34514 17728 34520 17740
rect 31726 17700 34520 17728
rect 30837 17663 30895 17669
rect 30837 17629 30849 17663
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 31021 17663 31079 17669
rect 31021 17629 31033 17663
rect 31067 17660 31079 17663
rect 31726 17660 31754 17700
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 36262 17688 36268 17740
rect 36320 17688 36326 17740
rect 36357 17731 36415 17737
rect 36357 17697 36369 17731
rect 36403 17728 36415 17731
rect 36403 17700 37780 17728
rect 36403 17697 36415 17700
rect 36357 17691 36415 17697
rect 37752 17672 37780 17700
rect 37826 17688 37832 17740
rect 37884 17688 37890 17740
rect 31067 17632 31754 17660
rect 32769 17663 32827 17669
rect 31067 17629 31079 17632
rect 31021 17623 31079 17629
rect 32769 17629 32781 17663
rect 32815 17629 32827 17663
rect 32769 17623 32827 17629
rect 30193 17595 30251 17601
rect 30193 17592 30205 17595
rect 28920 17564 30205 17592
rect 28813 17555 28871 17561
rect 30193 17561 30205 17564
rect 30239 17592 30251 17595
rect 30929 17595 30987 17601
rect 30929 17592 30941 17595
rect 30239 17564 30941 17592
rect 30239 17561 30251 17564
rect 30193 17555 30251 17561
rect 30929 17561 30941 17564
rect 30975 17561 30987 17595
rect 32784 17592 32812 17623
rect 32858 17620 32864 17672
rect 32916 17660 32922 17672
rect 32953 17663 33011 17669
rect 32953 17660 32965 17663
rect 32916 17632 32965 17660
rect 32916 17620 32922 17632
rect 32953 17629 32965 17632
rect 32999 17629 33011 17663
rect 32953 17623 33011 17629
rect 33042 17620 33048 17672
rect 33100 17620 33106 17672
rect 34146 17620 34152 17672
rect 34204 17620 34210 17672
rect 34330 17620 34336 17672
rect 34388 17620 34394 17672
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 34480 17635 35080 17660
rect 34480 17632 35081 17635
rect 34480 17620 34486 17632
rect 35023 17629 35081 17632
rect 35023 17595 35035 17629
rect 35069 17595 35081 17629
rect 36630 17620 36636 17672
rect 36688 17620 36694 17672
rect 36725 17663 36783 17669
rect 36725 17629 36737 17663
rect 36771 17629 36783 17663
rect 36725 17623 36783 17629
rect 37001 17663 37059 17669
rect 37001 17629 37013 17663
rect 37047 17660 37059 17663
rect 37461 17663 37519 17669
rect 37461 17660 37473 17663
rect 37047 17632 37473 17660
rect 37047 17629 37059 17632
rect 37001 17623 37059 17629
rect 37461 17629 37473 17632
rect 37507 17629 37519 17663
rect 37461 17623 37519 17629
rect 32784 17564 34836 17592
rect 35023 17589 35081 17595
rect 35253 17595 35311 17601
rect 30929 17555 30987 17561
rect 27982 17524 27988 17536
rect 27724 17496 27988 17524
rect 22955 17493 22967 17496
rect 22909 17487 22967 17493
rect 27982 17484 27988 17496
rect 28040 17524 28046 17536
rect 28166 17524 28172 17536
rect 28040 17496 28172 17524
rect 28040 17484 28046 17496
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 28626 17533 28632 17536
rect 28613 17527 28632 17533
rect 28613 17493 28625 17527
rect 28613 17487 28632 17493
rect 28626 17484 28632 17487
rect 28684 17484 28690 17536
rect 28828 17524 28856 17555
rect 34808 17536 34836 17564
rect 35253 17561 35265 17595
rect 35299 17592 35311 17595
rect 35894 17592 35900 17604
rect 35299 17564 35900 17592
rect 35299 17561 35311 17564
rect 35253 17555 35311 17561
rect 35894 17552 35900 17564
rect 35952 17592 35958 17604
rect 36740 17592 36768 17623
rect 37642 17620 37648 17672
rect 37700 17620 37706 17672
rect 37734 17620 37740 17672
rect 37792 17620 37798 17672
rect 37918 17620 37924 17672
rect 37976 17660 37982 17672
rect 38013 17663 38071 17669
rect 38013 17660 38025 17663
rect 37976 17632 38025 17660
rect 37976 17620 37982 17632
rect 38013 17629 38025 17632
rect 38059 17629 38071 17663
rect 38120 17660 38148 17768
rect 38197 17765 38209 17799
rect 38243 17796 38255 17799
rect 39114 17796 39120 17808
rect 38243 17768 39120 17796
rect 38243 17765 38255 17768
rect 38197 17759 38255 17765
rect 39114 17756 39120 17768
rect 39172 17756 39178 17808
rect 41414 17688 41420 17740
rect 41472 17728 41478 17740
rect 41966 17728 41972 17740
rect 41472 17700 41972 17728
rect 41472 17688 41478 17700
rect 41966 17688 41972 17700
rect 42024 17688 42030 17740
rect 38120 17632 38792 17660
rect 38013 17623 38071 17629
rect 35952 17564 36768 17592
rect 38028 17592 38056 17623
rect 38470 17592 38476 17604
rect 38028 17564 38476 17592
rect 35952 17552 35958 17564
rect 38470 17552 38476 17564
rect 38528 17552 38534 17604
rect 38657 17595 38715 17601
rect 38657 17561 38669 17595
rect 38703 17561 38715 17595
rect 38764 17592 38792 17632
rect 38838 17620 38844 17672
rect 38896 17620 38902 17672
rect 38933 17663 38991 17669
rect 38933 17629 38945 17663
rect 38979 17660 38991 17663
rect 40218 17660 40224 17672
rect 38979 17632 40224 17660
rect 38979 17629 38991 17632
rect 38933 17623 38991 17629
rect 40218 17620 40224 17632
rect 40276 17620 40282 17672
rect 40310 17620 40316 17672
rect 40368 17620 40374 17672
rect 41138 17620 41144 17672
rect 41196 17620 41202 17672
rect 42242 17669 42248 17672
rect 42236 17660 42248 17669
rect 42203 17632 42248 17660
rect 42236 17623 42248 17632
rect 42242 17620 42248 17623
rect 42300 17620 42306 17672
rect 43530 17592 43536 17604
rect 38764 17564 43536 17592
rect 38657 17555 38715 17561
rect 28902 17524 28908 17536
rect 28828 17496 28908 17524
rect 28902 17484 28908 17496
rect 28960 17484 28966 17536
rect 32122 17484 32128 17536
rect 32180 17524 32186 17536
rect 32585 17527 32643 17533
rect 32585 17524 32597 17527
rect 32180 17496 32597 17524
rect 32180 17484 32186 17496
rect 32585 17493 32597 17496
rect 32631 17493 32643 17527
rect 32585 17487 32643 17493
rect 34790 17484 34796 17536
rect 34848 17524 34854 17536
rect 34885 17527 34943 17533
rect 34885 17524 34897 17527
rect 34848 17496 34897 17524
rect 34848 17484 34854 17496
rect 34885 17493 34897 17496
rect 34931 17493 34943 17527
rect 34885 17487 34943 17493
rect 36538 17484 36544 17536
rect 36596 17484 36602 17536
rect 37734 17484 37740 17536
rect 37792 17524 37798 17536
rect 37918 17524 37924 17536
rect 37792 17496 37924 17524
rect 37792 17484 37798 17496
rect 37918 17484 37924 17496
rect 37976 17484 37982 17536
rect 38672 17524 38700 17555
rect 43530 17552 43536 17564
rect 43588 17552 43594 17604
rect 38746 17524 38752 17536
rect 38672 17496 38752 17524
rect 38746 17484 38752 17496
rect 38804 17484 38810 17536
rect 39117 17527 39175 17533
rect 39117 17493 39129 17527
rect 39163 17524 39175 17527
rect 39482 17524 39488 17536
rect 39163 17496 39488 17524
rect 39163 17493 39175 17496
rect 39117 17487 39175 17493
rect 39482 17484 39488 17496
rect 39540 17484 39546 17536
rect 1104 17434 43884 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 43884 17434
rect 1104 17360 43884 17382
rect 14829 17323 14887 17329
rect 14829 17289 14841 17323
rect 14875 17320 14887 17323
rect 14918 17320 14924 17332
rect 14875 17292 14924 17320
rect 14875 17289 14887 17292
rect 14829 17283 14887 17289
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15657 17323 15715 17329
rect 15657 17320 15669 17323
rect 15620 17292 15669 17320
rect 15620 17280 15626 17292
rect 15657 17289 15669 17292
rect 15703 17289 15715 17323
rect 15657 17283 15715 17289
rect 18230 17280 18236 17332
rect 18288 17320 18294 17332
rect 18690 17320 18696 17332
rect 18288 17292 18696 17320
rect 18288 17280 18294 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 20530 17280 20536 17332
rect 20588 17280 20594 17332
rect 24026 17320 24032 17332
rect 20640 17292 24032 17320
rect 14274 17252 14280 17264
rect 12820 17224 14280 17252
rect 12820 17193 12848 17224
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 14642 17212 14648 17264
rect 14700 17252 14706 17264
rect 15473 17255 15531 17261
rect 15473 17252 15485 17255
rect 14700 17224 15485 17252
rect 14700 17212 14706 17224
rect 15473 17221 15485 17224
rect 15519 17221 15531 17255
rect 15473 17215 15531 17221
rect 16960 17224 19196 17252
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13705 17187 13763 17193
rect 13705 17184 13717 17187
rect 13596 17156 13717 17184
rect 13596 17144 13602 17156
rect 13705 17153 13717 17156
rect 13751 17153 13763 17187
rect 13705 17147 13763 17153
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 16960 17184 16988 17224
rect 19168 17196 19196 17224
rect 19242 17212 19248 17264
rect 19300 17252 19306 17264
rect 20640 17252 20668 17292
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 28350 17320 28356 17332
rect 25363 17292 28356 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 28350 17280 28356 17292
rect 28408 17280 28414 17332
rect 28534 17280 28540 17332
rect 28592 17280 28598 17332
rect 31846 17320 31852 17332
rect 31312 17292 31852 17320
rect 24578 17252 24584 17264
rect 19300 17224 20668 17252
rect 22020 17224 24584 17252
rect 19300 17212 19306 17224
rect 17126 17193 17132 17196
rect 17120 17184 17132 17193
rect 16908 17156 16988 17184
rect 17087 17156 17132 17184
rect 16908 17144 16914 17156
rect 17120 17147 17132 17156
rect 17126 17144 17132 17147
rect 17184 17144 17190 17196
rect 19150 17144 19156 17196
rect 19208 17144 19214 17196
rect 19420 17187 19478 17193
rect 19420 17153 19432 17187
rect 19466 17184 19478 17187
rect 20898 17184 20904 17196
rect 19466 17156 20904 17184
rect 19466 17153 19478 17156
rect 19420 17147 19478 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 22020 17193 22048 17224
rect 24578 17212 24584 17224
rect 24636 17252 24642 17264
rect 25130 17252 25136 17264
rect 24636 17224 25136 17252
rect 24636 17212 24642 17224
rect 25130 17212 25136 17224
rect 25188 17212 25194 17264
rect 29086 17252 29092 17264
rect 25700 17224 29092 17252
rect 25700 17196 25728 17224
rect 29086 17212 29092 17224
rect 29144 17212 29150 17264
rect 30742 17212 30748 17264
rect 30800 17212 30806 17264
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22261 17187 22319 17193
rect 22261 17184 22273 17187
rect 22005 17147 22063 17153
rect 22112 17156 22273 17184
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13412 17088 13461 17116
rect 13412 17076 13418 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 12986 16940 12992 16992
rect 13044 16940 13050 16992
rect 21284 16980 21312 17147
rect 22112 17116 22140 17156
rect 22261 17153 22273 17156
rect 22307 17153 22319 17187
rect 22261 17147 22319 17153
rect 25314 17187 25372 17193
rect 25314 17153 25326 17187
rect 25360 17184 25372 17187
rect 25682 17184 25688 17196
rect 25360 17156 25688 17184
rect 25360 17153 25372 17156
rect 25314 17147 25372 17153
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 25774 17144 25780 17196
rect 25832 17144 25838 17196
rect 27430 17193 27436 17196
rect 27424 17147 27436 17193
rect 27430 17144 27436 17147
rect 27488 17144 27494 17196
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29730 17184 29736 17196
rect 29052 17156 29736 17184
rect 29052 17144 29058 17156
rect 29730 17144 29736 17156
rect 29788 17144 29794 17196
rect 31312 17193 31340 17292
rect 31846 17280 31852 17292
rect 31904 17280 31910 17332
rect 32858 17280 32864 17332
rect 32916 17320 32922 17332
rect 33689 17323 33747 17329
rect 33689 17320 33701 17323
rect 32916 17292 33701 17320
rect 32916 17280 32922 17292
rect 33689 17289 33701 17292
rect 33735 17289 33747 17323
rect 33689 17283 33747 17289
rect 34609 17323 34667 17329
rect 34609 17289 34621 17323
rect 34655 17320 34667 17323
rect 36170 17320 36176 17332
rect 34655 17292 36176 17320
rect 34655 17289 34667 17292
rect 34609 17283 34667 17289
rect 36170 17280 36176 17292
rect 36228 17280 36234 17332
rect 36817 17323 36875 17329
rect 36817 17289 36829 17323
rect 36863 17320 36875 17323
rect 37642 17320 37648 17332
rect 36863 17292 37648 17320
rect 36863 17289 36875 17292
rect 36817 17283 36875 17289
rect 37642 17280 37648 17292
rect 37700 17280 37706 17332
rect 39117 17323 39175 17329
rect 39117 17289 39129 17323
rect 39163 17320 39175 17323
rect 39390 17320 39396 17332
rect 39163 17292 39396 17320
rect 39163 17289 39175 17292
rect 39117 17283 39175 17289
rect 39390 17280 39396 17292
rect 39448 17280 39454 17332
rect 41046 17280 41052 17332
rect 41104 17320 41110 17332
rect 41141 17323 41199 17329
rect 41141 17320 41153 17323
rect 41104 17292 41153 17320
rect 41104 17280 41110 17292
rect 41141 17289 41153 17292
rect 41187 17320 41199 17323
rect 41874 17320 41880 17332
rect 41187 17292 41880 17320
rect 41187 17289 41199 17292
rect 41141 17283 41199 17289
rect 41874 17280 41880 17292
rect 41932 17280 41938 17332
rect 43070 17280 43076 17332
rect 43128 17320 43134 17332
rect 43165 17323 43223 17329
rect 43165 17320 43177 17323
rect 43128 17292 43177 17320
rect 43128 17280 43134 17292
rect 43165 17289 43177 17292
rect 43211 17289 43223 17323
rect 43165 17283 43223 17289
rect 31757 17255 31815 17261
rect 31757 17221 31769 17255
rect 31803 17252 31815 17255
rect 32554 17255 32612 17261
rect 32554 17252 32566 17255
rect 31803 17224 32566 17252
rect 31803 17221 31815 17224
rect 31757 17215 31815 17221
rect 32554 17221 32566 17224
rect 32600 17221 32612 17255
rect 32554 17215 32612 17221
rect 34514 17212 34520 17264
rect 34572 17252 34578 17264
rect 35345 17255 35403 17261
rect 34572 17224 34744 17252
rect 34572 17212 34578 17224
rect 31297 17187 31355 17193
rect 31297 17153 31309 17187
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31386 17144 31392 17196
rect 31444 17144 31450 17196
rect 31573 17187 31631 17193
rect 31573 17153 31585 17187
rect 31619 17184 31631 17187
rect 32122 17184 32128 17196
rect 31619 17156 32128 17184
rect 31619 17153 31631 17156
rect 31573 17147 31631 17153
rect 32122 17144 32128 17156
rect 32180 17144 32186 17196
rect 34422 17144 34428 17196
rect 34480 17144 34486 17196
rect 34606 17144 34612 17196
rect 34664 17144 34670 17196
rect 34716 17184 34744 17224
rect 35345 17221 35357 17255
rect 35391 17252 35403 17255
rect 35986 17252 35992 17264
rect 35391 17224 35992 17252
rect 35391 17221 35403 17224
rect 35345 17215 35403 17221
rect 35986 17212 35992 17224
rect 36044 17212 36050 17264
rect 37090 17212 37096 17264
rect 37148 17252 37154 17264
rect 38657 17255 38715 17261
rect 37148 17224 37780 17252
rect 37148 17212 37154 17224
rect 35529 17187 35587 17193
rect 35529 17184 35541 17187
rect 34716 17156 35541 17184
rect 35529 17153 35541 17156
rect 35575 17184 35587 17187
rect 36449 17187 36507 17193
rect 36449 17184 36461 17187
rect 35575 17156 36461 17184
rect 35575 17153 35587 17156
rect 35529 17147 35587 17153
rect 36449 17153 36461 17156
rect 36495 17153 36507 17187
rect 36449 17147 36507 17153
rect 36633 17187 36691 17193
rect 36633 17153 36645 17187
rect 36679 17184 36691 17187
rect 36722 17184 36728 17196
rect 36679 17156 36728 17184
rect 36679 17153 36691 17156
rect 36633 17147 36691 17153
rect 36722 17144 36728 17156
rect 36780 17144 36786 17196
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37752 17193 37780 17224
rect 38657 17221 38669 17255
rect 38703 17252 38715 17255
rect 38746 17252 38752 17264
rect 38703 17224 38752 17252
rect 38703 17221 38715 17224
rect 38657 17215 38715 17221
rect 38746 17212 38752 17224
rect 38804 17212 38810 17264
rect 41506 17212 41512 17264
rect 41564 17252 41570 17264
rect 41601 17255 41659 17261
rect 41601 17252 41613 17255
rect 41564 17224 41613 17252
rect 41564 17212 41570 17224
rect 41601 17221 41613 17224
rect 41647 17221 41659 17255
rect 41601 17215 41659 17221
rect 41690 17212 41696 17264
rect 41748 17252 41754 17264
rect 43257 17255 43315 17261
rect 43257 17252 43269 17255
rect 41748 17224 43269 17252
rect 41748 17212 41754 17224
rect 43257 17221 43269 17224
rect 43303 17221 43315 17255
rect 43257 17215 43315 17221
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37424 17156 37657 17184
rect 37424 17144 37430 17156
rect 37645 17153 37657 17156
rect 37691 17153 37703 17187
rect 37645 17147 37703 17153
rect 37737 17187 37795 17193
rect 37737 17153 37749 17187
rect 37783 17153 37795 17187
rect 37737 17147 37795 17153
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 38378 17184 38384 17196
rect 37967 17156 38384 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38378 17144 38384 17156
rect 38436 17144 38442 17196
rect 38930 17144 38936 17196
rect 38988 17144 38994 17196
rect 39945 17187 40003 17193
rect 39945 17153 39957 17187
rect 39991 17184 40003 17187
rect 40034 17184 40040 17196
rect 39991 17156 40040 17184
rect 39991 17153 40003 17156
rect 39945 17147 40003 17153
rect 40034 17144 40040 17156
rect 40092 17144 40098 17196
rect 40126 17144 40132 17196
rect 40184 17193 40190 17196
rect 40184 17187 40199 17193
rect 40187 17184 40199 17187
rect 41969 17187 42027 17193
rect 40187 17156 40448 17184
rect 40187 17153 40199 17156
rect 40184 17147 40199 17153
rect 40184 17144 40190 17147
rect 21468 17088 22140 17116
rect 21468 17057 21496 17088
rect 27154 17076 27160 17128
rect 27212 17076 27218 17128
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 29273 17119 29331 17125
rect 29273 17116 29285 17119
rect 28776 17088 29285 17116
rect 28776 17076 28782 17088
rect 29273 17085 29285 17088
rect 29319 17085 29331 17119
rect 29273 17079 29331 17085
rect 21453 17051 21511 17057
rect 21453 17017 21465 17051
rect 21499 17017 21511 17051
rect 21453 17011 21511 17017
rect 25038 17008 25044 17060
rect 25096 17048 25102 17060
rect 25133 17051 25191 17057
rect 25133 17048 25145 17051
rect 25096 17020 25145 17048
rect 25096 17008 25102 17020
rect 25133 17017 25145 17020
rect 25179 17017 25191 17051
rect 25133 17011 25191 17017
rect 29089 17051 29147 17057
rect 29089 17017 29101 17051
rect 29135 17017 29147 17051
rect 29288 17048 29316 17079
rect 29546 17076 29552 17128
rect 29604 17116 29610 17128
rect 29917 17119 29975 17125
rect 29917 17116 29929 17119
rect 29604 17088 29929 17116
rect 29604 17076 29610 17088
rect 29917 17085 29929 17088
rect 29963 17116 29975 17119
rect 32309 17119 32367 17125
rect 32309 17116 32321 17119
rect 29963 17088 32321 17116
rect 29963 17085 29975 17088
rect 29917 17079 29975 17085
rect 32309 17085 32321 17088
rect 32355 17085 32367 17119
rect 32309 17079 32367 17085
rect 34330 17076 34336 17128
rect 34388 17116 34394 17128
rect 36357 17119 36415 17125
rect 36357 17116 36369 17119
rect 34388 17088 36369 17116
rect 34388 17076 34394 17088
rect 36357 17085 36369 17088
rect 36403 17116 36415 17119
rect 36906 17116 36912 17128
rect 36403 17088 36912 17116
rect 36403 17085 36415 17088
rect 36357 17079 36415 17085
rect 36906 17076 36912 17088
rect 36964 17116 36970 17128
rect 36964 17088 37688 17116
rect 36964 17076 36970 17088
rect 31938 17048 31944 17060
rect 29288 17020 31944 17048
rect 29089 17011 29147 17017
rect 22186 16980 22192 16992
rect 21284 16952 22192 16980
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 23382 16940 23388 16992
rect 23440 16940 23446 16992
rect 25685 16983 25743 16989
rect 25685 16949 25697 16983
rect 25731 16980 25743 16983
rect 26510 16980 26516 16992
rect 25731 16952 26516 16980
rect 25731 16949 25743 16952
rect 25685 16943 25743 16949
rect 26510 16940 26516 16952
rect 26568 16940 26574 16992
rect 28626 16940 28632 16992
rect 28684 16980 28690 16992
rect 28997 16983 29055 16989
rect 28997 16980 29009 16983
rect 28684 16952 29009 16980
rect 28684 16940 28690 16952
rect 28997 16949 29009 16952
rect 29043 16949 29055 16983
rect 29104 16980 29132 17011
rect 31938 17008 31944 17020
rect 31996 17008 32002 17060
rect 37458 17008 37464 17060
rect 37516 17008 37522 17060
rect 29178 16980 29184 16992
rect 29104 16952 29184 16980
rect 28997 16943 29055 16949
rect 29178 16940 29184 16952
rect 29236 16980 29242 16992
rect 31018 16980 31024 16992
rect 29236 16952 31024 16980
rect 29236 16940 29242 16952
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 34606 16940 34612 16992
rect 34664 16980 34670 16992
rect 35161 16983 35219 16989
rect 35161 16980 35173 16983
rect 34664 16952 35173 16980
rect 34664 16940 34670 16952
rect 35161 16949 35173 16952
rect 35207 16980 35219 16983
rect 37550 16980 37556 16992
rect 35207 16952 37556 16980
rect 35207 16949 35219 16952
rect 35161 16943 35219 16949
rect 37550 16940 37556 16952
rect 37608 16940 37614 16992
rect 37660 16980 37688 17088
rect 38838 17076 38844 17128
rect 38896 17116 38902 17128
rect 39114 17116 39120 17128
rect 38896 17088 39120 17116
rect 38896 17076 38902 17088
rect 39114 17076 39120 17088
rect 39172 17076 39178 17128
rect 40420 17116 40448 17156
rect 41969 17153 41981 17187
rect 42015 17184 42027 17187
rect 42242 17184 42248 17196
rect 42015 17156 42248 17184
rect 42015 17153 42027 17156
rect 41969 17147 42027 17153
rect 42242 17144 42248 17156
rect 42300 17184 42306 17196
rect 43990 17184 43996 17196
rect 42300 17156 43996 17184
rect 42300 17144 42306 17156
rect 43990 17144 43996 17156
rect 44048 17144 44054 17196
rect 43165 17119 43223 17125
rect 40420 17088 42748 17116
rect 39942 17008 39948 17060
rect 40000 17008 40006 17060
rect 42720 17057 42748 17088
rect 43165 17085 43177 17119
rect 43211 17116 43223 17119
rect 43530 17116 43536 17128
rect 43211 17088 43536 17116
rect 43211 17085 43223 17088
rect 43165 17079 43223 17085
rect 43530 17076 43536 17088
rect 43588 17076 43594 17128
rect 42705 17051 42763 17057
rect 42705 17017 42717 17051
rect 42751 17017 42763 17051
rect 42705 17011 42763 17017
rect 37829 16983 37887 16989
rect 37829 16980 37841 16983
rect 37660 16952 37841 16980
rect 37829 16949 37841 16952
rect 37875 16980 37887 16983
rect 38286 16980 38292 16992
rect 37875 16952 38292 16980
rect 37875 16949 37887 16952
rect 37829 16943 37887 16949
rect 38286 16940 38292 16952
rect 38344 16940 38350 16992
rect 38470 16940 38476 16992
rect 38528 16980 38534 16992
rect 38657 16983 38715 16989
rect 38657 16980 38669 16983
rect 38528 16952 38669 16980
rect 38528 16940 38534 16952
rect 38657 16949 38669 16952
rect 38703 16949 38715 16983
rect 38657 16943 38715 16949
rect 1104 16890 43884 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 43884 16890
rect 1104 16816 43884 16838
rect 13538 16736 13544 16788
rect 13596 16736 13602 16788
rect 19812 16748 20760 16776
rect 14734 16708 14740 16720
rect 14660 16680 14740 16708
rect 14660 16640 14688 16680
rect 14734 16668 14740 16680
rect 14792 16708 14798 16720
rect 17954 16708 17960 16720
rect 14792 16680 17960 16708
rect 14792 16668 14798 16680
rect 14568 16612 14688 16640
rect 14829 16643 14887 16649
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 13771 16544 14320 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14292 16445 14320 16544
rect 14568 16504 14596 16612
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 15194 16640 15200 16652
rect 14875 16612 15200 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 15194 16600 15200 16612
rect 15252 16640 15258 16652
rect 15470 16640 15476 16652
rect 15252 16612 15476 16640
rect 15252 16600 15258 16612
rect 15470 16600 15476 16612
rect 15528 16640 15534 16652
rect 17604 16649 17632 16680
rect 17954 16668 17960 16680
rect 18012 16708 18018 16720
rect 19242 16708 19248 16720
rect 18012 16680 19248 16708
rect 18012 16668 18018 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15528 16612 16313 16640
rect 15528 16600 15534 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 17678 16600 17684 16652
rect 17736 16600 17742 16652
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19812 16649 19840 16748
rect 20162 16708 20168 16720
rect 19996 16680 20168 16708
rect 19996 16649 20024 16680
rect 20162 16668 20168 16680
rect 20220 16668 20226 16720
rect 20441 16711 20499 16717
rect 20441 16677 20453 16711
rect 20487 16708 20499 16711
rect 20487 16680 20668 16708
rect 20487 16677 20499 16680
rect 20441 16671 20499 16677
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19116 16612 19809 16640
rect 19116 16600 19122 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19981 16643 20039 16649
rect 19981 16609 19993 16643
rect 20027 16609 20039 16643
rect 20530 16640 20536 16652
rect 19981 16603 20039 16609
rect 20088 16612 20536 16640
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 14918 16572 14924 16584
rect 14691 16544 14924 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15620 16544 15853 16572
rect 15620 16532 15626 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 18230 16572 18236 16584
rect 17543 16544 18236 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16572 18383 16575
rect 18598 16572 18604 16584
rect 18371 16544 18604 16572
rect 18371 16541 18383 16544
rect 18325 16535 18383 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 20088 16581 20116 16612
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16541 20131 16575
rect 20640 16572 20668 16680
rect 20732 16640 20760 16748
rect 20898 16736 20904 16788
rect 20956 16736 20962 16788
rect 22186 16736 22192 16788
rect 22244 16736 22250 16788
rect 24578 16736 24584 16788
rect 24636 16776 24642 16788
rect 24636 16748 26464 16776
rect 24636 16736 24642 16748
rect 21634 16668 21640 16720
rect 21692 16668 21698 16720
rect 26436 16649 26464 16748
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 27525 16779 27583 16785
rect 27525 16776 27537 16779
rect 27488 16748 27537 16776
rect 27488 16736 27494 16748
rect 27525 16745 27537 16748
rect 27571 16745 27583 16779
rect 27525 16739 27583 16745
rect 27798 16736 27804 16788
rect 27856 16776 27862 16788
rect 28537 16779 28595 16785
rect 28537 16776 28549 16779
rect 27856 16748 28549 16776
rect 27856 16736 27862 16748
rect 28537 16745 28549 16748
rect 28583 16745 28595 16779
rect 28994 16776 29000 16788
rect 28537 16739 28595 16745
rect 28644 16748 29000 16776
rect 28644 16708 28672 16748
rect 28994 16736 29000 16748
rect 29052 16736 29058 16788
rect 30190 16736 30196 16788
rect 30248 16736 30254 16788
rect 30374 16736 30380 16788
rect 30432 16776 30438 16788
rect 31573 16779 31631 16785
rect 31573 16776 31585 16779
rect 30432 16748 31585 16776
rect 30432 16736 30438 16748
rect 31573 16745 31585 16748
rect 31619 16745 31631 16779
rect 31573 16739 31631 16745
rect 31757 16779 31815 16785
rect 31757 16745 31769 16779
rect 31803 16745 31815 16779
rect 31757 16739 31815 16745
rect 30650 16708 30656 16720
rect 27724 16680 28672 16708
rect 28736 16680 30656 16708
rect 22741 16643 22799 16649
rect 22741 16640 22753 16643
rect 20732 16612 22753 16640
rect 22741 16609 22753 16612
rect 22787 16609 22799 16643
rect 22741 16603 22799 16609
rect 26421 16643 26479 16649
rect 26421 16609 26433 16643
rect 26467 16609 26479 16643
rect 26421 16603 26479 16609
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20640 16544 21097 16572
rect 20073 16535 20131 16541
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16572 22615 16575
rect 23382 16572 23388 16584
rect 22603 16544 23388 16572
rect 22603 16541 22615 16544
rect 22557 16535 22615 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 25130 16532 25136 16584
rect 25188 16572 25194 16584
rect 25961 16575 26019 16581
rect 25961 16572 25973 16575
rect 25188 16544 25973 16572
rect 25188 16532 25194 16544
rect 25961 16541 25973 16544
rect 26007 16541 26019 16575
rect 25961 16535 26019 16541
rect 26510 16532 26516 16584
rect 26568 16532 26574 16584
rect 26697 16575 26755 16581
rect 26697 16541 26709 16575
rect 26743 16572 26755 16575
rect 27614 16572 27620 16584
rect 26743 16544 27620 16572
rect 26743 16541 26755 16544
rect 26697 16535 26755 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 27724 16581 27752 16680
rect 28534 16640 28540 16652
rect 27816 16612 28540 16640
rect 27816 16581 27844 16612
rect 28534 16600 28540 16612
rect 28592 16600 28598 16652
rect 28736 16649 28764 16680
rect 30650 16668 30656 16680
rect 30708 16668 30714 16720
rect 31772 16708 31800 16739
rect 32398 16736 32404 16788
rect 32456 16736 32462 16788
rect 32585 16779 32643 16785
rect 32585 16745 32597 16779
rect 32631 16776 32643 16779
rect 33410 16776 33416 16788
rect 32631 16748 33416 16776
rect 32631 16745 32643 16748
rect 32585 16739 32643 16745
rect 33410 16736 33416 16748
rect 33468 16736 33474 16788
rect 35066 16776 35072 16788
rect 34072 16748 35072 16776
rect 33505 16711 33563 16717
rect 31772 16680 33456 16708
rect 28721 16643 28779 16649
rect 28721 16609 28733 16643
rect 28767 16609 28779 16643
rect 28721 16603 28779 16609
rect 28997 16643 29055 16649
rect 28997 16609 29009 16643
rect 29043 16640 29055 16643
rect 29086 16640 29092 16652
rect 29043 16612 29092 16640
rect 29043 16609 29055 16612
rect 28997 16603 29055 16609
rect 29086 16600 29092 16612
rect 29144 16600 29150 16652
rect 30745 16643 30803 16649
rect 30745 16640 30757 16643
rect 30392 16612 30757 16640
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 28077 16575 28135 16581
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28626 16572 28632 16584
rect 28123 16544 28632 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 28626 16532 28632 16544
rect 28684 16532 28690 16584
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 14737 16507 14795 16513
rect 14737 16504 14749 16507
rect 14568 16476 14749 16504
rect 14737 16473 14749 16476
rect 14783 16473 14795 16507
rect 14737 16467 14795 16473
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17000 16476 22094 16504
rect 17000 16464 17006 16476
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16405 14335 16439
rect 14277 16399 14335 16405
rect 15654 16396 15660 16448
rect 15712 16396 15718 16448
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 17092 16408 17141 16436
rect 17092 16396 17098 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 22066 16436 22094 16476
rect 22370 16464 22376 16516
rect 22428 16504 22434 16516
rect 22649 16507 22707 16513
rect 22649 16504 22661 16507
rect 22428 16476 22661 16504
rect 22428 16464 22434 16476
rect 22649 16473 22661 16476
rect 22695 16473 22707 16507
rect 22649 16467 22707 16473
rect 25716 16507 25774 16513
rect 25716 16473 25728 16507
rect 25762 16504 25774 16507
rect 26881 16507 26939 16513
rect 26881 16504 26893 16507
rect 25762 16476 26893 16504
rect 25762 16473 25774 16476
rect 25716 16467 25774 16473
rect 26881 16473 26893 16476
rect 26927 16473 26939 16507
rect 26881 16467 26939 16473
rect 27893 16507 27951 16513
rect 27893 16473 27905 16507
rect 27939 16473 27951 16507
rect 28828 16504 28856 16535
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 30392 16572 30420 16612
rect 30745 16609 30757 16612
rect 30791 16640 30803 16643
rect 32490 16640 32496 16652
rect 30791 16612 32496 16640
rect 30791 16609 30803 16612
rect 30745 16603 30803 16609
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 33428 16640 33456 16680
rect 33505 16677 33517 16711
rect 33551 16708 33563 16711
rect 34072 16708 34100 16748
rect 35066 16736 35072 16748
rect 35124 16736 35130 16788
rect 35161 16779 35219 16785
rect 35161 16745 35173 16779
rect 35207 16776 35219 16779
rect 35526 16776 35532 16788
rect 35207 16748 35532 16776
rect 35207 16745 35219 16748
rect 35161 16739 35219 16745
rect 35176 16708 35204 16739
rect 35526 16736 35532 16748
rect 35584 16736 35590 16788
rect 36262 16736 36268 16788
rect 36320 16736 36326 16788
rect 37461 16779 37519 16785
rect 37461 16745 37473 16779
rect 37507 16776 37519 16779
rect 37734 16776 37740 16788
rect 37507 16748 37740 16776
rect 37507 16745 37519 16748
rect 37461 16739 37519 16745
rect 37734 16736 37740 16748
rect 37792 16736 37798 16788
rect 37826 16736 37832 16788
rect 37884 16776 37890 16788
rect 37921 16779 37979 16785
rect 37921 16776 37933 16779
rect 37884 16748 37933 16776
rect 37884 16736 37890 16748
rect 37921 16745 37933 16748
rect 37967 16745 37979 16779
rect 37921 16739 37979 16745
rect 38378 16736 38384 16788
rect 38436 16776 38442 16788
rect 39025 16779 39083 16785
rect 39025 16776 39037 16779
rect 38436 16748 39037 16776
rect 38436 16736 38442 16748
rect 39025 16745 39037 16748
rect 39071 16745 39083 16779
rect 39025 16739 39083 16745
rect 39850 16736 39856 16788
rect 39908 16776 39914 16788
rect 40129 16779 40187 16785
rect 40129 16776 40141 16779
rect 39908 16748 40141 16776
rect 39908 16736 39914 16748
rect 40129 16745 40141 16748
rect 40175 16745 40187 16779
rect 40129 16739 40187 16745
rect 33551 16680 34100 16708
rect 34164 16680 35204 16708
rect 33551 16677 33563 16680
rect 33505 16671 33563 16677
rect 34164 16640 34192 16680
rect 37182 16668 37188 16720
rect 37240 16708 37246 16720
rect 37240 16680 39988 16708
rect 37240 16668 37246 16680
rect 33428 16612 34192 16640
rect 34974 16600 34980 16652
rect 35032 16600 35038 16652
rect 36173 16643 36231 16649
rect 36173 16640 36185 16643
rect 35084 16612 36185 16640
rect 28960 16544 30420 16572
rect 30469 16575 30527 16581
rect 28960 16532 28966 16544
rect 30469 16541 30481 16575
rect 30515 16572 30527 16575
rect 32306 16572 32312 16584
rect 30515 16544 32312 16572
rect 30515 16541 30527 16544
rect 30469 16535 30527 16541
rect 32306 16532 32312 16544
rect 32364 16532 32370 16584
rect 34057 16575 34115 16581
rect 34057 16541 34069 16575
rect 34103 16541 34115 16575
rect 34057 16535 34115 16541
rect 34241 16575 34299 16581
rect 34241 16541 34253 16575
rect 34287 16572 34299 16575
rect 34330 16572 34336 16584
rect 34287 16544 34336 16572
rect 34287 16541 34299 16544
rect 34241 16535 34299 16541
rect 29178 16504 29184 16516
rect 28828 16476 29184 16504
rect 27893 16467 27951 16473
rect 26970 16436 26976 16448
rect 22066 16408 26976 16436
rect 26970 16396 26976 16408
rect 27028 16396 27034 16448
rect 27908 16436 27936 16467
rect 29178 16464 29184 16476
rect 29236 16464 29242 16516
rect 30377 16507 30435 16513
rect 30377 16473 30389 16507
rect 30423 16504 30435 16507
rect 30650 16504 30656 16516
rect 30423 16476 30656 16504
rect 30423 16473 30435 16476
rect 30377 16467 30435 16473
rect 30650 16464 30656 16476
rect 30708 16464 30714 16516
rect 31294 16464 31300 16516
rect 31352 16504 31358 16516
rect 31725 16507 31783 16513
rect 31725 16504 31737 16507
rect 31352 16476 31737 16504
rect 31352 16464 31358 16476
rect 31725 16473 31737 16476
rect 31771 16504 31783 16507
rect 31771 16476 31892 16504
rect 31771 16473 31783 16476
rect 31725 16467 31783 16473
rect 28810 16436 28816 16448
rect 27908 16408 28816 16436
rect 28810 16396 28816 16408
rect 28868 16396 28874 16448
rect 30006 16396 30012 16448
rect 30064 16436 30070 16448
rect 30561 16439 30619 16445
rect 30561 16436 30573 16439
rect 30064 16408 30573 16436
rect 30064 16396 30070 16408
rect 30561 16405 30573 16408
rect 30607 16436 30619 16439
rect 31478 16436 31484 16448
rect 30607 16408 31484 16436
rect 30607 16405 30619 16408
rect 30561 16399 30619 16405
rect 31478 16396 31484 16408
rect 31536 16396 31542 16448
rect 31864 16436 31892 16476
rect 31938 16464 31944 16516
rect 31996 16464 32002 16516
rect 32769 16507 32827 16513
rect 32769 16473 32781 16507
rect 32815 16504 32827 16507
rect 32858 16504 32864 16516
rect 32815 16476 32864 16504
rect 32815 16473 32827 16476
rect 32769 16467 32827 16473
rect 32858 16464 32864 16476
rect 32916 16464 32922 16516
rect 33778 16464 33784 16516
rect 33836 16504 33842 16516
rect 34072 16504 34100 16535
rect 34330 16532 34336 16544
rect 34388 16572 34394 16584
rect 35084 16572 35112 16612
rect 36173 16609 36185 16612
rect 36219 16640 36231 16643
rect 37366 16640 37372 16652
rect 36219 16612 37372 16640
rect 36219 16609 36231 16612
rect 36173 16603 36231 16609
rect 37366 16600 37372 16612
rect 37424 16640 37430 16652
rect 38470 16640 38476 16652
rect 37424 16612 38476 16640
rect 37424 16600 37430 16612
rect 38470 16600 38476 16612
rect 38528 16640 38534 16652
rect 39117 16643 39175 16649
rect 39117 16640 39129 16643
rect 38528 16612 39129 16640
rect 38528 16600 38534 16612
rect 39117 16609 39129 16612
rect 39163 16609 39175 16643
rect 39117 16603 39175 16609
rect 34388 16544 35112 16572
rect 34388 16532 34394 16544
rect 35158 16532 35164 16584
rect 35216 16532 35222 16584
rect 35250 16532 35256 16584
rect 35308 16572 35314 16584
rect 35989 16575 36047 16581
rect 35989 16572 36001 16575
rect 35308 16544 36001 16572
rect 35308 16532 35314 16544
rect 35989 16541 36001 16544
rect 36035 16541 36047 16575
rect 35989 16535 36047 16541
rect 36096 16544 36400 16572
rect 33836 16476 34100 16504
rect 33836 16464 33842 16476
rect 34882 16464 34888 16516
rect 34940 16504 34946 16516
rect 36096 16504 36124 16544
rect 34940 16476 36124 16504
rect 36265 16507 36323 16513
rect 34940 16464 34946 16476
rect 36265 16473 36277 16507
rect 36311 16473 36323 16507
rect 36372 16504 36400 16544
rect 37182 16532 37188 16584
rect 37240 16532 37246 16584
rect 37274 16532 37280 16584
rect 37332 16532 37338 16584
rect 38102 16532 38108 16584
rect 38160 16532 38166 16584
rect 38381 16575 38439 16581
rect 38381 16541 38393 16575
rect 38427 16572 38439 16575
rect 38746 16572 38752 16584
rect 38427 16544 38752 16572
rect 38427 16541 38439 16544
rect 38381 16535 38439 16541
rect 38746 16532 38752 16544
rect 38804 16532 38810 16584
rect 39206 16532 39212 16584
rect 39264 16532 39270 16584
rect 39960 16572 39988 16680
rect 41524 16680 42564 16708
rect 41524 16649 41552 16680
rect 41509 16643 41567 16649
rect 41509 16609 41521 16643
rect 41555 16609 41567 16643
rect 41509 16603 41567 16609
rect 41690 16600 41696 16652
rect 41748 16600 41754 16652
rect 42536 16649 42564 16680
rect 42429 16643 42487 16649
rect 42429 16609 42441 16643
rect 42475 16609 42487 16643
rect 42429 16603 42487 16609
rect 42521 16643 42579 16649
rect 42521 16609 42533 16643
rect 42567 16640 42579 16643
rect 42886 16640 42892 16652
rect 42567 16612 42892 16640
rect 42567 16609 42579 16612
rect 42521 16603 42579 16609
rect 40218 16572 40224 16584
rect 39960 16544 40224 16572
rect 40218 16532 40224 16544
rect 40276 16532 40282 16584
rect 40310 16532 40316 16584
rect 40368 16572 40374 16584
rect 40405 16575 40463 16581
rect 40405 16572 40417 16575
rect 40368 16544 40417 16572
rect 40368 16532 40374 16544
rect 40405 16541 40417 16544
rect 40451 16541 40463 16575
rect 42444 16572 42472 16603
rect 42886 16600 42892 16612
rect 42944 16600 42950 16652
rect 42978 16572 42984 16584
rect 42444 16544 42984 16572
rect 40405 16535 40463 16541
rect 42978 16532 42984 16544
rect 43036 16532 43042 16584
rect 36446 16504 36452 16516
rect 36372 16476 36452 16504
rect 36265 16467 36323 16473
rect 32559 16439 32617 16445
rect 32559 16436 32571 16439
rect 31864 16408 32571 16436
rect 32559 16405 32571 16408
rect 32605 16436 32617 16439
rect 34057 16439 34115 16445
rect 34057 16436 34069 16439
rect 32605 16408 34069 16436
rect 32605 16405 32617 16408
rect 32559 16399 32617 16405
rect 34057 16405 34069 16408
rect 34103 16436 34115 16439
rect 34422 16436 34428 16448
rect 34103 16408 34428 16436
rect 34103 16405 34115 16408
rect 34057 16399 34115 16405
rect 34422 16396 34428 16408
rect 34480 16396 34486 16448
rect 35342 16396 35348 16448
rect 35400 16396 35406 16448
rect 35618 16396 35624 16448
rect 35676 16436 35682 16448
rect 35805 16439 35863 16445
rect 35805 16436 35817 16439
rect 35676 16408 35817 16436
rect 35676 16396 35682 16408
rect 35805 16405 35817 16408
rect 35851 16405 35863 16439
rect 35805 16399 35863 16405
rect 35986 16396 35992 16448
rect 36044 16436 36050 16448
rect 36280 16436 36308 16467
rect 36446 16464 36452 16476
rect 36504 16504 36510 16516
rect 37461 16507 37519 16513
rect 37461 16504 37473 16507
rect 36504 16476 37473 16504
rect 36504 16464 36510 16476
rect 37461 16473 37473 16476
rect 37507 16504 37519 16507
rect 37642 16504 37648 16516
rect 37507 16476 37648 16504
rect 37507 16473 37519 16476
rect 37461 16467 37519 16473
rect 37642 16464 37648 16476
rect 37700 16464 37706 16516
rect 38010 16464 38016 16516
rect 38068 16504 38074 16516
rect 41417 16507 41475 16513
rect 38068 16476 38884 16504
rect 38068 16464 38074 16476
rect 36044 16408 36308 16436
rect 36044 16396 36050 16408
rect 36814 16396 36820 16448
rect 36872 16436 36878 16448
rect 37001 16439 37059 16445
rect 37001 16436 37013 16439
rect 36872 16408 37013 16436
rect 36872 16396 36878 16408
rect 37001 16405 37013 16408
rect 37047 16405 37059 16439
rect 37001 16399 37059 16405
rect 37918 16396 37924 16448
rect 37976 16436 37982 16448
rect 38856 16445 38884 16476
rect 41417 16473 41429 16507
rect 41463 16504 41475 16507
rect 41506 16504 41512 16516
rect 41463 16476 41512 16504
rect 41463 16473 41475 16476
rect 41417 16467 41475 16473
rect 41506 16464 41512 16476
rect 41564 16504 41570 16516
rect 42613 16507 42671 16513
rect 42613 16504 42625 16507
rect 41564 16476 42625 16504
rect 41564 16464 41570 16476
rect 42613 16473 42625 16476
rect 42659 16473 42671 16507
rect 42613 16467 42671 16473
rect 38289 16439 38347 16445
rect 38289 16436 38301 16439
rect 37976 16408 38301 16436
rect 37976 16396 37982 16408
rect 38289 16405 38301 16408
rect 38335 16405 38347 16439
rect 38289 16399 38347 16405
rect 38841 16439 38899 16445
rect 38841 16405 38853 16439
rect 38887 16405 38899 16439
rect 38841 16399 38899 16405
rect 41046 16396 41052 16448
rect 41104 16396 41110 16448
rect 42794 16396 42800 16448
rect 42852 16436 42858 16448
rect 42981 16439 43039 16445
rect 42981 16436 42993 16439
rect 42852 16408 42993 16436
rect 42852 16396 42858 16408
rect 42981 16405 42993 16408
rect 43027 16405 43039 16439
rect 42981 16399 43039 16405
rect 1104 16346 43884 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 43884 16346
rect 1104 16272 43884 16294
rect 14642 16192 14648 16244
rect 14700 16192 14706 16244
rect 15562 16192 15568 16244
rect 15620 16192 15626 16244
rect 15933 16235 15991 16241
rect 15933 16201 15945 16235
rect 15979 16232 15991 16235
rect 17310 16232 17316 16244
rect 15979 16204 17316 16232
rect 15979 16201 15991 16204
rect 15933 16195 15991 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 18138 16232 18144 16244
rect 17451 16204 18144 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 19484 16204 19625 16232
rect 19484 16192 19490 16204
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 19613 16195 19671 16201
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 21450 16232 21456 16244
rect 21131 16204 21456 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 22186 16192 22192 16244
rect 22244 16232 22250 16244
rect 22373 16235 22431 16241
rect 22373 16232 22385 16235
rect 22244 16204 22385 16232
rect 22244 16192 22250 16204
rect 22373 16201 22385 16204
rect 22419 16232 22431 16235
rect 22738 16232 22744 16244
rect 22419 16204 22744 16232
rect 22419 16201 22431 16204
rect 22373 16195 22431 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 26602 16192 26608 16244
rect 26660 16192 26666 16244
rect 27614 16192 27620 16244
rect 27672 16192 27678 16244
rect 34974 16232 34980 16244
rect 28092 16204 34980 16232
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 13510 16167 13568 16173
rect 13510 16164 13522 16167
rect 13044 16136 13522 16164
rect 13044 16124 13050 16136
rect 13510 16133 13522 16136
rect 13556 16133 13568 16167
rect 13510 16127 13568 16133
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15804 16136 16037 16164
rect 15804 16124 15810 16136
rect 16025 16133 16037 16136
rect 16071 16164 16083 16167
rect 16942 16164 16948 16176
rect 16071 16136 16948 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 18506 16124 18512 16176
rect 18564 16173 18570 16176
rect 18564 16164 18576 16173
rect 22465 16167 22523 16173
rect 18564 16136 18609 16164
rect 18564 16127 18576 16136
rect 22465 16133 22477 16167
rect 22511 16164 22523 16167
rect 22646 16164 22652 16176
rect 22511 16136 22652 16164
rect 22511 16133 22523 16136
rect 22465 16127 22523 16133
rect 18564 16124 18570 16127
rect 22646 16124 22652 16136
rect 22704 16124 22710 16176
rect 28092 16173 28120 16204
rect 34974 16192 34980 16204
rect 35032 16192 35038 16244
rect 36357 16235 36415 16241
rect 36357 16201 36369 16235
rect 36403 16232 36415 16235
rect 36722 16232 36728 16244
rect 36403 16204 36728 16232
rect 36403 16201 36415 16204
rect 36357 16195 36415 16201
rect 36722 16192 36728 16204
rect 36780 16192 36786 16244
rect 36909 16235 36967 16241
rect 36909 16201 36921 16235
rect 36955 16232 36967 16235
rect 37182 16232 37188 16244
rect 36955 16204 37188 16232
rect 36955 16201 36967 16204
rect 36909 16195 36967 16201
rect 37182 16192 37188 16204
rect 37240 16192 37246 16244
rect 38654 16192 38660 16244
rect 38712 16192 38718 16244
rect 40954 16192 40960 16244
rect 41012 16232 41018 16244
rect 42061 16235 42119 16241
rect 42061 16232 42073 16235
rect 41012 16204 42073 16232
rect 41012 16192 41018 16204
rect 42061 16201 42073 16204
rect 42107 16232 42119 16235
rect 43073 16235 43131 16241
rect 43073 16232 43085 16235
rect 42107 16204 43085 16232
rect 42107 16201 42119 16204
rect 42061 16195 42119 16201
rect 43073 16201 43085 16204
rect 43119 16201 43131 16235
rect 43073 16195 43131 16201
rect 25492 16167 25550 16173
rect 25492 16133 25504 16167
rect 25538 16164 25550 16167
rect 28077 16167 28135 16173
rect 25538 16136 28028 16164
rect 25538 16133 25550 16136
rect 25492 16127 25550 16133
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13354 16096 13360 16108
rect 13311 16068 13360 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13354 16056 13360 16068
rect 13412 16096 13418 16108
rect 15102 16096 15108 16108
rect 13412 16068 15108 16096
rect 13412 16056 13418 16068
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18785 16099 18843 16105
rect 17736 16068 18736 16096
rect 17736 16056 17742 16068
rect 16206 15988 16212 16040
rect 16264 15988 16270 16040
rect 18708 16028 18736 16068
rect 18785 16065 18797 16099
rect 18831 16096 18843 16099
rect 19150 16096 19156 16108
rect 18831 16068 19156 16096
rect 18831 16065 18843 16068
rect 18785 16059 18843 16065
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 21177 16099 21235 16105
rect 21177 16065 21189 16099
rect 21223 16096 21235 16099
rect 22370 16096 22376 16108
rect 21223 16068 22376 16096
rect 21223 16065 21235 16068
rect 21177 16059 21235 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 23201 16099 23259 16105
rect 23201 16065 23213 16099
rect 23247 16096 23259 16099
rect 23382 16096 23388 16108
rect 23247 16068 23388 16096
rect 23247 16065 23259 16068
rect 23201 16059 23259 16065
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 27798 16056 27804 16108
rect 27856 16056 27862 16108
rect 28000 16096 28028 16136
rect 28077 16133 28089 16167
rect 28123 16133 28135 16167
rect 32493 16167 32551 16173
rect 32493 16164 32505 16167
rect 28077 16127 28135 16133
rect 28920 16136 32505 16164
rect 28920 16105 28948 16136
rect 32493 16133 32505 16136
rect 32539 16164 32551 16167
rect 33321 16167 33379 16173
rect 33321 16164 33333 16167
rect 32539 16136 33333 16164
rect 32539 16133 32551 16136
rect 32493 16127 32551 16133
rect 33321 16133 33333 16136
rect 33367 16133 33379 16167
rect 33321 16127 33379 16133
rect 34606 16124 34612 16176
rect 34664 16124 34670 16176
rect 36170 16124 36176 16176
rect 36228 16124 36234 16176
rect 36740 16164 36768 16192
rect 39206 16164 39212 16176
rect 36740 16136 39212 16164
rect 39206 16124 39212 16136
rect 39264 16124 39270 16176
rect 42981 16167 43039 16173
rect 42981 16133 42993 16167
rect 43027 16164 43039 16167
rect 43162 16164 43168 16176
rect 43027 16136 43168 16164
rect 43027 16133 43039 16136
rect 42981 16127 43039 16133
rect 43162 16124 43168 16136
rect 43220 16124 43226 16176
rect 28905 16099 28963 16105
rect 28905 16096 28917 16099
rect 28000 16068 28917 16096
rect 28905 16065 28917 16068
rect 28951 16065 28963 16099
rect 28905 16059 28963 16065
rect 28997 16099 29055 16105
rect 28997 16065 29009 16099
rect 29043 16096 29055 16099
rect 29178 16096 29184 16108
rect 29043 16068 29184 16096
rect 29043 16065 29055 16068
rect 28997 16059 29055 16065
rect 29178 16056 29184 16068
rect 29236 16056 29242 16108
rect 29816 16099 29874 16105
rect 29816 16065 29828 16099
rect 29862 16096 29874 16099
rect 30098 16096 30104 16108
rect 29862 16068 30104 16096
rect 29862 16065 29874 16068
rect 29816 16059 29874 16065
rect 30098 16056 30104 16068
rect 30156 16056 30162 16108
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 30576 16068 31585 16096
rect 21266 16028 21272 16040
rect 18708 16000 21272 16028
rect 21266 15988 21272 16000
rect 21324 15988 21330 16040
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 19392 15932 20085 15960
rect 19392 15920 19398 15932
rect 20073 15929 20085 15932
rect 20119 15960 20131 15963
rect 21634 15960 21640 15972
rect 20119 15932 21640 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 21634 15920 21640 15932
rect 21692 15960 21698 15972
rect 22572 15960 22600 15991
rect 25130 15988 25136 16040
rect 25188 16028 25194 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 25188 16000 25237 16028
rect 25188 15988 25194 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 27246 15988 27252 16040
rect 27304 16028 27310 16040
rect 27893 16031 27951 16037
rect 27893 16028 27905 16031
rect 27304 16000 27905 16028
rect 27304 15988 27310 16000
rect 27893 15997 27905 16000
rect 27939 16028 27951 16031
rect 27939 16000 29500 16028
rect 27939 15997 27951 16000
rect 27893 15991 27951 15997
rect 21692 15932 22600 15960
rect 21692 15920 21698 15932
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 20312 15864 20729 15892
rect 20312 15852 20318 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 22002 15852 22008 15904
rect 22060 15852 22066 15904
rect 23385 15895 23443 15901
rect 23385 15861 23397 15895
rect 23431 15892 23443 15895
rect 23658 15892 23664 15904
rect 23431 15864 23664 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 28074 15852 28080 15904
rect 28132 15852 28138 15904
rect 29472 15892 29500 16000
rect 29546 15988 29552 16040
rect 29604 15988 29610 16040
rect 30576 15892 30604 16068
rect 31573 16065 31585 16068
rect 31619 16096 31631 16099
rect 31662 16096 31668 16108
rect 31619 16068 31668 16096
rect 31619 16065 31631 16068
rect 31573 16059 31631 16065
rect 31662 16056 31668 16068
rect 31720 16056 31726 16108
rect 31757 16099 31815 16105
rect 31757 16065 31769 16099
rect 31803 16065 31815 16099
rect 31757 16059 31815 16065
rect 30929 15963 30987 15969
rect 30929 15929 30941 15963
rect 30975 15960 30987 15963
rect 31570 15960 31576 15972
rect 30975 15932 31576 15960
rect 30975 15929 30987 15932
rect 30929 15923 30987 15929
rect 31570 15920 31576 15932
rect 31628 15960 31634 15972
rect 31772 15960 31800 16059
rect 32306 16056 32312 16108
rect 32364 16056 32370 16108
rect 33137 16099 33195 16105
rect 33137 16065 33149 16099
rect 33183 16096 33195 16099
rect 33226 16096 33232 16108
rect 33183 16068 33232 16096
rect 33183 16065 33195 16068
rect 33137 16059 33195 16065
rect 33226 16056 33232 16068
rect 33284 16056 33290 16108
rect 33410 16056 33416 16108
rect 33468 16096 33474 16108
rect 33870 16096 33876 16108
rect 33468 16068 33876 16096
rect 33468 16056 33474 16068
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 35986 16056 35992 16108
rect 36044 16056 36050 16108
rect 38194 16056 38200 16108
rect 38252 16056 38258 16108
rect 38378 16056 38384 16108
rect 38436 16056 38442 16108
rect 38470 16056 38476 16108
rect 38528 16056 38534 16108
rect 39298 16056 39304 16108
rect 39356 16056 39362 16108
rect 40948 16099 41006 16105
rect 40948 16065 40960 16099
rect 40994 16096 41006 16099
rect 41230 16096 41236 16108
rect 40994 16068 41236 16096
rect 40994 16065 41006 16068
rect 40948 16059 41006 16065
rect 41230 16056 41236 16068
rect 41288 16056 41294 16108
rect 31938 15988 31944 16040
rect 31996 16028 32002 16040
rect 34241 16031 34299 16037
rect 34241 16028 34253 16031
rect 31996 16000 34253 16028
rect 31996 15988 32002 16000
rect 34241 15997 34253 16000
rect 34287 15997 34299 16031
rect 34241 15991 34299 15997
rect 34330 15988 34336 16040
rect 34388 16028 34394 16040
rect 34425 16031 34483 16037
rect 34425 16028 34437 16031
rect 34388 16000 34437 16028
rect 34388 15988 34394 16000
rect 34425 15997 34437 16000
rect 34471 15997 34483 16031
rect 34425 15991 34483 15997
rect 35894 15988 35900 16040
rect 35952 16028 35958 16040
rect 37461 16031 37519 16037
rect 37461 16028 37473 16031
rect 35952 16000 37473 16028
rect 35952 15988 35958 16000
rect 37461 15997 37473 16000
rect 37507 15997 37519 16031
rect 37461 15991 37519 15997
rect 38289 16031 38347 16037
rect 38289 15997 38301 16031
rect 38335 16028 38347 16031
rect 39117 16031 39175 16037
rect 39117 16028 39129 16031
rect 38335 16000 39129 16028
rect 38335 15997 38347 16000
rect 38289 15991 38347 15997
rect 39117 15997 39129 16000
rect 39163 15997 39175 16031
rect 39117 15991 39175 15997
rect 39577 16031 39635 16037
rect 39577 15997 39589 16031
rect 39623 16028 39635 16031
rect 39850 16028 39856 16040
rect 39623 16000 39856 16028
rect 39623 15997 39635 16000
rect 39577 15991 39635 15997
rect 39850 15988 39856 16000
rect 39908 15988 39914 16040
rect 40681 16031 40739 16037
rect 40681 15997 40693 16031
rect 40727 15997 40739 16031
rect 40681 15991 40739 15997
rect 43165 16031 43223 16037
rect 43165 15997 43177 16031
rect 43211 15997 43223 16031
rect 43165 15991 43223 15997
rect 31628 15932 31800 15960
rect 31628 15920 31634 15932
rect 33226 15920 33232 15972
rect 33284 15960 33290 15972
rect 34348 15960 34376 15988
rect 34790 15960 34796 15972
rect 33284 15932 34376 15960
rect 34532 15932 34796 15960
rect 33284 15920 33290 15932
rect 29472 15864 30604 15892
rect 31386 15852 31392 15904
rect 31444 15852 31450 15904
rect 32677 15895 32735 15901
rect 32677 15861 32689 15895
rect 32723 15892 32735 15895
rect 32766 15892 32772 15904
rect 32723 15864 32772 15892
rect 32723 15861 32735 15864
rect 32677 15855 32735 15861
rect 32766 15852 32772 15864
rect 32824 15852 32830 15904
rect 33134 15852 33140 15904
rect 33192 15852 33198 15904
rect 34333 15895 34391 15901
rect 34333 15861 34345 15895
rect 34379 15892 34391 15895
rect 34532 15892 34560 15932
rect 34790 15920 34796 15932
rect 34848 15920 34854 15972
rect 34974 15920 34980 15972
rect 35032 15960 35038 15972
rect 36722 15960 36728 15972
rect 35032 15932 36728 15960
rect 35032 15920 35038 15932
rect 36722 15920 36728 15932
rect 36780 15960 36786 15972
rect 37274 15960 37280 15972
rect 36780 15932 37280 15960
rect 36780 15920 36786 15932
rect 37274 15920 37280 15932
rect 37332 15960 37338 15972
rect 37918 15960 37924 15972
rect 37332 15932 37924 15960
rect 37332 15920 37338 15932
rect 37918 15920 37924 15932
rect 37976 15920 37982 15972
rect 34379 15864 34560 15892
rect 34379 15861 34391 15864
rect 34333 15855 34391 15861
rect 34606 15852 34612 15904
rect 34664 15852 34670 15904
rect 35158 15852 35164 15904
rect 35216 15892 35222 15904
rect 35529 15895 35587 15901
rect 35529 15892 35541 15895
rect 35216 15864 35541 15892
rect 35216 15852 35222 15864
rect 35529 15861 35541 15864
rect 35575 15892 35587 15895
rect 37182 15892 37188 15904
rect 35575 15864 37188 15892
rect 35575 15861 35587 15864
rect 35529 15855 35587 15861
rect 37182 15852 37188 15864
rect 37240 15852 37246 15904
rect 39022 15852 39028 15904
rect 39080 15892 39086 15904
rect 39485 15895 39543 15901
rect 39485 15892 39497 15895
rect 39080 15864 39497 15892
rect 39080 15852 39086 15864
rect 39485 15861 39497 15864
rect 39531 15861 39543 15895
rect 39485 15855 39543 15861
rect 40129 15895 40187 15901
rect 40129 15861 40141 15895
rect 40175 15892 40187 15895
rect 40218 15892 40224 15904
rect 40175 15864 40224 15892
rect 40175 15861 40187 15864
rect 40129 15855 40187 15861
rect 40218 15852 40224 15864
rect 40276 15852 40282 15904
rect 40696 15892 40724 15991
rect 42978 15920 42984 15972
rect 43036 15960 43042 15972
rect 43180 15960 43208 15991
rect 43036 15932 43208 15960
rect 43036 15920 43042 15932
rect 41322 15892 41328 15904
rect 40696 15864 41328 15892
rect 41322 15852 41328 15864
rect 41380 15852 41386 15904
rect 41598 15852 41604 15904
rect 41656 15892 41662 15904
rect 42613 15895 42671 15901
rect 42613 15892 42625 15895
rect 41656 15864 42625 15892
rect 41656 15852 41662 15864
rect 42613 15861 42625 15864
rect 42659 15861 42671 15895
rect 42613 15855 42671 15861
rect 1104 15802 43884 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 43884 15802
rect 1104 15728 43884 15750
rect 16485 15691 16543 15697
rect 16485 15657 16497 15691
rect 16531 15688 16543 15691
rect 17310 15688 17316 15700
rect 16531 15660 17316 15688
rect 16531 15657 16543 15660
rect 16485 15651 16543 15657
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 18598 15648 18604 15700
rect 18656 15648 18662 15700
rect 22186 15648 22192 15700
rect 22244 15648 22250 15700
rect 23382 15648 23388 15700
rect 23440 15648 23446 15700
rect 27246 15648 27252 15700
rect 27304 15688 27310 15700
rect 27433 15691 27491 15697
rect 27433 15688 27445 15691
rect 27304 15660 27445 15688
rect 27304 15648 27310 15660
rect 27433 15657 27445 15660
rect 27479 15657 27491 15691
rect 27433 15651 27491 15657
rect 27890 15648 27896 15700
rect 27948 15688 27954 15700
rect 28169 15691 28227 15697
rect 28169 15688 28181 15691
rect 27948 15660 28181 15688
rect 27948 15648 27954 15660
rect 28169 15657 28181 15660
rect 28215 15657 28227 15691
rect 28169 15651 28227 15657
rect 30098 15648 30104 15700
rect 30156 15648 30162 15700
rect 31205 15691 31263 15697
rect 31205 15657 31217 15691
rect 31251 15688 31263 15691
rect 31478 15688 31484 15700
rect 31251 15660 31484 15688
rect 31251 15657 31263 15660
rect 31205 15651 31263 15657
rect 31478 15648 31484 15660
rect 31536 15648 31542 15700
rect 31754 15648 31760 15700
rect 31812 15648 31818 15700
rect 32858 15688 32864 15700
rect 32600 15660 32864 15688
rect 26234 15620 26240 15632
rect 25976 15592 26240 15620
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 16264 15524 17969 15552
rect 16264 15512 16270 15524
rect 17957 15521 17969 15524
rect 18003 15552 18015 15555
rect 19058 15552 19064 15564
rect 18003 15524 19064 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 20254 15552 20260 15564
rect 19536 15524 20260 15552
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14476 15416 14504 15447
rect 15102 15444 15108 15496
rect 15160 15444 15166 15496
rect 15372 15487 15430 15493
rect 15372 15453 15384 15487
rect 15418 15484 15430 15487
rect 15654 15484 15660 15496
rect 15418 15456 15660 15484
rect 15418 15453 15430 15456
rect 15372 15447 15430 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 16942 15444 16948 15496
rect 17000 15444 17006 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 19536 15493 19564 15524
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20809 15555 20867 15561
rect 20809 15552 20821 15555
rect 20772 15524 20821 15552
rect 20772 15512 20778 15524
rect 20809 15521 20821 15524
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 22370 15512 22376 15564
rect 22428 15552 22434 15564
rect 22741 15555 22799 15561
rect 22741 15552 22753 15555
rect 22428 15524 22753 15552
rect 22428 15512 22434 15524
rect 22741 15521 22753 15524
rect 22787 15552 22799 15555
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 22787 15524 23857 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 25976 15561 26004 15592
rect 26234 15580 26240 15592
rect 26292 15620 26298 15632
rect 26513 15623 26571 15629
rect 26513 15620 26525 15623
rect 26292 15592 26525 15620
rect 26292 15580 26298 15592
rect 26513 15589 26525 15592
rect 26559 15620 26571 15623
rect 30006 15620 30012 15632
rect 26559 15592 30012 15620
rect 26559 15589 26571 15592
rect 26513 15583 26571 15589
rect 30006 15580 30012 15592
rect 30064 15580 30070 15632
rect 32600 15620 32628 15660
rect 32858 15648 32864 15660
rect 32916 15688 32922 15700
rect 35805 15691 35863 15697
rect 32916 15660 33732 15688
rect 32916 15648 32922 15660
rect 33134 15620 33140 15632
rect 30484 15592 32628 15620
rect 32692 15592 33140 15620
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 25740 15524 25789 15552
rect 25740 15512 25746 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 25961 15555 26019 15561
rect 25961 15521 25973 15555
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 28074 15512 28080 15564
rect 28132 15552 28138 15564
rect 29914 15552 29920 15564
rect 28132 15524 29920 15552
rect 28132 15512 28138 15524
rect 29914 15512 29920 15524
rect 29972 15552 29978 15564
rect 30484 15552 30512 15592
rect 29972 15524 30512 15552
rect 30561 15555 30619 15561
rect 29972 15512 29978 15524
rect 30561 15521 30573 15555
rect 30607 15552 30619 15555
rect 31386 15552 31392 15564
rect 30607 15524 31392 15552
rect 30607 15521 30619 15524
rect 30561 15515 30619 15521
rect 31386 15512 31392 15524
rect 31444 15512 31450 15564
rect 32692 15561 32720 15592
rect 33134 15580 33140 15592
rect 33192 15580 33198 15632
rect 32677 15555 32735 15561
rect 32677 15521 32689 15555
rect 32723 15521 32735 15555
rect 32677 15515 32735 15521
rect 32766 15512 32772 15564
rect 32824 15512 32830 15564
rect 32858 15512 32864 15564
rect 32916 15552 32922 15564
rect 33597 15555 33655 15561
rect 33597 15552 33609 15555
rect 32916 15524 33609 15552
rect 32916 15512 32922 15524
rect 33597 15521 33609 15524
rect 33643 15521 33655 15555
rect 33597 15515 33655 15521
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18196 15456 18245 15484
rect 18196 15444 18202 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15484 20223 15487
rect 22002 15484 22008 15496
rect 20211 15456 22008 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22830 15444 22836 15496
rect 22888 15484 22894 15496
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22888 15456 23029 15484
rect 22888 15444 22894 15456
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15484 28411 15487
rect 28534 15484 28540 15496
rect 28399 15456 28540 15484
rect 28399 15453 28411 15456
rect 28353 15447 28411 15453
rect 28534 15444 28540 15456
rect 28592 15484 28598 15496
rect 28902 15484 28908 15496
rect 28592 15456 28908 15484
rect 28592 15444 28598 15456
rect 28902 15444 28908 15456
rect 28960 15444 28966 15496
rect 30282 15444 30288 15496
rect 30340 15444 30346 15496
rect 30377 15487 30435 15493
rect 30377 15453 30389 15487
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 30469 15487 30527 15493
rect 30469 15453 30481 15487
rect 30515 15484 30527 15487
rect 31110 15484 31116 15496
rect 30515 15456 31116 15484
rect 30515 15453 30527 15456
rect 30469 15447 30527 15453
rect 15286 15416 15292 15428
rect 14476 15388 15292 15416
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 21054 15419 21112 15425
rect 21054 15416 21066 15419
rect 20364 15388 21066 15416
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 17126 15308 17132 15360
rect 17184 15308 17190 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18141 15351 18199 15357
rect 18141 15348 18153 15351
rect 18012 15320 18153 15348
rect 18012 15308 18018 15320
rect 18141 15317 18153 15320
rect 18187 15317 18199 15351
rect 18141 15311 18199 15317
rect 19705 15351 19763 15357
rect 19705 15317 19717 15351
rect 19751 15348 19763 15351
rect 20070 15348 20076 15360
rect 19751 15320 20076 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20364 15357 20392 15388
rect 21054 15385 21066 15388
rect 21100 15385 21112 15419
rect 21054 15379 21112 15385
rect 22646 15376 22652 15428
rect 22704 15416 22710 15428
rect 22925 15419 22983 15425
rect 22925 15416 22937 15419
rect 22704 15388 22937 15416
rect 22704 15376 22710 15388
rect 22925 15385 22937 15388
rect 22971 15385 22983 15419
rect 30392 15416 30420 15447
rect 31110 15444 31116 15456
rect 31168 15444 31174 15496
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 32953 15487 33011 15493
rect 32953 15484 32965 15487
rect 31812 15456 32965 15484
rect 31812 15444 31818 15456
rect 32953 15453 32965 15456
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 33502 15444 33508 15496
rect 33560 15444 33566 15496
rect 33704 15493 33732 15660
rect 35805 15657 35817 15691
rect 35851 15688 35863 15691
rect 35894 15688 35900 15700
rect 35851 15660 35900 15688
rect 35851 15657 35863 15660
rect 35805 15651 35863 15657
rect 35894 15648 35900 15660
rect 35952 15648 35958 15700
rect 36357 15691 36415 15697
rect 36357 15657 36369 15691
rect 36403 15688 36415 15691
rect 36630 15688 36636 15700
rect 36403 15660 36636 15688
rect 36403 15657 36415 15660
rect 36357 15651 36415 15657
rect 36630 15648 36636 15660
rect 36688 15648 36694 15700
rect 38194 15648 38200 15700
rect 38252 15648 38258 15700
rect 42886 15648 42892 15700
rect 42944 15688 42950 15700
rect 43349 15691 43407 15697
rect 43349 15688 43361 15691
rect 42944 15660 43361 15688
rect 42944 15648 42950 15660
rect 43349 15657 43361 15660
rect 43395 15657 43407 15691
rect 43349 15651 43407 15657
rect 38930 15620 38936 15632
rect 36188 15592 38936 15620
rect 35342 15552 35348 15564
rect 35084 15524 35348 15552
rect 33689 15487 33747 15493
rect 33689 15453 33701 15487
rect 33735 15484 33747 15487
rect 34149 15487 34207 15493
rect 34149 15484 34161 15487
rect 33735 15456 34161 15484
rect 33735 15453 33747 15456
rect 33689 15447 33747 15453
rect 34149 15453 34161 15456
rect 34195 15484 34207 15487
rect 34238 15484 34244 15496
rect 34195 15456 34244 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 34238 15444 34244 15456
rect 34296 15444 34302 15496
rect 34333 15487 34391 15493
rect 34333 15453 34345 15487
rect 34379 15484 34391 15487
rect 34514 15484 34520 15496
rect 34379 15456 34520 15484
rect 34379 15453 34391 15456
rect 34333 15447 34391 15453
rect 34514 15444 34520 15456
rect 34572 15444 34578 15496
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 35084 15493 35112 15524
rect 35342 15512 35348 15524
rect 35400 15512 35406 15564
rect 35069 15487 35127 15493
rect 34756 15456 35020 15484
rect 34756 15444 34762 15456
rect 34790 15416 34796 15428
rect 30392 15388 34796 15416
rect 22925 15379 22983 15385
rect 34790 15376 34796 15388
rect 34848 15416 34854 15428
rect 34885 15419 34943 15425
rect 34885 15416 34897 15419
rect 34848 15388 34897 15416
rect 34848 15376 34854 15388
rect 34885 15385 34897 15388
rect 34931 15385 34943 15419
rect 34992 15416 35020 15456
rect 35069 15453 35081 15487
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15453 35311 15487
rect 35253 15447 35311 15453
rect 35268 15416 35296 15447
rect 35526 15444 35532 15496
rect 35584 15484 35590 15496
rect 36188 15484 36216 15592
rect 36262 15512 36268 15564
rect 36320 15552 36326 15564
rect 36725 15555 36783 15561
rect 36725 15552 36737 15555
rect 36320 15524 36737 15552
rect 36320 15512 36326 15524
rect 36725 15521 36737 15524
rect 36771 15552 36783 15555
rect 37182 15552 37188 15564
rect 36771 15524 37188 15552
rect 36771 15521 36783 15524
rect 36725 15515 36783 15521
rect 37182 15512 37188 15524
rect 37240 15512 37246 15564
rect 36541 15487 36599 15493
rect 36541 15484 36553 15487
rect 35584 15456 36553 15484
rect 35584 15444 35590 15456
rect 36541 15453 36553 15456
rect 36587 15453 36599 15487
rect 36541 15447 36599 15453
rect 36630 15444 36636 15496
rect 36688 15444 36694 15496
rect 36814 15444 36820 15496
rect 36872 15444 36878 15496
rect 37660 15493 37688 15592
rect 38930 15580 38936 15592
rect 38988 15580 38994 15632
rect 38378 15552 38384 15564
rect 37752 15524 38384 15552
rect 37752 15493 37780 15524
rect 38378 15512 38384 15524
rect 38436 15512 38442 15564
rect 40954 15512 40960 15564
rect 41012 15512 41018 15564
rect 41138 15512 41144 15564
rect 41196 15552 41202 15564
rect 41690 15552 41696 15564
rect 41196 15524 41696 15552
rect 41196 15512 41202 15524
rect 41690 15512 41696 15524
rect 41748 15512 41754 15564
rect 41966 15512 41972 15564
rect 42024 15512 42030 15564
rect 37645 15487 37703 15493
rect 37645 15453 37657 15487
rect 37691 15453 37703 15487
rect 37645 15447 37703 15453
rect 37737 15487 37795 15493
rect 37737 15453 37749 15487
rect 37783 15453 37795 15487
rect 37737 15447 37795 15453
rect 37918 15444 37924 15496
rect 37976 15444 37982 15496
rect 38013 15487 38071 15493
rect 38013 15453 38025 15487
rect 38059 15453 38071 15487
rect 38013 15447 38071 15453
rect 39117 15487 39175 15493
rect 39117 15453 39129 15487
rect 39163 15453 39175 15487
rect 39117 15447 39175 15453
rect 35618 15416 35624 15428
rect 34992 15388 35624 15416
rect 34885 15379 34943 15385
rect 35618 15376 35624 15388
rect 35676 15376 35682 15428
rect 36078 15376 36084 15428
rect 36136 15416 36142 15428
rect 38028 15416 38056 15447
rect 36136 15388 38056 15416
rect 39132 15416 39160 15447
rect 39206 15444 39212 15496
rect 39264 15444 39270 15496
rect 41322 15444 41328 15496
rect 41380 15484 41386 15496
rect 41984 15484 42012 15512
rect 43162 15484 43168 15496
rect 41380 15456 42012 15484
rect 42168 15456 43168 15484
rect 41380 15444 41386 15456
rect 40865 15419 40923 15425
rect 39132 15388 40632 15416
rect 36136 15376 36142 15388
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15317 20407 15351
rect 20349 15311 20407 15317
rect 25222 15308 25228 15360
rect 25280 15348 25286 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 25280 15320 25329 15348
rect 25280 15308 25286 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 26050 15348 26056 15360
rect 25731 15320 26056 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 26050 15308 26056 15320
rect 26108 15308 26114 15360
rect 27614 15308 27620 15360
rect 27672 15348 27678 15360
rect 27982 15348 27988 15360
rect 27672 15320 27988 15348
rect 27672 15308 27678 15320
rect 27982 15308 27988 15320
rect 28040 15348 28046 15360
rect 28813 15351 28871 15357
rect 28813 15348 28825 15351
rect 28040 15320 28825 15348
rect 28040 15308 28046 15320
rect 28813 15317 28825 15320
rect 28859 15317 28871 15351
rect 28813 15311 28871 15317
rect 32398 15308 32404 15360
rect 32456 15348 32462 15360
rect 32493 15351 32551 15357
rect 32493 15348 32505 15351
rect 32456 15320 32505 15348
rect 32456 15308 32462 15320
rect 32493 15317 32505 15320
rect 32539 15317 32551 15351
rect 32493 15311 32551 15317
rect 34146 15308 34152 15360
rect 34204 15308 34210 15360
rect 40494 15308 40500 15360
rect 40552 15308 40558 15360
rect 40604 15348 40632 15388
rect 40865 15385 40877 15419
rect 40911 15416 40923 15419
rect 42168 15416 42196 15456
rect 43162 15444 43168 15456
rect 43220 15444 43226 15496
rect 40911 15388 42196 15416
rect 42236 15419 42294 15425
rect 40911 15385 40923 15388
rect 40865 15379 40923 15385
rect 42236 15385 42248 15419
rect 42282 15416 42294 15419
rect 42610 15416 42616 15428
rect 42282 15388 42616 15416
rect 42282 15385 42294 15388
rect 42236 15379 42294 15385
rect 42610 15376 42616 15388
rect 42668 15376 42674 15428
rect 41046 15348 41052 15360
rect 40604 15320 41052 15348
rect 41046 15308 41052 15320
rect 41104 15308 41110 15360
rect 1104 15258 43884 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 43884 15258
rect 1104 15184 43884 15206
rect 14826 15104 14832 15156
rect 14884 15104 14890 15156
rect 15286 15104 15292 15156
rect 15344 15104 15350 15156
rect 15746 15104 15752 15156
rect 15804 15104 15810 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18104 15116 18245 15144
rect 18104 15104 18110 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 19153 15147 19211 15153
rect 19153 15113 19165 15147
rect 19199 15144 19211 15147
rect 19978 15144 19984 15156
rect 19199 15116 19984 15144
rect 19199 15113 19211 15116
rect 19153 15107 19211 15113
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 21361 15147 21419 15153
rect 21361 15113 21373 15147
rect 21407 15144 21419 15147
rect 21450 15144 21456 15156
rect 21407 15116 21456 15144
rect 21407 15113 21419 15116
rect 21361 15107 21419 15113
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 22557 15147 22615 15153
rect 22557 15113 22569 15147
rect 22603 15144 22615 15147
rect 22830 15144 22836 15156
rect 22603 15116 22836 15144
rect 22603 15113 22615 15116
rect 22557 15107 22615 15113
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 28718 15104 28724 15156
rect 28776 15144 28782 15156
rect 28905 15147 28963 15153
rect 28905 15144 28917 15147
rect 28776 15116 28917 15144
rect 28776 15104 28782 15116
rect 28905 15113 28917 15116
rect 28951 15113 28963 15147
rect 28905 15107 28963 15113
rect 29086 15104 29092 15156
rect 29144 15144 29150 15156
rect 29457 15147 29515 15153
rect 29457 15144 29469 15147
rect 29144 15116 29469 15144
rect 29144 15104 29150 15116
rect 29457 15113 29469 15116
rect 29503 15113 29515 15147
rect 29457 15107 29515 15113
rect 31754 15104 31760 15156
rect 31812 15144 31818 15156
rect 32309 15147 32367 15153
rect 32309 15144 32321 15147
rect 31812 15116 32321 15144
rect 31812 15104 31818 15116
rect 32309 15113 32321 15116
rect 32355 15113 32367 15147
rect 32309 15107 32367 15113
rect 35161 15147 35219 15153
rect 35161 15113 35173 15147
rect 35207 15144 35219 15147
rect 35434 15144 35440 15156
rect 35207 15116 35440 15144
rect 35207 15113 35219 15116
rect 35161 15107 35219 15113
rect 35434 15104 35440 15116
rect 35492 15104 35498 15156
rect 36814 15104 36820 15156
rect 36872 15144 36878 15156
rect 36909 15147 36967 15153
rect 36909 15144 36921 15147
rect 36872 15116 36921 15144
rect 36872 15104 36878 15116
rect 36909 15113 36921 15116
rect 36955 15113 36967 15147
rect 36909 15107 36967 15113
rect 37090 15104 37096 15156
rect 37148 15144 37154 15156
rect 38289 15147 38347 15153
rect 37148 15116 38056 15144
rect 37148 15104 37154 15116
rect 15102 15036 15108 15088
rect 15160 15076 15166 15088
rect 20714 15076 20720 15088
rect 15160 15048 19196 15076
rect 15160 15036 15166 15048
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 13412 14980 13461 15008
rect 13412 14968 13418 14980
rect 13449 14977 13461 14980
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13716 15011 13774 15017
rect 13716 14977 13728 15011
rect 13762 15008 13774 15011
rect 14274 15008 14280 15020
rect 13762 14980 14280 15008
rect 13762 14977 13774 14980
rect 13716 14971 13774 14977
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 16868 15017 16896 15048
rect 19168 15020 19196 15048
rect 19996 15048 20720 15076
rect 17126 15017 17132 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 14884 14980 15669 15008
rect 14884 14968 14890 14980
rect 15657 14977 15669 14980
rect 15703 14977 15715 15011
rect 15657 14971 15715 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 17120 15008 17132 15017
rect 17087 14980 17132 15008
rect 16853 14971 16911 14977
rect 17120 14971 17132 14980
rect 17126 14968 17132 14971
rect 17184 14968 17190 15020
rect 19150 14968 19156 15020
rect 19208 15008 19214 15020
rect 19996 15017 20024 15048
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 23658 15036 23664 15088
rect 23716 15085 23722 15088
rect 23716 15076 23728 15085
rect 23716 15048 23761 15076
rect 23716 15039 23728 15048
rect 23716 15036 23722 15039
rect 27338 15036 27344 15088
rect 27396 15076 27402 15088
rect 27801 15079 27859 15085
rect 27801 15076 27813 15079
rect 27396 15048 27813 15076
rect 27396 15036 27402 15048
rect 27801 15045 27813 15048
rect 27847 15045 27859 15079
rect 27801 15039 27859 15045
rect 27893 15079 27951 15085
rect 27893 15045 27905 15079
rect 27939 15076 27951 15079
rect 29270 15076 29276 15088
rect 27939 15048 29276 15076
rect 27939 15045 27951 15048
rect 27893 15039 27951 15045
rect 29270 15036 29276 15048
rect 29328 15036 29334 15088
rect 32766 15036 32772 15088
rect 32824 15076 32830 15088
rect 33318 15076 33324 15088
rect 32824 15048 33324 15076
rect 32824 15036 32830 15048
rect 33318 15036 33324 15048
rect 33376 15036 33382 15088
rect 34698 15085 34704 15088
rect 34675 15079 34704 15085
rect 34675 15045 34687 15079
rect 34675 15039 34704 15045
rect 34698 15036 34704 15039
rect 34756 15036 34762 15088
rect 35066 15076 35072 15088
rect 34808 15048 35072 15076
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19208 14980 19993 15008
rect 19208 14968 19214 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 24946 15017 24952 15020
rect 20237 15011 20295 15017
rect 20237 15008 20249 15011
rect 20128 14980 20249 15008
rect 20128 14968 20134 14980
rect 20237 14977 20249 14980
rect 20283 14977 20295 15011
rect 20237 14971 20295 14977
rect 24940 14971 24952 15017
rect 24946 14968 24952 14971
rect 25004 14968 25010 15020
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 27709 15011 27767 15017
rect 27709 15008 27721 15011
rect 27672 14980 27721 15008
rect 27672 14968 27678 14980
rect 27709 14977 27721 14980
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28537 15011 28595 15017
rect 28537 15008 28549 15011
rect 28123 14980 28549 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28537 14977 28549 14980
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28721 15011 28779 15017
rect 28721 14977 28733 15011
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 15010 14900 15016 14952
rect 15068 14940 15074 14952
rect 15930 14940 15936 14952
rect 15068 14912 15936 14940
rect 15068 14900 15074 14912
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18064 14912 18889 14940
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 18064 14804 18092 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14940 19119 14943
rect 19107 14912 19932 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 18892 14872 18920 14903
rect 19334 14872 19340 14884
rect 18892 14844 19340 14872
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 15528 14776 18092 14804
rect 15528 14764 15534 14776
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19521 14807 19579 14813
rect 19521 14804 19533 14807
rect 19484 14776 19533 14804
rect 19484 14764 19490 14776
rect 19521 14773 19533 14776
rect 19567 14773 19579 14807
rect 19904 14804 19932 14912
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 23992 14912 24685 14940
rect 23992 14900 23998 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 28736 14940 28764 14971
rect 28994 14968 29000 15020
rect 29052 14968 29058 15020
rect 29178 14968 29184 15020
rect 29236 15008 29242 15020
rect 29641 15011 29699 15017
rect 29641 15008 29653 15011
rect 29236 14980 29653 15008
rect 29236 14968 29242 14980
rect 29641 14977 29653 14980
rect 29687 14977 29699 15011
rect 29641 14971 29699 14977
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 15008 29975 15011
rect 31478 15008 31484 15020
rect 29963 14980 31484 15008
rect 29963 14977 29975 14980
rect 29917 14971 29975 14977
rect 31478 14968 31484 14980
rect 31536 14968 31542 15020
rect 33226 14968 33232 15020
rect 33284 15008 33290 15020
rect 34808 15017 34836 15048
rect 35066 15036 35072 15048
rect 35124 15036 35130 15088
rect 35894 15036 35900 15088
rect 35952 15076 35958 15088
rect 37918 15076 37924 15088
rect 35952 15048 37924 15076
rect 35952 15036 35958 15048
rect 37918 15036 37924 15048
rect 37976 15036 37982 15088
rect 33689 15011 33747 15017
rect 33689 15008 33701 15011
rect 33284 14980 33701 15008
rect 33284 14968 33290 14980
rect 33689 14977 33701 14980
rect 33735 14977 33747 15011
rect 33689 14971 33747 14977
rect 34793 15011 34851 15017
rect 34793 14977 34805 15011
rect 34839 14977 34851 15011
rect 34793 14971 34851 14977
rect 34882 14968 34888 15020
rect 34940 14968 34946 15020
rect 34977 15011 35035 15017
rect 34977 14977 34989 15011
rect 35023 14977 35035 15011
rect 34977 14971 35035 14977
rect 35813 15011 35871 15017
rect 35813 14977 35825 15011
rect 35859 15008 35871 15011
rect 35912 15008 35940 15036
rect 35859 14980 35940 15008
rect 35989 15011 36047 15017
rect 35859 14977 35871 14980
rect 35813 14971 35871 14977
rect 35989 14977 36001 15011
rect 36035 15008 36047 15011
rect 36354 15008 36360 15020
rect 36035 14980 36360 15008
rect 36035 14977 36047 14980
rect 35989 14971 36047 14977
rect 28736 14912 28994 14940
rect 24673 14903 24731 14909
rect 28966 14872 28994 14912
rect 29086 14900 29092 14952
rect 29144 14940 29150 14952
rect 29825 14943 29883 14949
rect 29825 14940 29837 14943
rect 29144 14912 29837 14940
rect 29144 14900 29150 14912
rect 29825 14909 29837 14912
rect 29871 14940 29883 14943
rect 29871 14912 31156 14940
rect 29871 14909 29883 14912
rect 29825 14903 29883 14909
rect 31128 14872 31156 14912
rect 34514 14900 34520 14952
rect 34572 14900 34578 14952
rect 34606 14872 34612 14884
rect 28966 14844 30328 14872
rect 31128 14844 34612 14872
rect 30300 14816 30328 14844
rect 34606 14832 34612 14844
rect 34664 14832 34670 14884
rect 34900 14872 34928 14968
rect 34992 14940 35020 14971
rect 36354 14968 36360 14980
rect 36412 14968 36418 15020
rect 36446 14968 36452 15020
rect 36504 14968 36510 15020
rect 36722 14968 36728 15020
rect 36780 15008 36786 15020
rect 36780 14980 37412 15008
rect 36780 14968 36786 14980
rect 35897 14943 35955 14949
rect 35897 14940 35909 14943
rect 34992 14912 35909 14940
rect 35897 14909 35909 14912
rect 35943 14909 35955 14943
rect 35897 14903 35955 14909
rect 35526 14872 35532 14884
rect 34900 14844 35532 14872
rect 35526 14832 35532 14844
rect 35584 14832 35590 14884
rect 36464 14872 36492 14968
rect 36633 14943 36691 14949
rect 36633 14909 36645 14943
rect 36679 14940 36691 14943
rect 37274 14940 37280 14952
rect 36679 14912 37280 14940
rect 36679 14909 36691 14912
rect 36633 14903 36691 14909
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 37384 14940 37412 14980
rect 37458 14968 37464 15020
rect 37516 14968 37522 15020
rect 37642 14968 37648 15020
rect 37700 14968 37706 15020
rect 38028 15008 38056 15116
rect 38289 15113 38301 15147
rect 38335 15144 38347 15147
rect 38378 15144 38384 15156
rect 38335 15116 38384 15144
rect 38335 15113 38347 15116
rect 38289 15107 38347 15113
rect 38378 15104 38384 15116
rect 38436 15104 38442 15156
rect 41230 15104 41236 15156
rect 41288 15144 41294 15156
rect 41325 15147 41383 15153
rect 41325 15144 41337 15147
rect 41288 15116 41337 15144
rect 41288 15104 41294 15116
rect 41325 15113 41337 15116
rect 41371 15113 41383 15147
rect 41325 15107 41383 15113
rect 41874 15104 41880 15156
rect 41932 15144 41938 15156
rect 41969 15147 42027 15153
rect 41969 15144 41981 15147
rect 41932 15116 41981 15144
rect 41932 15104 41938 15116
rect 41969 15113 41981 15116
rect 42015 15113 42027 15147
rect 41969 15107 42027 15113
rect 42610 15104 42616 15156
rect 42668 15104 42674 15156
rect 43346 15104 43352 15156
rect 43404 15104 43410 15156
rect 38102 15036 38108 15088
rect 38160 15076 38166 15088
rect 38473 15079 38531 15085
rect 38473 15076 38485 15079
rect 38160 15048 38485 15076
rect 38160 15036 38166 15048
rect 38473 15045 38485 15048
rect 38519 15045 38531 15079
rect 38473 15039 38531 15045
rect 38657 15079 38715 15085
rect 38657 15045 38669 15079
rect 38703 15076 38715 15079
rect 38746 15076 38752 15088
rect 38703 15048 38752 15076
rect 38703 15045 38715 15048
rect 38657 15039 38715 15045
rect 38746 15036 38752 15048
rect 38804 15036 38810 15088
rect 39577 15079 39635 15085
rect 39577 15045 39589 15079
rect 39623 15076 39635 15079
rect 40126 15076 40132 15088
rect 39623 15048 40132 15076
rect 39623 15045 39635 15048
rect 39577 15039 39635 15045
rect 40126 15036 40132 15048
rect 40184 15036 40190 15088
rect 39393 15011 39451 15017
rect 39393 15008 39405 15011
rect 38028 14980 39405 15008
rect 39393 14977 39405 14980
rect 39439 14977 39451 15011
rect 39393 14971 39451 14977
rect 39758 14968 39764 15020
rect 39816 14968 39822 15020
rect 40497 15011 40555 15017
rect 40497 14977 40509 15011
rect 40543 15008 40555 15011
rect 41046 15008 41052 15020
rect 40543 14980 41052 15008
rect 40543 14977 40555 14980
rect 40497 14971 40555 14977
rect 41046 14968 41052 14980
rect 41104 14968 41110 15020
rect 41509 15011 41567 15017
rect 41509 14977 41521 15011
rect 41555 15008 41567 15011
rect 41598 15008 41604 15020
rect 41555 14980 41604 15008
rect 41555 14977 41567 14980
rect 41509 14971 41567 14977
rect 41598 14968 41604 14980
rect 41656 14968 41662 15020
rect 42794 14968 42800 15020
rect 42852 14968 42858 15020
rect 39850 14940 39856 14952
rect 37384 14912 39856 14940
rect 39850 14900 39856 14912
rect 39908 14900 39914 14952
rect 36722 14872 36728 14884
rect 36464 14844 36728 14872
rect 36722 14832 36728 14844
rect 36780 14832 36786 14884
rect 39022 14872 39028 14884
rect 36832 14844 39028 14872
rect 20162 14804 20168 14816
rect 19904 14776 20168 14804
rect 19521 14767 19579 14773
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 27522 14764 27528 14816
rect 27580 14764 27586 14816
rect 28718 14764 28724 14816
rect 28776 14804 28782 14816
rect 29086 14804 29092 14816
rect 28776 14776 29092 14804
rect 28776 14764 28782 14776
rect 29086 14764 29092 14776
rect 29144 14764 29150 14816
rect 29730 14764 29736 14816
rect 29788 14764 29794 14816
rect 30282 14764 30288 14816
rect 30340 14804 30346 14816
rect 33137 14807 33195 14813
rect 33137 14804 33149 14807
rect 30340 14776 33149 14804
rect 30340 14764 30346 14776
rect 33137 14773 33149 14776
rect 33183 14773 33195 14807
rect 33137 14767 33195 14773
rect 33321 14807 33379 14813
rect 33321 14773 33333 14807
rect 33367 14804 33379 14807
rect 33410 14804 33416 14816
rect 33367 14776 33416 14804
rect 33367 14773 33379 14776
rect 33321 14767 33379 14773
rect 33410 14764 33416 14776
rect 33468 14804 33474 14816
rect 33778 14804 33784 14816
rect 33468 14776 33784 14804
rect 33468 14764 33474 14776
rect 33778 14764 33784 14776
rect 33836 14804 33842 14816
rect 36262 14804 36268 14816
rect 33836 14776 36268 14804
rect 33836 14764 33842 14776
rect 36262 14764 36268 14776
rect 36320 14764 36326 14816
rect 36446 14764 36452 14816
rect 36504 14804 36510 14816
rect 36832 14804 36860 14844
rect 39022 14832 39028 14844
rect 39080 14872 39086 14884
rect 40313 14875 40371 14881
rect 40313 14872 40325 14875
rect 39080 14844 40325 14872
rect 39080 14832 39086 14844
rect 40313 14841 40325 14844
rect 40359 14841 40371 14875
rect 40313 14835 40371 14841
rect 36504 14776 36860 14804
rect 37737 14807 37795 14813
rect 36504 14764 36510 14776
rect 37737 14773 37749 14807
rect 37783 14804 37795 14807
rect 37826 14804 37832 14816
rect 37783 14776 37832 14804
rect 37783 14773 37795 14776
rect 37737 14767 37795 14773
rect 37826 14764 37832 14776
rect 37884 14764 37890 14816
rect 1104 14714 43884 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 43884 14714
rect 1104 14640 43884 14662
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 17000 14572 17049 14600
rect 17000 14560 17006 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 20070 14600 20076 14612
rect 17037 14563 17095 14569
rect 17144 14572 20076 14600
rect 14461 14535 14519 14541
rect 14461 14501 14473 14535
rect 14507 14532 14519 14535
rect 14507 14504 15792 14532
rect 14507 14501 14519 14504
rect 14461 14495 14519 14501
rect 15396 14473 15424 14504
rect 15764 14476 15792 14504
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 16393 14535 16451 14541
rect 16393 14532 16405 14535
rect 15988 14504 16405 14532
rect 15988 14492 15994 14504
rect 16393 14501 16405 14504
rect 16439 14532 16451 14535
rect 17144 14532 17172 14572
rect 20070 14560 20076 14572
rect 20128 14600 20134 14612
rect 20346 14600 20352 14612
rect 20128 14572 20352 14600
rect 20128 14560 20134 14572
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 20806 14560 20812 14612
rect 20864 14560 20870 14612
rect 22370 14560 22376 14612
rect 22428 14560 22434 14612
rect 24946 14560 24952 14612
rect 25004 14600 25010 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 25004 14572 25053 14600
rect 25004 14560 25010 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25041 14563 25099 14569
rect 27249 14603 27307 14609
rect 27249 14569 27261 14603
rect 27295 14600 27307 14603
rect 27430 14600 27436 14612
rect 27295 14572 27436 14600
rect 27295 14569 27307 14572
rect 27249 14563 27307 14569
rect 27430 14560 27436 14572
rect 27488 14600 27494 14612
rect 27706 14600 27712 14612
rect 27488 14572 27712 14600
rect 27488 14560 27494 14572
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 29178 14560 29184 14612
rect 29236 14560 29242 14612
rect 29730 14560 29736 14612
rect 29788 14560 29794 14612
rect 30006 14560 30012 14612
rect 30064 14600 30070 14612
rect 30064 14572 31984 14600
rect 30064 14560 30070 14572
rect 16439 14504 17172 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 28902 14492 28908 14544
rect 28960 14492 28966 14544
rect 28994 14492 29000 14544
rect 29052 14532 29058 14544
rect 31294 14532 31300 14544
rect 29052 14504 31300 14532
rect 29052 14492 29058 14504
rect 31294 14492 31300 14504
rect 31352 14532 31358 14544
rect 31956 14532 31984 14572
rect 34514 14560 34520 14612
rect 34572 14600 34578 14612
rect 34885 14603 34943 14609
rect 34885 14600 34897 14603
rect 34572 14572 34897 14600
rect 34572 14560 34578 14572
rect 34885 14569 34897 14572
rect 34931 14569 34943 14603
rect 34885 14563 34943 14569
rect 35066 14560 35072 14612
rect 35124 14560 35130 14612
rect 36265 14603 36323 14609
rect 36265 14569 36277 14603
rect 36311 14600 36323 14603
rect 36538 14600 36544 14612
rect 36311 14572 36544 14600
rect 36311 14569 36323 14572
rect 36265 14563 36323 14569
rect 36538 14560 36544 14572
rect 36596 14560 36602 14612
rect 38102 14560 38108 14612
rect 38160 14600 38166 14612
rect 38565 14603 38623 14609
rect 38565 14600 38577 14603
rect 38160 14572 38577 14600
rect 38160 14560 38166 14572
rect 38565 14569 38577 14572
rect 38611 14569 38623 14603
rect 38565 14563 38623 14569
rect 39301 14603 39359 14609
rect 39301 14569 39313 14603
rect 39347 14600 39359 14603
rect 40126 14600 40132 14612
rect 39347 14572 40132 14600
rect 39347 14569 39359 14572
rect 39301 14563 39359 14569
rect 40126 14560 40132 14572
rect 40184 14560 40190 14612
rect 40218 14560 40224 14612
rect 40276 14600 40282 14612
rect 41233 14603 41291 14609
rect 41233 14600 41245 14603
rect 40276 14572 41245 14600
rect 40276 14560 40282 14572
rect 41233 14569 41245 14572
rect 41279 14569 41291 14603
rect 41233 14563 41291 14569
rect 41782 14560 41788 14612
rect 41840 14560 41846 14612
rect 33321 14535 33379 14541
rect 33321 14532 33333 14535
rect 31352 14504 31800 14532
rect 31352 14492 31358 14504
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14433 15439 14467
rect 15381 14427 15439 14433
rect 15470 14424 15476 14476
rect 15528 14424 15534 14476
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 16206 14464 16212 14476
rect 15804 14436 16212 14464
rect 15804 14424 15810 14436
rect 16206 14424 16212 14436
rect 16264 14464 16270 14476
rect 17494 14464 17500 14476
rect 16264 14436 17500 14464
rect 16264 14424 16270 14436
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 17678 14424 17684 14476
rect 17736 14424 17742 14476
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 19208 14436 19441 14464
rect 19208 14424 19214 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 23934 14424 23940 14476
rect 23992 14464 23998 14476
rect 25130 14464 25136 14476
rect 23992 14436 25136 14464
rect 23992 14424 23998 14436
rect 25130 14424 25136 14436
rect 25188 14464 25194 14476
rect 25869 14467 25927 14473
rect 25869 14464 25881 14467
rect 25188 14436 25881 14464
rect 25188 14424 25194 14436
rect 25869 14433 25881 14436
rect 25915 14433 25927 14467
rect 28920 14464 28948 14492
rect 31772 14476 31800 14504
rect 31956 14504 33333 14532
rect 29822 14464 29828 14476
rect 25869 14427 25927 14433
rect 28736 14436 29828 14464
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14396 15347 14399
rect 15838 14396 15844 14408
rect 15335 14368 15844 14396
rect 15335 14365 15347 14368
rect 15289 14359 15347 14365
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14396 17463 14399
rect 18046 14396 18052 14408
rect 17451 14368 18052 14396
rect 17451 14365 17463 14368
rect 17405 14359 17463 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 20254 14396 20260 14408
rect 18739 14368 20260 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 25222 14356 25228 14408
rect 25280 14356 25286 14408
rect 28534 14356 28540 14408
rect 28592 14356 28598 14408
rect 28736 14405 28764 14436
rect 29822 14424 29828 14436
rect 29880 14464 29886 14476
rect 30009 14467 30067 14473
rect 30558 14472 30564 14476
rect 29880 14436 29960 14464
rect 29880 14424 29886 14436
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28721 14359 28779 14365
rect 28810 14356 28816 14408
rect 28868 14356 28874 14408
rect 29932 14405 29960 14436
rect 30009 14433 30021 14467
rect 30055 14464 30067 14467
rect 30392 14464 30564 14472
rect 30055 14444 30564 14464
rect 30055 14436 30420 14444
rect 30055 14433 30067 14436
rect 30009 14427 30067 14433
rect 30558 14424 30564 14444
rect 30616 14424 30622 14476
rect 31662 14424 31668 14476
rect 31720 14424 31726 14476
rect 31754 14424 31760 14476
rect 31812 14424 31818 14476
rect 31956 14473 31984 14504
rect 33321 14501 33333 14504
rect 33367 14501 33379 14535
rect 33321 14495 33379 14501
rect 35894 14492 35900 14544
rect 35952 14532 35958 14544
rect 39117 14535 39175 14541
rect 39117 14532 39129 14535
rect 35952 14504 39129 14532
rect 35952 14492 35958 14504
rect 39117 14501 39129 14504
rect 39163 14501 39175 14535
rect 39117 14495 39175 14501
rect 31941 14467 31999 14473
rect 31941 14433 31953 14467
rect 31987 14433 31999 14467
rect 31941 14427 31999 14433
rect 32582 14424 32588 14476
rect 32640 14464 32646 14476
rect 32640 14436 33180 14464
rect 32640 14424 32646 14436
rect 28905 14399 28963 14405
rect 28905 14365 28917 14399
rect 28951 14365 28963 14399
rect 28905 14359 28963 14365
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 19674 14331 19732 14337
rect 19674 14328 19686 14331
rect 18892 14300 19686 14328
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 18892 14269 18920 14300
rect 19674 14297 19686 14300
rect 19720 14297 19732 14331
rect 19674 14291 19732 14297
rect 26136 14331 26194 14337
rect 26136 14297 26148 14331
rect 26182 14328 26194 14331
rect 26786 14328 26792 14340
rect 26182 14300 26792 14328
rect 26182 14297 26194 14300
rect 26136 14291 26194 14297
rect 26786 14288 26792 14300
rect 26844 14288 26850 14340
rect 28626 14288 28632 14340
rect 28684 14328 28690 14340
rect 28920 14328 28948 14359
rect 30098 14356 30104 14408
rect 30156 14356 30162 14408
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14396 30251 14399
rect 30926 14396 30932 14408
rect 30239 14368 30932 14396
rect 30239 14365 30251 14368
rect 30193 14359 30251 14365
rect 30926 14356 30932 14368
rect 30984 14356 30990 14408
rect 31849 14399 31907 14405
rect 31849 14365 31861 14399
rect 31895 14365 31907 14399
rect 31849 14359 31907 14365
rect 30466 14328 30472 14340
rect 28684 14300 30472 14328
rect 28684 14288 28690 14300
rect 30466 14288 30472 14300
rect 30524 14288 30530 14340
rect 31864 14328 31892 14359
rect 32490 14356 32496 14408
rect 32548 14356 32554 14408
rect 32677 14399 32735 14405
rect 32677 14365 32689 14399
rect 32723 14396 32735 14399
rect 32766 14396 32772 14408
rect 32723 14368 32772 14396
rect 32723 14365 32735 14368
rect 32677 14359 32735 14365
rect 32692 14328 32720 14359
rect 32766 14356 32772 14368
rect 32824 14356 32830 14408
rect 33152 14405 33180 14436
rect 33980 14436 36308 14464
rect 33137 14399 33195 14405
rect 33137 14365 33149 14399
rect 33183 14365 33195 14399
rect 33137 14359 33195 14365
rect 33321 14399 33379 14405
rect 33321 14365 33333 14399
rect 33367 14390 33379 14399
rect 33502 14396 33508 14408
rect 33428 14390 33508 14396
rect 33367 14368 33508 14390
rect 33367 14365 33456 14368
rect 33321 14362 33456 14365
rect 33321 14359 33379 14362
rect 33502 14356 33508 14368
rect 33560 14356 33566 14408
rect 33980 14405 34008 14436
rect 33781 14399 33839 14405
rect 33781 14365 33793 14399
rect 33827 14365 33839 14399
rect 33781 14359 33839 14365
rect 33965 14399 34023 14405
rect 33965 14365 33977 14399
rect 34011 14365 34023 14399
rect 33965 14359 34023 14365
rect 31864 14300 32720 14328
rect 33042 14288 33048 14340
rect 33100 14328 33106 14340
rect 33796 14328 33824 14359
rect 35802 14356 35808 14408
rect 35860 14396 35866 14408
rect 36081 14399 36139 14405
rect 36081 14396 36093 14399
rect 35860 14368 36093 14396
rect 35860 14356 35866 14368
rect 36081 14365 36093 14368
rect 36127 14365 36139 14399
rect 36081 14359 36139 14365
rect 36173 14399 36231 14405
rect 36173 14365 36185 14399
rect 36219 14365 36231 14399
rect 36280 14396 36308 14436
rect 36354 14424 36360 14476
rect 36412 14464 36418 14476
rect 38102 14464 38108 14476
rect 36412 14436 38108 14464
rect 36412 14424 36418 14436
rect 37016 14405 37044 14436
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 38194 14424 38200 14476
rect 38252 14464 38258 14476
rect 39758 14464 39764 14476
rect 38252 14436 39764 14464
rect 38252 14424 38258 14436
rect 39758 14424 39764 14436
rect 39816 14424 39822 14476
rect 39850 14424 39856 14476
rect 39908 14464 39914 14476
rect 40405 14467 40463 14473
rect 40405 14464 40417 14467
rect 39908 14436 40417 14464
rect 39908 14424 39914 14436
rect 40405 14433 40417 14436
rect 40451 14433 40463 14467
rect 40405 14427 40463 14433
rect 37001 14399 37059 14405
rect 36280 14368 36952 14396
rect 36173 14359 36231 14365
rect 33100 14300 33824 14328
rect 33100 14288 33106 14300
rect 33870 14288 33876 14340
rect 33928 14288 33934 14340
rect 35253 14331 35311 14337
rect 35253 14297 35265 14331
rect 35299 14328 35311 14331
rect 35342 14328 35348 14340
rect 35299 14300 35348 14328
rect 35299 14297 35311 14300
rect 35253 14291 35311 14297
rect 35342 14288 35348 14300
rect 35400 14288 35406 14340
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14884 14232 14933 14260
rect 14884 14220 14890 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 18877 14263 18935 14269
rect 18877 14229 18889 14263
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 24394 14220 24400 14272
rect 24452 14260 24458 14272
rect 25222 14260 25228 14272
rect 24452 14232 25228 14260
rect 24452 14220 24458 14232
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 30742 14220 30748 14272
rect 30800 14220 30806 14272
rect 31478 14220 31484 14272
rect 31536 14220 31542 14272
rect 31570 14220 31576 14272
rect 31628 14260 31634 14272
rect 32493 14263 32551 14269
rect 32493 14260 32505 14263
rect 31628 14232 32505 14260
rect 31628 14220 31634 14232
rect 32493 14229 32505 14232
rect 32539 14229 32551 14263
rect 32493 14223 32551 14229
rect 33778 14220 33784 14272
rect 33836 14260 33842 14272
rect 35043 14263 35101 14269
rect 35043 14260 35055 14263
rect 33836 14232 35055 14260
rect 33836 14220 33842 14232
rect 35043 14229 35055 14232
rect 35089 14260 35101 14263
rect 35158 14260 35164 14272
rect 35089 14232 35164 14260
rect 35089 14229 35101 14232
rect 35043 14223 35101 14229
rect 35158 14220 35164 14232
rect 35216 14220 35222 14272
rect 35360 14260 35388 14288
rect 35802 14260 35808 14272
rect 35360 14232 35808 14260
rect 35802 14220 35808 14232
rect 35860 14220 35866 14272
rect 36096 14260 36124 14359
rect 36188 14328 36216 14359
rect 36814 14328 36820 14340
rect 36188 14300 36820 14328
rect 36814 14288 36820 14300
rect 36872 14288 36878 14340
rect 36170 14260 36176 14272
rect 36096 14232 36176 14260
rect 36170 14220 36176 14232
rect 36228 14220 36234 14272
rect 36924 14260 36952 14368
rect 37001 14365 37013 14399
rect 37047 14365 37059 14399
rect 37001 14359 37059 14365
rect 37182 14356 37188 14408
rect 37240 14396 37246 14408
rect 37550 14396 37556 14408
rect 37240 14368 37556 14396
rect 37240 14356 37246 14368
rect 37550 14356 37556 14368
rect 37608 14356 37614 14408
rect 37734 14356 37740 14408
rect 37792 14356 37798 14408
rect 38473 14399 38531 14405
rect 38473 14365 38485 14399
rect 38519 14365 38531 14399
rect 38473 14359 38531 14365
rect 38657 14399 38715 14405
rect 38657 14365 38669 14399
rect 38703 14396 38715 14399
rect 39114 14396 39120 14408
rect 38703 14368 39120 14396
rect 38703 14365 38715 14368
rect 38657 14359 38715 14365
rect 38286 14328 38292 14340
rect 37292 14300 38292 14328
rect 37292 14260 37320 14300
rect 38286 14288 38292 14300
rect 38344 14288 38350 14340
rect 38488 14328 38516 14359
rect 39114 14356 39120 14368
rect 39172 14356 39178 14408
rect 39574 14396 39580 14408
rect 39500 14368 39580 14396
rect 39500 14337 39528 14368
rect 39574 14356 39580 14368
rect 39632 14396 39638 14408
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 39632 14368 40049 14396
rect 39632 14356 39638 14368
rect 40037 14365 40049 14368
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 40126 14356 40132 14408
rect 40184 14396 40190 14408
rect 40497 14399 40555 14405
rect 40497 14396 40509 14399
rect 40184 14368 40509 14396
rect 40184 14356 40190 14368
rect 40497 14365 40509 14368
rect 40543 14365 40555 14399
rect 40497 14359 40555 14365
rect 43346 14356 43352 14408
rect 43404 14356 43410 14408
rect 39485 14331 39543 14337
rect 39485 14328 39497 14331
rect 38488 14300 39497 14328
rect 39485 14297 39497 14300
rect 39531 14297 39543 14331
rect 39485 14291 39543 14297
rect 40310 14288 40316 14340
rect 40368 14328 40374 14340
rect 40586 14328 40592 14340
rect 40368 14300 40592 14328
rect 40368 14288 40374 14300
rect 40586 14288 40592 14300
rect 40644 14328 40650 14340
rect 42337 14331 42395 14337
rect 42337 14328 42349 14331
rect 40644 14300 42349 14328
rect 40644 14288 40650 14300
rect 42337 14297 42349 14300
rect 42383 14297 42395 14331
rect 42337 14291 42395 14297
rect 43070 14288 43076 14340
rect 43128 14288 43134 14340
rect 36924 14232 37320 14260
rect 37918 14220 37924 14272
rect 37976 14260 37982 14272
rect 38562 14260 38568 14272
rect 37976 14232 38568 14260
rect 37976 14220 37982 14232
rect 38562 14220 38568 14232
rect 38620 14220 38626 14272
rect 39285 14263 39343 14269
rect 39285 14229 39297 14263
rect 39331 14260 39343 14263
rect 40494 14260 40500 14272
rect 39331 14232 40500 14260
rect 39331 14229 39343 14232
rect 39285 14223 39343 14229
rect 40494 14220 40500 14232
rect 40552 14220 40558 14272
rect 1104 14170 43884 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 43884 14170
rect 1104 14096 43884 14118
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 15838 14056 15844 14068
rect 15611 14028 15844 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16206 14016 16212 14068
rect 16264 14016 16270 14068
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 17865 14059 17923 14065
rect 17865 14056 17877 14059
rect 17552 14028 17877 14056
rect 17552 14016 17558 14028
rect 17865 14025 17877 14028
rect 17911 14025 17923 14059
rect 17865 14019 17923 14025
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 19978 14056 19984 14068
rect 19843 14028 19984 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20625 14059 20683 14065
rect 20625 14025 20637 14059
rect 20671 14056 20683 14059
rect 20806 14056 20812 14068
rect 20671 14028 20812 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 22833 14059 22891 14065
rect 22833 14025 22845 14059
rect 22879 14056 22891 14059
rect 23750 14056 23756 14068
rect 22879 14028 23756 14056
rect 22879 14025 22891 14028
rect 22833 14019 22891 14025
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 24857 14059 24915 14065
rect 24857 14025 24869 14059
rect 24903 14025 24915 14059
rect 24857 14019 24915 14025
rect 15102 13988 15108 14000
rect 14200 13960 15108 13988
rect 14200 13929 14228 13960
rect 15102 13948 15108 13960
rect 15160 13948 15166 14000
rect 19150 13988 19156 14000
rect 18432 13960 19156 13988
rect 14458 13929 14464 13932
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14452 13883 14464 13929
rect 14458 13880 14464 13883
rect 14516 13880 14522 13932
rect 18432 13929 18460 13960
rect 19150 13948 19156 13960
rect 19208 13948 19214 14000
rect 20162 13948 20168 14000
rect 20220 13988 20226 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 20220 13960 20729 13988
rect 20220 13948 20226 13960
rect 20717 13957 20729 13960
rect 20763 13957 20775 13991
rect 20717 13951 20775 13957
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22462 13988 22468 14000
rect 22244 13960 22468 13988
rect 22244 13948 22250 13960
rect 22462 13948 22468 13960
rect 22520 13988 22526 14000
rect 22925 13991 22983 13997
rect 22925 13988 22937 13991
rect 22520 13960 22937 13988
rect 22520 13948 22526 13960
rect 22925 13957 22937 13960
rect 22971 13957 22983 13991
rect 22925 13951 22983 13957
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18684 13923 18742 13929
rect 18684 13889 18696 13923
rect 18730 13920 18742 13923
rect 19518 13920 19524 13932
rect 18730 13892 19524 13920
rect 18730 13889 18742 13892
rect 18684 13883 18742 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13920 24271 13923
rect 24872 13920 24900 14019
rect 25222 14016 25228 14068
rect 25280 14016 25286 14068
rect 25317 14059 25375 14065
rect 25317 14025 25329 14059
rect 25363 14025 25375 14059
rect 25317 14019 25375 14025
rect 27157 14059 27215 14065
rect 27157 14025 27169 14059
rect 27203 14056 27215 14059
rect 27338 14056 27344 14068
rect 27203 14028 27344 14056
rect 27203 14025 27215 14028
rect 27157 14019 27215 14025
rect 25332 13988 25360 14019
rect 27338 14016 27344 14028
rect 27396 14016 27402 14068
rect 30006 14056 30012 14068
rect 27448 14028 30012 14056
rect 27448 13988 27476 14028
rect 30006 14016 30012 14028
rect 30064 14016 30070 14068
rect 30098 14016 30104 14068
rect 30156 14016 30162 14068
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 31478 14056 31484 14068
rect 30524 14028 31484 14056
rect 30524 14016 30530 14028
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 31570 14016 31576 14068
rect 31628 14016 31634 14068
rect 34146 14056 34152 14068
rect 31680 14028 34152 14056
rect 25332 13960 27476 13988
rect 27522 13948 27528 14000
rect 27580 13988 27586 14000
rect 28270 13991 28328 13997
rect 28270 13988 28282 13991
rect 27580 13960 28282 13988
rect 27580 13948 27586 13960
rect 28270 13957 28282 13960
rect 28316 13957 28328 13991
rect 29638 13988 29644 14000
rect 28270 13951 28328 13957
rect 29380 13960 29644 13988
rect 24259 13892 24900 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 26418 13880 26424 13932
rect 26476 13880 26482 13932
rect 26605 13923 26663 13929
rect 26605 13889 26617 13923
rect 26651 13920 26663 13923
rect 28994 13920 29000 13932
rect 26651 13892 29000 13920
rect 26651 13889 26663 13892
rect 26605 13883 26663 13889
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 29086 13880 29092 13932
rect 29144 13880 29150 13932
rect 29270 13880 29276 13932
rect 29328 13880 29334 13932
rect 29380 13929 29408 13960
rect 29638 13948 29644 13960
rect 29696 13948 29702 14000
rect 29730 13948 29736 14000
rect 29788 13988 29794 14000
rect 31680 13988 31708 14028
rect 34146 14016 34152 14028
rect 34204 14016 34210 14068
rect 34422 14016 34428 14068
rect 34480 14056 34486 14068
rect 34701 14059 34759 14065
rect 34701 14056 34713 14059
rect 34480 14028 34713 14056
rect 34480 14016 34486 14028
rect 34701 14025 34713 14028
rect 34747 14025 34759 14059
rect 36078 14056 36084 14068
rect 34701 14019 34759 14025
rect 35360 14028 36084 14056
rect 29788 13960 31708 13988
rect 29788 13948 29794 13960
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29365 13883 29423 13889
rect 29457 13923 29515 13929
rect 29457 13889 29469 13923
rect 29503 13920 29515 13923
rect 29503 13892 29776 13920
rect 29503 13889 29515 13892
rect 29457 13883 29515 13889
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 23017 13855 23075 13861
rect 23017 13821 23029 13855
rect 23063 13821 23075 13855
rect 24854 13852 24860 13864
rect 23017 13815 23075 13821
rect 24412 13824 24860 13852
rect 20162 13744 20168 13796
rect 20220 13784 20226 13796
rect 20916 13784 20944 13815
rect 22370 13784 22376 13796
rect 20220 13756 22376 13784
rect 20220 13744 20226 13756
rect 22370 13744 22376 13756
rect 22428 13784 22434 13796
rect 23032 13784 23060 13815
rect 24412 13793 24440 13824
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25501 13855 25559 13861
rect 25501 13821 25513 13855
rect 25547 13821 25559 13855
rect 25501 13815 25559 13821
rect 28537 13855 28595 13861
rect 28537 13821 28549 13855
rect 28583 13852 28595 13855
rect 29178 13852 29184 13864
rect 28583 13824 29184 13852
rect 28583 13821 28595 13824
rect 28537 13815 28595 13821
rect 22428 13756 23060 13784
rect 24397 13787 24455 13793
rect 22428 13744 22434 13756
rect 24397 13753 24409 13787
rect 24443 13753 24455 13787
rect 25516 13784 25544 13815
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 29748 13852 29776 13892
rect 30282 13880 30288 13932
rect 30340 13880 30346 13932
rect 30374 13880 30380 13932
rect 30432 13920 30438 13932
rect 31496 13929 31524 13960
rect 31754 13948 31760 14000
rect 31812 13988 31818 14000
rect 33042 13988 33048 14000
rect 31812 13960 33048 13988
rect 31812 13948 31818 13960
rect 33042 13948 33048 13960
rect 33100 13988 33106 14000
rect 33229 13991 33287 13997
rect 33229 13988 33241 13991
rect 33100 13960 33241 13988
rect 33100 13948 33106 13960
rect 33229 13957 33241 13960
rect 33275 13957 33287 13991
rect 33229 13951 33287 13957
rect 33410 13948 33416 14000
rect 33468 13948 33474 14000
rect 33502 13948 33508 14000
rect 33560 13988 33566 14000
rect 35360 13988 35388 14028
rect 36078 14016 36084 14028
rect 36136 14056 36142 14068
rect 37090 14056 37096 14068
rect 36136 14028 37096 14056
rect 36136 14016 36142 14028
rect 37090 14016 37096 14028
rect 37148 14016 37154 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37645 14059 37703 14065
rect 37645 14056 37657 14059
rect 37424 14028 37657 14056
rect 37424 14016 37430 14028
rect 37645 14025 37657 14028
rect 37691 14025 37703 14059
rect 37645 14019 37703 14025
rect 38286 14016 38292 14068
rect 38344 14016 38350 14068
rect 41141 14059 41199 14065
rect 41141 14025 41153 14059
rect 41187 14056 41199 14059
rect 41230 14056 41236 14068
rect 41187 14028 41236 14056
rect 41187 14025 41199 14028
rect 41141 14019 41199 14025
rect 41230 14016 41236 14028
rect 41288 14016 41294 14068
rect 42613 14059 42671 14065
rect 42613 14056 42625 14059
rect 41386 14028 42625 14056
rect 33560 13960 35388 13988
rect 33560 13948 33566 13960
rect 30561 13923 30619 13929
rect 30561 13920 30573 13923
rect 30432 13892 30573 13920
rect 30432 13880 30438 13892
rect 30561 13889 30573 13892
rect 30607 13920 30619 13923
rect 31481 13923 31539 13929
rect 30607 13892 31432 13920
rect 30607 13889 30619 13892
rect 30561 13883 30619 13889
rect 30742 13852 30748 13864
rect 29748 13824 30748 13852
rect 26234 13784 26240 13796
rect 25516 13756 26240 13784
rect 24397 13747 24455 13753
rect 26234 13744 26240 13756
rect 26292 13744 26298 13796
rect 29748 13784 29776 13824
rect 30742 13812 30748 13824
rect 30800 13812 30806 13864
rect 28920 13756 29776 13784
rect 31404 13784 31432 13892
rect 31481 13889 31493 13923
rect 31527 13889 31539 13923
rect 31481 13883 31539 13889
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 33612 13929 33640 13960
rect 32493 13923 32551 13929
rect 32493 13920 32505 13923
rect 31720 13892 32505 13920
rect 31720 13880 31726 13892
rect 32493 13889 32505 13892
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 33597 13923 33655 13929
rect 33597 13889 33609 13923
rect 33643 13889 33655 13923
rect 33597 13883 33655 13889
rect 34882 13880 34888 13932
rect 34940 13880 34946 13932
rect 35360 13929 35388 13960
rect 35618 13948 35624 14000
rect 35676 13988 35682 14000
rect 38654 13988 38660 14000
rect 35676 13960 38660 13988
rect 35676 13948 35682 13960
rect 35526 13929 35532 13932
rect 35345 13923 35403 13929
rect 35345 13889 35357 13923
rect 35391 13889 35403 13923
rect 35345 13883 35403 13889
rect 35523 13883 35532 13929
rect 35584 13920 35590 13932
rect 35584 13892 35756 13920
rect 35526 13880 35532 13883
rect 35584 13880 35590 13892
rect 32677 13855 32735 13861
rect 32677 13821 32689 13855
rect 32723 13852 32735 13855
rect 32766 13852 32772 13864
rect 32723 13824 32772 13852
rect 32723 13821 32735 13824
rect 32677 13815 32735 13821
rect 32766 13812 32772 13824
rect 32824 13812 32830 13864
rect 34698 13812 34704 13864
rect 34756 13852 34762 13864
rect 35437 13855 35495 13861
rect 35437 13852 35449 13855
rect 34756 13824 35449 13852
rect 34756 13812 34762 13824
rect 35437 13821 35449 13824
rect 35483 13821 35495 13855
rect 35437 13815 35495 13821
rect 34716 13784 34744 13812
rect 31404 13756 34744 13784
rect 22462 13676 22468 13728
rect 22520 13676 22526 13728
rect 26510 13676 26516 13728
rect 26568 13676 26574 13728
rect 27614 13676 27620 13728
rect 27672 13716 27678 13728
rect 28920 13716 28948 13756
rect 34882 13744 34888 13796
rect 34940 13784 34946 13796
rect 35618 13784 35624 13796
rect 34940 13756 35624 13784
rect 34940 13744 34946 13756
rect 35618 13744 35624 13756
rect 35676 13744 35682 13796
rect 35728 13784 35756 13892
rect 36354 13880 36360 13932
rect 36412 13924 36418 13932
rect 36449 13924 36507 13929
rect 36412 13923 36507 13924
rect 36412 13896 36461 13923
rect 36412 13880 36418 13896
rect 36449 13889 36461 13896
rect 36495 13889 36507 13923
rect 36449 13883 36507 13889
rect 36633 13923 36691 13929
rect 36633 13889 36645 13923
rect 36679 13920 36691 13923
rect 36679 13892 37044 13920
rect 36679 13889 36691 13892
rect 36633 13883 36691 13889
rect 36541 13855 36599 13861
rect 36541 13821 36553 13855
rect 36587 13852 36599 13855
rect 36722 13852 36728 13864
rect 36587 13824 36728 13852
rect 36587 13821 36599 13824
rect 36541 13815 36599 13821
rect 36722 13812 36728 13824
rect 36780 13812 36786 13864
rect 37016 13784 37044 13892
rect 37458 13880 37464 13932
rect 37516 13880 37522 13932
rect 38212 13929 38240 13960
rect 38654 13948 38660 13960
rect 38712 13948 38718 14000
rect 38933 13991 38991 13997
rect 38933 13988 38945 13991
rect 38764 13960 38945 13988
rect 38197 13923 38255 13929
rect 38197 13889 38209 13923
rect 38243 13889 38255 13923
rect 38197 13883 38255 13889
rect 38381 13923 38439 13929
rect 38381 13889 38393 13923
rect 38427 13920 38439 13923
rect 38764 13920 38792 13960
rect 38933 13957 38945 13960
rect 38979 13957 38991 13991
rect 38933 13951 38991 13957
rect 39114 13948 39120 14000
rect 39172 13988 39178 14000
rect 41386 13988 41414 14028
rect 42613 14025 42625 14028
rect 42659 14025 42671 14059
rect 42613 14019 42671 14025
rect 42981 14059 43039 14065
rect 42981 14025 42993 14059
rect 43027 14056 43039 14059
rect 43070 14056 43076 14068
rect 43027 14028 43076 14056
rect 43027 14025 43039 14028
rect 42981 14019 43039 14025
rect 43070 14016 43076 14028
rect 43128 14016 43134 14068
rect 39172 13960 41414 13988
rect 39172 13948 39178 13960
rect 41874 13948 41880 14000
rect 41932 13988 41938 14000
rect 41969 13991 42027 13997
rect 41969 13988 41981 13991
rect 41932 13960 41981 13988
rect 41932 13948 41938 13960
rect 41969 13957 41981 13960
rect 42015 13957 42027 13991
rect 41969 13951 42027 13957
rect 38427 13892 38792 13920
rect 38841 13923 38899 13929
rect 38427 13889 38439 13892
rect 38381 13883 38439 13889
rect 38841 13889 38853 13923
rect 38887 13889 38899 13923
rect 38841 13883 38899 13889
rect 37734 13812 37740 13864
rect 37792 13852 37798 13864
rect 38396 13852 38424 13883
rect 37792 13824 38424 13852
rect 37792 13812 37798 13824
rect 38562 13812 38568 13864
rect 38620 13852 38626 13864
rect 38856 13852 38884 13883
rect 39022 13880 39028 13932
rect 39080 13880 39086 13932
rect 39574 13880 39580 13932
rect 39632 13880 39638 13932
rect 39758 13880 39764 13932
rect 39816 13920 39822 13932
rect 39945 13923 40003 13929
rect 39945 13920 39957 13923
rect 39816 13892 39957 13920
rect 39816 13880 39822 13892
rect 39945 13889 39957 13892
rect 39991 13889 40003 13923
rect 39945 13883 40003 13889
rect 40313 13923 40371 13929
rect 40313 13889 40325 13923
rect 40359 13920 40371 13923
rect 40494 13920 40500 13932
rect 40359 13892 40500 13920
rect 40359 13889 40371 13892
rect 40313 13883 40371 13889
rect 40494 13880 40500 13892
rect 40552 13880 40558 13932
rect 39592 13852 39620 13880
rect 38620 13824 39620 13852
rect 38620 13812 38626 13824
rect 41046 13812 41052 13864
rect 41104 13852 41110 13864
rect 41233 13855 41291 13861
rect 41233 13852 41245 13855
rect 41104 13824 41245 13852
rect 41104 13812 41110 13824
rect 41233 13821 41245 13824
rect 41279 13821 41291 13855
rect 41233 13815 41291 13821
rect 41417 13855 41475 13861
rect 41417 13821 41429 13855
rect 41463 13852 41475 13855
rect 42886 13852 42892 13864
rect 41463 13824 42892 13852
rect 41463 13821 41475 13824
rect 41417 13815 41475 13821
rect 42886 13812 42892 13824
rect 42944 13812 42950 13864
rect 43070 13812 43076 13864
rect 43128 13812 43134 13864
rect 43257 13855 43315 13861
rect 43257 13821 43269 13855
rect 43303 13821 43315 13855
rect 43257 13815 43315 13821
rect 38746 13784 38752 13796
rect 35728 13756 38752 13784
rect 38746 13744 38752 13756
rect 38804 13744 38810 13796
rect 40034 13744 40040 13796
rect 40092 13784 40098 13796
rect 40773 13787 40831 13793
rect 40773 13784 40785 13787
rect 40092 13756 40785 13784
rect 40092 13744 40098 13756
rect 40773 13753 40785 13756
rect 40819 13753 40831 13787
rect 40773 13747 40831 13753
rect 41138 13744 41144 13796
rect 41196 13784 41202 13796
rect 43162 13784 43168 13796
rect 41196 13756 43168 13784
rect 41196 13744 41202 13756
rect 43162 13744 43168 13756
rect 43220 13784 43226 13796
rect 43272 13784 43300 13815
rect 43220 13756 43300 13784
rect 43220 13744 43226 13756
rect 27672 13688 28948 13716
rect 27672 13676 27678 13688
rect 29178 13676 29184 13728
rect 29236 13716 29242 13728
rect 29454 13716 29460 13728
rect 29236 13688 29460 13716
rect 29236 13676 29242 13688
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 29546 13676 29552 13728
rect 29604 13716 29610 13728
rect 29641 13719 29699 13725
rect 29641 13716 29653 13719
rect 29604 13688 29653 13716
rect 29604 13676 29610 13688
rect 29641 13685 29653 13688
rect 29687 13685 29699 13719
rect 29641 13679 29699 13685
rect 31757 13719 31815 13725
rect 31757 13685 31769 13719
rect 31803 13716 31815 13719
rect 32214 13716 32220 13728
rect 31803 13688 32220 13716
rect 31803 13685 31815 13688
rect 31757 13679 31815 13685
rect 32214 13676 32220 13688
rect 32272 13676 32278 13728
rect 32309 13719 32367 13725
rect 32309 13685 32321 13719
rect 32355 13716 32367 13719
rect 32490 13716 32496 13728
rect 32355 13688 32496 13716
rect 32355 13685 32367 13688
rect 32309 13679 32367 13685
rect 32490 13676 32496 13688
rect 32548 13676 32554 13728
rect 33134 13676 33140 13728
rect 33192 13716 33198 13728
rect 34698 13716 34704 13728
rect 33192 13688 34704 13716
rect 33192 13676 33198 13688
rect 34698 13676 34704 13688
rect 34756 13716 34762 13728
rect 35434 13716 35440 13728
rect 34756 13688 35440 13716
rect 34756 13676 34762 13688
rect 35434 13676 35440 13688
rect 35492 13676 35498 13728
rect 1104 13626 43884 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 43884 13626
rect 1104 13552 43884 13574
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14516 13484 14657 13512
rect 14516 13472 14522 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15933 13515 15991 13521
rect 15933 13512 15945 13515
rect 15528 13484 15945 13512
rect 15528 13472 15534 13484
rect 15933 13481 15945 13484
rect 15979 13481 15991 13515
rect 15933 13475 15991 13481
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19518 13512 19524 13524
rect 19475 13484 19524 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 23661 13515 23719 13521
rect 23661 13481 23673 13515
rect 23707 13512 23719 13515
rect 23750 13512 23756 13524
rect 23707 13484 23756 13512
rect 23707 13481 23719 13484
rect 23661 13475 23719 13481
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 25222 13472 25228 13524
rect 25280 13512 25286 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25280 13484 25973 13512
rect 25280 13472 25286 13484
rect 25961 13481 25973 13484
rect 26007 13481 26019 13515
rect 25961 13475 26019 13481
rect 26786 13472 26792 13524
rect 26844 13472 26850 13524
rect 29086 13472 29092 13524
rect 29144 13512 29150 13524
rect 29825 13515 29883 13521
rect 29825 13512 29837 13515
rect 29144 13484 29837 13512
rect 29144 13472 29150 13484
rect 29825 13481 29837 13484
rect 29871 13481 29883 13515
rect 29825 13475 29883 13481
rect 31757 13515 31815 13521
rect 31757 13481 31769 13515
rect 31803 13512 31815 13515
rect 31846 13512 31852 13524
rect 31803 13484 31852 13512
rect 31803 13481 31815 13484
rect 31757 13475 31815 13481
rect 31846 13472 31852 13484
rect 31904 13472 31910 13524
rect 33505 13515 33563 13521
rect 33505 13481 33517 13515
rect 33551 13512 33563 13515
rect 34790 13512 34796 13524
rect 33551 13484 34796 13512
rect 33551 13481 33563 13484
rect 33505 13475 33563 13481
rect 34790 13472 34796 13484
rect 34848 13472 34854 13524
rect 35710 13472 35716 13524
rect 35768 13472 35774 13524
rect 37458 13472 37464 13524
rect 37516 13472 37522 13524
rect 38654 13472 38660 13524
rect 38712 13472 38718 13524
rect 43070 13472 43076 13524
rect 43128 13512 43134 13524
rect 43257 13515 43315 13521
rect 43257 13512 43269 13515
rect 43128 13484 43269 13512
rect 43128 13472 43134 13484
rect 43257 13481 43269 13484
rect 43303 13481 43315 13515
rect 43257 13475 43315 13481
rect 19334 13404 19340 13456
rect 19392 13444 19398 13456
rect 20533 13447 20591 13453
rect 20533 13444 20545 13447
rect 19392 13416 20545 13444
rect 19392 13404 19398 13416
rect 20533 13413 20545 13416
rect 20579 13444 20591 13447
rect 29181 13447 29239 13453
rect 20579 13416 21680 13444
rect 20579 13413 20591 13416
rect 20533 13407 20591 13413
rect 21652 13385 21680 13416
rect 29181 13413 29193 13447
rect 29227 13444 29239 13447
rect 29270 13444 29276 13456
rect 29227 13416 29276 13444
rect 29227 13413 29239 13416
rect 29181 13407 29239 13413
rect 29270 13404 29276 13416
rect 29328 13404 29334 13456
rect 33134 13444 33140 13456
rect 32048 13416 33140 13444
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13345 21695 13379
rect 21637 13339 21695 13345
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 26973 13379 27031 13385
rect 26973 13376 26985 13379
rect 26568 13348 26985 13376
rect 26568 13336 26574 13348
rect 26973 13345 26985 13348
rect 27019 13345 27031 13379
rect 26973 13339 27031 13345
rect 27430 13336 27436 13388
rect 27488 13336 27494 13388
rect 29730 13376 29736 13388
rect 28828 13348 29736 13376
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19484 13280 19625 13308
rect 19484 13268 19490 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 21591 13280 21864 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 21453 13243 21511 13249
rect 21453 13209 21465 13243
rect 21499 13240 21511 13243
rect 21836 13240 21864 13280
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22281 13311 22339 13317
rect 22281 13308 22293 13311
rect 22060 13280 22293 13308
rect 22060 13268 22066 13280
rect 22281 13277 22293 13280
rect 22327 13308 22339 13311
rect 23934 13308 23940 13320
rect 22327 13280 23940 13308
rect 22327 13277 22339 13280
rect 22281 13271 22339 13277
rect 23934 13268 23940 13280
rect 23992 13308 23998 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 23992 13280 24593 13308
rect 23992 13268 23998 13280
rect 24581 13277 24593 13280
rect 24627 13308 24639 13311
rect 25130 13308 25136 13320
rect 24627 13280 25136 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 27065 13311 27123 13317
rect 27065 13277 27077 13311
rect 27111 13308 27123 13311
rect 28828 13308 28856 13348
rect 29730 13336 29736 13348
rect 29788 13336 29794 13388
rect 30834 13376 30840 13388
rect 29932 13348 30840 13376
rect 27111 13280 28856 13308
rect 27111 13277 27123 13280
rect 27065 13271 27123 13277
rect 28902 13268 28908 13320
rect 28960 13268 28966 13320
rect 28997 13311 29055 13317
rect 28997 13277 29009 13311
rect 29043 13308 29055 13311
rect 29932 13308 29960 13348
rect 30834 13336 30840 13348
rect 30892 13336 30898 13388
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13376 30987 13379
rect 31662 13376 31668 13388
rect 30975 13348 31668 13376
rect 30975 13345 30987 13348
rect 30929 13339 30987 13345
rect 31662 13336 31668 13348
rect 31720 13376 31726 13388
rect 32048 13385 32076 13416
rect 33134 13404 33140 13416
rect 33192 13404 33198 13456
rect 33226 13404 33232 13456
rect 33284 13444 33290 13456
rect 33597 13447 33655 13453
rect 33597 13444 33609 13447
rect 33284 13416 33609 13444
rect 33284 13404 33290 13416
rect 33597 13413 33609 13416
rect 33643 13413 33655 13447
rect 33597 13407 33655 13413
rect 34238 13404 34244 13456
rect 34296 13444 34302 13456
rect 34977 13447 35035 13453
rect 34977 13444 34989 13447
rect 34296 13416 34989 13444
rect 34296 13404 34302 13416
rect 34977 13413 34989 13416
rect 35023 13413 35035 13447
rect 34977 13407 35035 13413
rect 35342 13404 35348 13456
rect 35400 13444 35406 13456
rect 35989 13447 36047 13453
rect 35989 13444 36001 13447
rect 35400 13416 36001 13444
rect 35400 13404 35406 13416
rect 35989 13413 36001 13416
rect 36035 13444 36047 13447
rect 36446 13444 36452 13456
rect 36035 13416 36452 13444
rect 36035 13413 36047 13416
rect 35989 13407 36047 13413
rect 36446 13404 36452 13416
rect 36504 13404 36510 13456
rect 40034 13404 40040 13456
rect 40092 13404 40098 13456
rect 31941 13379 31999 13385
rect 31941 13376 31953 13379
rect 31720 13348 31953 13376
rect 31720 13336 31726 13348
rect 31941 13345 31953 13348
rect 31987 13345 31999 13379
rect 31941 13339 31999 13345
rect 32033 13379 32091 13385
rect 32033 13345 32045 13379
rect 32079 13345 32091 13379
rect 33413 13379 33471 13385
rect 33413 13376 33425 13379
rect 32033 13339 32091 13345
rect 32140 13348 33425 13376
rect 29043 13280 29960 13308
rect 29043 13277 29055 13280
rect 28997 13271 29055 13277
rect 30006 13268 30012 13320
rect 30064 13268 30070 13320
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13308 30343 13311
rect 30374 13308 30380 13320
rect 30331 13280 30380 13308
rect 30331 13277 30343 13280
rect 30285 13271 30343 13277
rect 30374 13268 30380 13280
rect 30432 13268 30438 13320
rect 31018 13268 31024 13320
rect 31076 13268 31082 13320
rect 31113 13311 31171 13317
rect 31113 13277 31125 13311
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 31205 13311 31263 13317
rect 31205 13277 31217 13311
rect 31251 13308 31263 13311
rect 31846 13308 31852 13320
rect 31251 13280 31852 13308
rect 31251 13277 31263 13280
rect 31205 13271 31263 13277
rect 22186 13240 22192 13252
rect 21499 13212 21772 13240
rect 21836 13212 22192 13240
rect 21499 13209 21511 13212
rect 21453 13203 21511 13209
rect 21085 13175 21143 13181
rect 21085 13141 21097 13175
rect 21131 13172 21143 13175
rect 21266 13172 21272 13184
rect 21131 13144 21272 13172
rect 21131 13141 21143 13144
rect 21085 13135 21143 13141
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 21744 13172 21772 13212
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 22548 13243 22606 13249
rect 22548 13209 22560 13243
rect 22594 13240 22606 13243
rect 22646 13240 22652 13252
rect 22594 13212 22652 13240
rect 22594 13209 22606 13212
rect 22548 13203 22606 13209
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 24854 13249 24860 13252
rect 24848 13240 24860 13249
rect 24815 13212 24860 13240
rect 24848 13203 24860 13212
rect 24854 13200 24860 13203
rect 24912 13200 24918 13252
rect 27341 13243 27399 13249
rect 27341 13209 27353 13243
rect 27387 13240 27399 13243
rect 27614 13240 27620 13252
rect 27387 13212 27620 13240
rect 27387 13209 27399 13212
rect 27341 13203 27399 13209
rect 27614 13200 27620 13212
rect 27672 13240 27678 13252
rect 27893 13243 27951 13249
rect 27893 13240 27905 13243
rect 27672 13212 27905 13240
rect 27672 13200 27678 13212
rect 27893 13209 27905 13212
rect 27939 13209 27951 13243
rect 31128 13240 31156 13271
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 32140 13317 32168 13348
rect 33413 13345 33425 13348
rect 33459 13376 33471 13379
rect 34422 13376 34428 13388
rect 33459 13348 34428 13376
rect 33459 13345 33471 13348
rect 33413 13339 33471 13345
rect 34422 13336 34428 13348
rect 34480 13336 34486 13388
rect 35526 13376 35532 13388
rect 35084 13348 35532 13376
rect 32125 13311 32183 13317
rect 32125 13277 32137 13311
rect 32171 13277 32183 13311
rect 32125 13271 32183 13277
rect 27893 13203 27951 13209
rect 30208 13212 31156 13240
rect 23290 13172 23296 13184
rect 21744 13144 23296 13172
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 29914 13132 29920 13184
rect 29972 13172 29978 13184
rect 30208 13181 30236 13212
rect 31478 13200 31484 13252
rect 31536 13240 31542 13252
rect 32140 13240 32168 13271
rect 32214 13268 32220 13320
rect 32272 13268 32278 13320
rect 33689 13311 33747 13317
rect 33689 13308 33701 13311
rect 32876 13280 33701 13308
rect 31536 13212 32168 13240
rect 31536 13200 31542 13212
rect 30193 13175 30251 13181
rect 30193 13172 30205 13175
rect 29972 13144 30205 13172
rect 29972 13132 29978 13144
rect 30193 13141 30205 13144
rect 30239 13141 30251 13175
rect 30193 13135 30251 13141
rect 30742 13132 30748 13184
rect 30800 13132 30806 13184
rect 31018 13132 31024 13184
rect 31076 13172 31082 13184
rect 32876 13172 32904 13280
rect 33689 13277 33701 13280
rect 33735 13308 33747 13311
rect 33778 13308 33784 13320
rect 33735 13280 33784 13308
rect 33735 13277 33747 13280
rect 33689 13271 33747 13277
rect 33778 13268 33784 13280
rect 33836 13268 33842 13320
rect 33873 13311 33931 13317
rect 33873 13277 33885 13311
rect 33919 13308 33931 13311
rect 35084 13308 35112 13348
rect 35526 13336 35532 13348
rect 35584 13336 35590 13388
rect 36081 13379 36139 13385
rect 36081 13345 36093 13379
rect 36127 13376 36139 13379
rect 40052 13376 40080 13404
rect 36127 13348 37136 13376
rect 36127 13345 36139 13348
rect 36081 13339 36139 13345
rect 33919 13280 35112 13308
rect 35161 13311 35219 13317
rect 33919 13277 33931 13280
rect 33873 13271 33931 13277
rect 35161 13277 35173 13311
rect 35207 13308 35219 13311
rect 35618 13308 35624 13320
rect 35207 13280 35624 13308
rect 35207 13277 35219 13280
rect 35161 13271 35219 13277
rect 35618 13268 35624 13280
rect 35676 13268 35682 13320
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 37108 13317 37136 13348
rect 39316 13348 40080 13376
rect 35897 13311 35955 13317
rect 35897 13308 35909 13311
rect 35860 13280 35909 13308
rect 35860 13268 35866 13280
rect 35897 13277 35909 13280
rect 35943 13277 35955 13311
rect 35897 13271 35955 13277
rect 36173 13311 36231 13317
rect 36173 13277 36185 13311
rect 36219 13277 36231 13311
rect 36173 13271 36231 13277
rect 37093 13311 37151 13317
rect 37093 13277 37105 13311
rect 37139 13308 37151 13311
rect 37366 13308 37372 13320
rect 37139 13280 37372 13308
rect 37139 13277 37151 13280
rect 37093 13271 37151 13277
rect 34514 13200 34520 13252
rect 34572 13240 34578 13252
rect 36188 13240 36216 13271
rect 37366 13268 37372 13280
rect 37424 13268 37430 13320
rect 37550 13268 37556 13320
rect 37608 13308 37614 13320
rect 37921 13311 37979 13317
rect 37921 13308 37933 13311
rect 37608 13280 37933 13308
rect 37608 13268 37614 13280
rect 37921 13277 37933 13280
rect 37967 13277 37979 13311
rect 37921 13271 37979 13277
rect 38105 13311 38163 13317
rect 38105 13277 38117 13311
rect 38151 13277 38163 13311
rect 38105 13271 38163 13277
rect 34572 13212 36216 13240
rect 34572 13200 34578 13212
rect 31076 13144 32904 13172
rect 31076 13132 31082 13144
rect 32950 13132 32956 13184
rect 33008 13172 33014 13184
rect 33137 13175 33195 13181
rect 33137 13172 33149 13175
rect 33008 13144 33149 13172
rect 33008 13132 33014 13144
rect 33137 13141 33149 13144
rect 33183 13141 33195 13175
rect 36188 13172 36216 13212
rect 37274 13200 37280 13252
rect 37332 13240 37338 13252
rect 38120 13240 38148 13271
rect 38562 13268 38568 13320
rect 38620 13268 38626 13320
rect 38746 13268 38752 13320
rect 38804 13268 38810 13320
rect 39316 13317 39344 13348
rect 39301 13311 39359 13317
rect 39301 13277 39313 13311
rect 39347 13277 39359 13311
rect 39301 13271 39359 13277
rect 40037 13311 40095 13317
rect 40037 13277 40049 13311
rect 40083 13308 40095 13311
rect 41322 13308 41328 13320
rect 40083 13280 41328 13308
rect 40083 13277 40095 13280
rect 40037 13271 40095 13277
rect 40420 13252 40448 13280
rect 41322 13268 41328 13280
rect 41380 13308 41386 13320
rect 41877 13311 41935 13317
rect 41877 13308 41889 13311
rect 41380 13280 41889 13308
rect 41380 13268 41386 13280
rect 41877 13277 41889 13280
rect 41923 13308 41935 13311
rect 41966 13308 41972 13320
rect 41923 13280 41972 13308
rect 41923 13277 41935 13280
rect 41877 13271 41935 13277
rect 41966 13268 41972 13280
rect 42024 13268 42030 13320
rect 40282 13243 40340 13249
rect 40282 13240 40294 13243
rect 37332 13212 38148 13240
rect 39500 13212 40294 13240
rect 37332 13200 37338 13212
rect 39500 13181 39528 13212
rect 40282 13209 40294 13212
rect 40328 13209 40340 13243
rect 40282 13203 40340 13209
rect 40402 13200 40408 13252
rect 40460 13200 40466 13252
rect 42150 13249 42156 13252
rect 42144 13203 42156 13249
rect 42150 13200 42156 13203
rect 42208 13200 42214 13252
rect 38013 13175 38071 13181
rect 38013 13172 38025 13175
rect 36188 13144 38025 13172
rect 33137 13135 33195 13141
rect 38013 13141 38025 13144
rect 38059 13141 38071 13175
rect 38013 13135 38071 13141
rect 39485 13175 39543 13181
rect 39485 13141 39497 13175
rect 39531 13141 39543 13175
rect 39485 13135 39543 13141
rect 41046 13132 41052 13184
rect 41104 13172 41110 13184
rect 41417 13175 41475 13181
rect 41417 13172 41429 13175
rect 41104 13144 41429 13172
rect 41104 13132 41110 13144
rect 41417 13141 41429 13144
rect 41463 13141 41475 13175
rect 41417 13135 41475 13141
rect 1104 13082 43884 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 43884 13082
rect 1104 13008 43884 13030
rect 20162 12928 20168 12980
rect 20220 12928 20226 12980
rect 21453 12971 21511 12977
rect 21453 12937 21465 12971
rect 21499 12968 21511 12971
rect 21499 12940 22094 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 22066 12900 22094 12940
rect 23290 12928 23296 12980
rect 23348 12968 23354 12980
rect 23385 12971 23443 12977
rect 23385 12968 23397 12971
rect 23348 12940 23397 12968
rect 23348 12928 23354 12940
rect 23385 12937 23397 12940
rect 23431 12937 23443 12971
rect 23385 12931 23443 12937
rect 25777 12971 25835 12977
rect 25777 12937 25789 12971
rect 25823 12968 25835 12971
rect 26234 12968 26240 12980
rect 25823 12940 26240 12968
rect 25823 12937 25835 12940
rect 25777 12931 25835 12937
rect 26234 12928 26240 12940
rect 26292 12968 26298 12980
rect 26513 12971 26571 12977
rect 26513 12968 26525 12971
rect 26292 12940 26525 12968
rect 26292 12928 26298 12940
rect 26513 12937 26525 12940
rect 26559 12968 26571 12971
rect 26602 12968 26608 12980
rect 26559 12940 26608 12968
rect 26559 12937 26571 12940
rect 26513 12931 26571 12937
rect 26602 12928 26608 12940
rect 26660 12928 26666 12980
rect 28445 12971 28503 12977
rect 28445 12937 28457 12971
rect 28491 12968 28503 12971
rect 29638 12968 29644 12980
rect 28491 12940 29644 12968
rect 28491 12937 28503 12940
rect 28445 12931 28503 12937
rect 29638 12928 29644 12940
rect 29696 12928 29702 12980
rect 31662 12928 31668 12980
rect 31720 12928 31726 12980
rect 31754 12928 31760 12980
rect 31812 12928 31818 12980
rect 31846 12928 31852 12980
rect 31904 12968 31910 12980
rect 32398 12968 32404 12980
rect 31904 12940 32404 12968
rect 31904 12928 31910 12940
rect 32398 12928 32404 12940
rect 32456 12928 32462 12980
rect 32950 12928 32956 12980
rect 33008 12928 33014 12980
rect 33318 12928 33324 12980
rect 33376 12968 33382 12980
rect 33689 12971 33747 12977
rect 33689 12968 33701 12971
rect 33376 12940 33701 12968
rect 33376 12928 33382 12940
rect 33689 12937 33701 12940
rect 33735 12937 33747 12971
rect 33689 12931 33747 12937
rect 33796 12940 36768 12968
rect 22250 12903 22308 12909
rect 22250 12900 22262 12903
rect 22066 12872 22262 12900
rect 22250 12869 22262 12872
rect 22296 12869 22308 12903
rect 22250 12863 22308 12869
rect 29178 12860 29184 12912
rect 29236 12900 29242 12912
rect 31772 12900 31800 12928
rect 29236 12872 29868 12900
rect 29236 12860 29242 12872
rect 21266 12792 21272 12844
rect 21324 12792 21330 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12832 27215 12835
rect 27338 12832 27344 12844
rect 27203 12804 27344 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 29546 12792 29552 12844
rect 29604 12841 29610 12844
rect 29604 12832 29616 12841
rect 29604 12804 29649 12832
rect 29604 12795 29616 12804
rect 29604 12792 29610 12795
rect 29840 12776 29868 12872
rect 31588 12872 31800 12900
rect 32416 12872 33640 12900
rect 30006 12792 30012 12844
rect 30064 12832 30070 12844
rect 30745 12835 30803 12841
rect 30745 12832 30757 12835
rect 30064 12804 30757 12832
rect 30064 12792 30070 12804
rect 30745 12801 30757 12804
rect 30791 12801 30803 12835
rect 30745 12795 30803 12801
rect 30929 12835 30987 12841
rect 30929 12801 30941 12835
rect 30975 12832 30987 12835
rect 31018 12832 31024 12844
rect 30975 12804 31024 12832
rect 30975 12801 30987 12804
rect 30929 12795 30987 12801
rect 29822 12724 29828 12776
rect 29880 12724 29886 12776
rect 30558 12724 30564 12776
rect 30616 12764 30622 12776
rect 30653 12767 30711 12773
rect 30653 12764 30665 12767
rect 30616 12736 30665 12764
rect 30616 12724 30622 12736
rect 30653 12733 30665 12736
rect 30699 12733 30711 12767
rect 30760 12764 30788 12795
rect 31018 12792 31024 12804
rect 31076 12792 31082 12844
rect 31588 12841 31616 12872
rect 31573 12835 31631 12841
rect 31573 12801 31585 12835
rect 31619 12801 31631 12835
rect 31573 12795 31631 12801
rect 31754 12792 31760 12844
rect 31812 12832 31818 12844
rect 32416 12832 32444 12872
rect 31812 12804 32444 12832
rect 31812 12792 31818 12804
rect 32490 12792 32496 12844
rect 32548 12792 32554 12844
rect 33612 12841 33640 12872
rect 33796 12841 33824 12940
rect 34701 12903 34759 12909
rect 34701 12869 34713 12903
rect 34747 12900 34759 12903
rect 34747 12872 34928 12900
rect 34747 12869 34759 12872
rect 34701 12863 34759 12869
rect 34900 12844 34928 12872
rect 35618 12860 35624 12912
rect 35676 12860 35682 12912
rect 36740 12900 36768 12940
rect 36814 12928 36820 12980
rect 36872 12968 36878 12980
rect 37829 12971 37887 12977
rect 37829 12968 37841 12971
rect 36872 12940 37841 12968
rect 36872 12928 36878 12940
rect 37829 12937 37841 12940
rect 37875 12937 37887 12971
rect 38746 12968 38752 12980
rect 37829 12931 37887 12937
rect 37936 12940 38752 12968
rect 37936 12900 37964 12940
rect 38746 12928 38752 12940
rect 38804 12968 38810 12980
rect 39945 12971 40003 12977
rect 39945 12968 39957 12971
rect 38804 12940 39957 12968
rect 38804 12928 38810 12940
rect 39945 12937 39957 12940
rect 39991 12937 40003 12971
rect 39945 12931 40003 12937
rect 40405 12971 40463 12977
rect 40405 12937 40417 12971
rect 40451 12968 40463 12971
rect 41046 12968 41052 12980
rect 40451 12940 41052 12968
rect 40451 12937 40463 12940
rect 40405 12931 40463 12937
rect 41046 12928 41052 12940
rect 41104 12928 41110 12980
rect 41414 12928 41420 12980
rect 41472 12968 41478 12980
rect 41874 12968 41880 12980
rect 41472 12940 41880 12968
rect 41472 12928 41478 12940
rect 41874 12928 41880 12940
rect 41932 12928 41938 12980
rect 42061 12971 42119 12977
rect 42061 12937 42073 12971
rect 42107 12968 42119 12971
rect 42150 12968 42156 12980
rect 42107 12940 42156 12968
rect 42107 12937 42119 12940
rect 42061 12931 42119 12937
rect 42150 12928 42156 12940
rect 42208 12928 42214 12980
rect 42613 12971 42671 12977
rect 42613 12937 42625 12971
rect 42659 12937 42671 12971
rect 42613 12931 42671 12937
rect 42518 12900 42524 12912
rect 36740 12872 37964 12900
rect 38028 12872 42524 12900
rect 33597 12835 33655 12841
rect 33597 12801 33609 12835
rect 33643 12801 33655 12835
rect 33597 12795 33655 12801
rect 33781 12835 33839 12841
rect 33781 12801 33793 12835
rect 33827 12801 33839 12835
rect 33781 12795 33839 12801
rect 32508 12764 32536 12792
rect 30760 12736 32536 12764
rect 32585 12767 32643 12773
rect 30653 12727 30711 12733
rect 32585 12733 32597 12767
rect 32631 12764 32643 12767
rect 32858 12764 32864 12776
rect 32631 12736 32864 12764
rect 32631 12733 32643 12736
rect 32585 12727 32643 12733
rect 30668 12696 30696 12727
rect 32858 12724 32864 12736
rect 32916 12724 32922 12776
rect 33612 12764 33640 12795
rect 34422 12792 34428 12844
rect 34480 12792 34486 12844
rect 34882 12832 34888 12844
rect 34532 12804 34888 12832
rect 34532 12764 34560 12804
rect 34882 12792 34888 12804
rect 34940 12792 34946 12844
rect 35342 12792 35348 12844
rect 35400 12832 35406 12844
rect 35805 12835 35863 12841
rect 35805 12832 35817 12835
rect 35400 12804 35817 12832
rect 35400 12792 35406 12804
rect 35805 12801 35817 12804
rect 35851 12801 35863 12835
rect 35805 12795 35863 12801
rect 36265 12835 36323 12841
rect 36265 12801 36277 12835
rect 36311 12801 36323 12835
rect 36265 12795 36323 12801
rect 36449 12835 36507 12841
rect 36449 12801 36461 12835
rect 36495 12832 36507 12835
rect 37458 12832 37464 12844
rect 36495 12804 37464 12832
rect 36495 12801 36507 12804
rect 36449 12795 36507 12801
rect 33612 12736 34560 12764
rect 34606 12724 34612 12776
rect 34664 12724 34670 12776
rect 35437 12767 35495 12773
rect 35437 12733 35449 12767
rect 35483 12764 35495 12767
rect 35986 12764 35992 12776
rect 35483 12736 35992 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35986 12724 35992 12736
rect 36044 12764 36050 12776
rect 36280 12764 36308 12795
rect 37458 12792 37464 12804
rect 37516 12792 37522 12844
rect 38028 12841 38056 12872
rect 38013 12835 38071 12841
rect 38013 12801 38025 12835
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 38197 12835 38255 12841
rect 38197 12801 38209 12835
rect 38243 12832 38255 12835
rect 38562 12832 38568 12844
rect 38243 12804 38568 12832
rect 38243 12801 38255 12804
rect 38197 12795 38255 12801
rect 38562 12792 38568 12804
rect 38620 12832 38626 12844
rect 39040 12841 39068 12872
rect 42518 12860 42524 12872
rect 42576 12860 42582 12912
rect 38749 12835 38807 12841
rect 38749 12832 38761 12835
rect 38620 12804 38761 12832
rect 38620 12792 38626 12804
rect 38749 12801 38761 12804
rect 38795 12801 38807 12835
rect 38749 12795 38807 12801
rect 39025 12835 39083 12841
rect 39025 12801 39037 12835
rect 39071 12801 39083 12835
rect 39025 12795 39083 12801
rect 40313 12835 40371 12841
rect 40313 12801 40325 12835
rect 40359 12832 40371 12835
rect 41230 12832 41236 12844
rect 40359 12804 41236 12832
rect 40359 12801 40371 12804
rect 40313 12795 40371 12801
rect 41230 12792 41236 12804
rect 41288 12792 41294 12844
rect 41877 12835 41935 12841
rect 41877 12801 41889 12835
rect 41923 12832 41935 12835
rect 42628 12832 42656 12931
rect 42978 12928 42984 12980
rect 43036 12928 43042 12980
rect 43070 12928 43076 12980
rect 43128 12928 43134 12980
rect 42996 12900 43024 12928
rect 43346 12900 43352 12912
rect 42996 12872 43352 12900
rect 43346 12860 43352 12872
rect 43404 12860 43410 12912
rect 41923 12804 42656 12832
rect 41923 12801 41935 12804
rect 41877 12795 41935 12801
rect 36044 12736 36308 12764
rect 36044 12724 36050 12736
rect 38654 12724 38660 12776
rect 38712 12724 38718 12776
rect 40589 12767 40647 12773
rect 40589 12733 40601 12767
rect 40635 12764 40647 12767
rect 41046 12764 41052 12776
rect 40635 12736 41052 12764
rect 40635 12733 40647 12736
rect 40589 12727 40647 12733
rect 41046 12724 41052 12736
rect 41104 12724 41110 12776
rect 42886 12724 42892 12776
rect 42944 12764 42950 12776
rect 43165 12767 43223 12773
rect 43165 12764 43177 12767
rect 42944 12736 43177 12764
rect 42944 12724 42950 12736
rect 43165 12733 43177 12736
rect 43211 12733 43223 12767
rect 43165 12727 43223 12733
rect 32766 12696 32772 12708
rect 30668 12668 32772 12696
rect 32766 12656 32772 12668
rect 32824 12656 32830 12708
rect 34698 12656 34704 12708
rect 34756 12696 34762 12708
rect 36265 12699 36323 12705
rect 36265 12696 36277 12699
rect 34756 12668 36277 12696
rect 34756 12656 34762 12668
rect 36265 12665 36277 12668
rect 36311 12665 36323 12699
rect 36265 12659 36323 12665
rect 27341 12631 27399 12637
rect 27341 12597 27353 12631
rect 27387 12628 27399 12631
rect 27430 12628 27436 12640
rect 27387 12600 27436 12628
rect 27387 12597 27399 12600
rect 27341 12591 27399 12597
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 30926 12588 30932 12640
rect 30984 12628 30990 12640
rect 31113 12631 31171 12637
rect 31113 12628 31125 12631
rect 30984 12600 31125 12628
rect 30984 12588 30990 12600
rect 31113 12597 31125 12600
rect 31159 12597 31171 12631
rect 31113 12591 31171 12597
rect 32122 12588 32128 12640
rect 32180 12628 32186 12640
rect 32309 12631 32367 12637
rect 32309 12628 32321 12631
rect 32180 12600 32321 12628
rect 32180 12588 32186 12600
rect 32309 12597 32321 12600
rect 32355 12597 32367 12631
rect 32309 12591 32367 12597
rect 34241 12631 34299 12637
rect 34241 12597 34253 12631
rect 34287 12628 34299 12631
rect 34330 12628 34336 12640
rect 34287 12600 34336 12628
rect 34287 12597 34299 12600
rect 34241 12591 34299 12597
rect 34330 12588 34336 12600
rect 34388 12588 34394 12640
rect 34609 12631 34667 12637
rect 34609 12597 34621 12631
rect 34655 12628 34667 12631
rect 34790 12628 34796 12640
rect 34655 12600 34796 12628
rect 34655 12597 34667 12600
rect 34609 12591 34667 12597
rect 34790 12588 34796 12600
rect 34848 12588 34854 12640
rect 1104 12538 43884 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 43884 12538
rect 1104 12464 43884 12486
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 26418 12384 26424 12436
rect 26476 12384 26482 12436
rect 27338 12384 27344 12436
rect 27396 12384 27402 12436
rect 30558 12424 30564 12436
rect 28920 12396 30564 12424
rect 26436 12356 26464 12384
rect 28920 12368 28948 12396
rect 30558 12384 30564 12396
rect 30616 12424 30622 12436
rect 31110 12424 31116 12436
rect 30616 12396 31116 12424
rect 30616 12384 30622 12396
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 32214 12384 32220 12436
rect 32272 12384 32278 12436
rect 37090 12384 37096 12436
rect 37148 12384 37154 12436
rect 38654 12384 38660 12436
rect 38712 12384 38718 12436
rect 40586 12384 40592 12436
rect 40644 12384 40650 12436
rect 41506 12384 41512 12436
rect 41564 12384 41570 12436
rect 28902 12356 28908 12368
rect 26436 12328 28908 12356
rect 28902 12316 28908 12328
rect 28960 12316 28966 12368
rect 29454 12316 29460 12368
rect 29512 12356 29518 12368
rect 29917 12359 29975 12365
rect 29917 12356 29929 12359
rect 29512 12328 29929 12356
rect 29512 12316 29518 12328
rect 29917 12325 29929 12328
rect 29963 12356 29975 12359
rect 31754 12356 31760 12368
rect 29963 12328 30604 12356
rect 29963 12325 29975 12328
rect 29917 12319 29975 12325
rect 26602 12288 26608 12300
rect 26160 12260 26608 12288
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 25590 12180 25596 12232
rect 25648 12180 25654 12232
rect 26160 12229 26188 12260
rect 26602 12248 26608 12260
rect 26660 12288 26666 12300
rect 27985 12291 28043 12297
rect 27985 12288 27997 12291
rect 26660 12260 27997 12288
rect 26660 12248 26666 12260
rect 27985 12257 27997 12260
rect 28031 12288 28043 12291
rect 30466 12288 30472 12300
rect 28031 12260 28948 12288
rect 28031 12257 28043 12260
rect 27985 12251 28043 12257
rect 26145 12223 26203 12229
rect 26145 12189 26157 12223
rect 26191 12189 26203 12223
rect 26145 12183 26203 12189
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12220 27859 12223
rect 28810 12220 28816 12232
rect 27847 12192 28816 12220
rect 27847 12189 27859 12192
rect 27801 12183 27859 12189
rect 28810 12180 28816 12192
rect 28868 12180 28874 12232
rect 25406 12044 25412 12096
rect 25464 12044 25470 12096
rect 27709 12087 27767 12093
rect 27709 12053 27721 12087
rect 27755 12084 27767 12087
rect 28442 12084 28448 12096
rect 27755 12056 28448 12084
rect 27755 12053 27767 12056
rect 27709 12047 27767 12053
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 28629 12087 28687 12093
rect 28629 12053 28641 12087
rect 28675 12084 28687 12087
rect 28920 12084 28948 12260
rect 29748 12260 30472 12288
rect 29748 12229 29776 12260
rect 30466 12248 30472 12260
rect 30524 12248 30530 12300
rect 30576 12229 30604 12328
rect 30760 12328 31760 12356
rect 29733 12223 29791 12229
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 29917 12223 29975 12229
rect 29917 12189 29929 12223
rect 29963 12189 29975 12223
rect 29917 12183 29975 12189
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 29932 12152 29960 12183
rect 30650 12180 30656 12232
rect 30708 12180 30714 12232
rect 30760 12152 30788 12328
rect 31754 12316 31760 12328
rect 31812 12316 31818 12368
rect 35805 12359 35863 12365
rect 35805 12325 35817 12359
rect 35851 12356 35863 12359
rect 39206 12356 39212 12368
rect 35851 12328 39212 12356
rect 35851 12325 35863 12328
rect 35805 12319 35863 12325
rect 32122 12288 32128 12300
rect 30852 12260 32128 12288
rect 30852 12229 30880 12260
rect 32122 12248 32128 12260
rect 32180 12248 32186 12300
rect 32306 12248 32312 12300
rect 32364 12248 32370 12300
rect 32858 12248 32864 12300
rect 32916 12288 32922 12300
rect 33965 12291 34023 12297
rect 33965 12288 33977 12291
rect 32916 12260 33977 12288
rect 32916 12248 32922 12260
rect 33965 12257 33977 12260
rect 34011 12257 34023 12291
rect 33965 12251 34023 12257
rect 34054 12248 34060 12300
rect 34112 12288 34118 12300
rect 34885 12291 34943 12297
rect 34885 12288 34897 12291
rect 34112 12260 34897 12288
rect 34112 12248 34118 12260
rect 34885 12257 34897 12260
rect 34931 12257 34943 12291
rect 36265 12291 36323 12297
rect 36265 12288 36277 12291
rect 34885 12251 34943 12257
rect 34992 12260 36277 12288
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 32214 12180 32220 12232
rect 32272 12180 32278 12232
rect 33781 12223 33839 12229
rect 33781 12189 33793 12223
rect 33827 12189 33839 12223
rect 33781 12183 33839 12189
rect 29932 12124 30788 12152
rect 32677 12155 32735 12161
rect 32677 12121 32689 12155
rect 32723 12152 32735 12155
rect 33597 12155 33655 12161
rect 33597 12152 33609 12155
rect 32723 12124 33609 12152
rect 32723 12121 32735 12124
rect 32677 12115 32735 12121
rect 33597 12121 33609 12124
rect 33643 12121 33655 12155
rect 33796 12152 33824 12183
rect 34146 12180 34152 12232
rect 34204 12180 34210 12232
rect 34330 12180 34336 12232
rect 34388 12180 34394 12232
rect 34992 12152 35020 12260
rect 36265 12257 36277 12260
rect 36311 12288 36323 12291
rect 36630 12288 36636 12300
rect 36311 12260 36636 12288
rect 36311 12257 36323 12260
rect 36265 12251 36323 12257
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12220 35311 12223
rect 35526 12220 35532 12232
rect 35299 12192 35532 12220
rect 35299 12189 35311 12192
rect 35253 12183 35311 12189
rect 35526 12180 35532 12192
rect 35584 12180 35590 12232
rect 36357 12223 36415 12229
rect 36357 12189 36369 12223
rect 36403 12189 36415 12223
rect 36357 12183 36415 12189
rect 36541 12223 36599 12229
rect 36541 12189 36553 12223
rect 36587 12220 36599 12223
rect 36587 12192 37504 12220
rect 36587 12189 36599 12192
rect 36541 12183 36599 12189
rect 33796 12124 35020 12152
rect 35069 12155 35127 12161
rect 33597 12115 33655 12121
rect 35069 12121 35081 12155
rect 35115 12152 35127 12155
rect 36372 12152 36400 12183
rect 37274 12152 37280 12164
rect 35115 12124 37280 12152
rect 35115 12121 35127 12124
rect 35069 12115 35127 12121
rect 29181 12087 29239 12093
rect 29181 12084 29193 12087
rect 28675 12056 29193 12084
rect 28675 12053 28687 12056
rect 28629 12047 28687 12053
rect 29181 12053 29193 12056
rect 29227 12084 29239 12087
rect 30006 12084 30012 12096
rect 29227 12056 30012 12084
rect 29227 12053 29239 12056
rect 29181 12047 29239 12053
rect 30006 12044 30012 12056
rect 30064 12044 30070 12096
rect 30377 12087 30435 12093
rect 30377 12053 30389 12087
rect 30423 12084 30435 12087
rect 30834 12084 30840 12096
rect 30423 12056 30840 12084
rect 30423 12053 30435 12056
rect 30377 12047 30435 12053
rect 30834 12044 30840 12056
rect 30892 12044 30898 12096
rect 32030 12044 32036 12096
rect 32088 12044 32094 12096
rect 32766 12044 32772 12096
rect 32824 12084 32830 12096
rect 33870 12084 33876 12096
rect 32824 12056 33876 12084
rect 32824 12044 32830 12056
rect 33870 12044 33876 12056
rect 33928 12044 33934 12096
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 35084 12084 35112 12115
rect 37274 12112 37280 12124
rect 37332 12112 37338 12164
rect 37476 12161 37504 12192
rect 38286 12180 38292 12232
rect 38344 12220 38350 12232
rect 38396 12229 38424 12328
rect 39206 12316 39212 12328
rect 39264 12356 39270 12368
rect 40037 12359 40095 12365
rect 40037 12356 40049 12359
rect 39264 12328 40049 12356
rect 39264 12316 39270 12328
rect 40037 12325 40049 12328
rect 40083 12325 40095 12359
rect 40037 12319 40095 12325
rect 41966 12248 41972 12300
rect 42024 12248 42030 12300
rect 38381 12223 38439 12229
rect 38381 12220 38393 12223
rect 38344 12192 38393 12220
rect 38344 12180 38350 12192
rect 38381 12189 38393 12192
rect 38427 12189 38439 12223
rect 38381 12183 38439 12189
rect 38654 12180 38660 12232
rect 38712 12220 38718 12232
rect 39209 12223 39267 12229
rect 39209 12220 39221 12223
rect 38712 12192 39221 12220
rect 38712 12180 38718 12192
rect 39209 12189 39221 12192
rect 39255 12189 39267 12223
rect 39209 12183 39267 12189
rect 39390 12180 39396 12232
rect 39448 12180 39454 12232
rect 37461 12155 37519 12161
rect 37461 12121 37473 12155
rect 37507 12121 37519 12155
rect 37461 12115 37519 12121
rect 34664 12056 35112 12084
rect 37476 12084 37504 12115
rect 42058 12112 42064 12164
rect 42116 12152 42122 12164
rect 42214 12155 42272 12161
rect 42214 12152 42226 12155
rect 42116 12124 42226 12152
rect 42116 12112 42122 12124
rect 42214 12121 42226 12124
rect 42260 12121 42272 12155
rect 42214 12115 42272 12121
rect 37642 12084 37648 12096
rect 37476 12056 37648 12084
rect 34664 12044 34670 12056
rect 37642 12044 37648 12056
rect 37700 12084 37706 12096
rect 39209 12087 39267 12093
rect 39209 12084 39221 12087
rect 37700 12056 39221 12084
rect 37700 12044 37706 12056
rect 39209 12053 39221 12056
rect 39255 12053 39267 12087
rect 39209 12047 39267 12053
rect 43070 12044 43076 12096
rect 43128 12084 43134 12096
rect 43349 12087 43407 12093
rect 43349 12084 43361 12087
rect 43128 12056 43361 12084
rect 43128 12044 43134 12056
rect 43349 12053 43361 12056
rect 43395 12053 43407 12087
rect 43349 12047 43407 12053
rect 1104 11994 43884 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 43884 11994
rect 1104 11920 43884 11942
rect 26142 11840 26148 11892
rect 26200 11880 26206 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26200 11852 26525 11880
rect 26200 11840 26206 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 26513 11843 26571 11849
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 28500 11852 28549 11880
rect 28500 11840 28506 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 28537 11843 28595 11849
rect 29454 11840 29460 11892
rect 29512 11840 29518 11892
rect 30834 11840 30840 11892
rect 30892 11840 30898 11892
rect 32214 11840 32220 11892
rect 32272 11880 32278 11892
rect 32582 11880 32588 11892
rect 32272 11852 32588 11880
rect 32272 11840 32278 11852
rect 32582 11840 32588 11852
rect 32640 11840 32646 11892
rect 34514 11880 34520 11892
rect 33152 11852 34520 11880
rect 25406 11821 25412 11824
rect 25400 11812 25412 11821
rect 25367 11784 25412 11812
rect 25400 11775 25412 11784
rect 25406 11772 25412 11775
rect 25464 11772 25470 11824
rect 27430 11821 27436 11824
rect 27424 11812 27436 11821
rect 27391 11784 27436 11812
rect 27424 11775 27436 11784
rect 27430 11772 27436 11775
rect 27488 11772 27494 11824
rect 27522 11772 27528 11824
rect 27580 11812 27586 11824
rect 32030 11812 32036 11824
rect 27580 11784 32036 11812
rect 27580 11772 27586 11784
rect 32030 11772 32036 11784
rect 32088 11772 32094 11824
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 27154 11704 27160 11756
rect 27212 11704 27218 11756
rect 29362 11704 29368 11756
rect 29420 11704 29426 11756
rect 30745 11747 30803 11753
rect 30745 11713 30757 11747
rect 30791 11744 30803 11747
rect 31754 11744 31760 11756
rect 30791 11716 31760 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 31754 11704 31760 11716
rect 31812 11744 31818 11756
rect 32674 11744 32680 11756
rect 31812 11716 32680 11744
rect 31812 11704 31818 11716
rect 32674 11704 32680 11716
rect 32732 11704 32738 11756
rect 32766 11704 32772 11756
rect 32824 11704 32830 11756
rect 33152 11753 33180 11852
rect 34514 11840 34520 11852
rect 34572 11840 34578 11892
rect 34974 11840 34980 11892
rect 35032 11880 35038 11892
rect 35894 11880 35900 11892
rect 35032 11852 35900 11880
rect 35032 11840 35038 11852
rect 35894 11840 35900 11852
rect 35952 11840 35958 11892
rect 37366 11840 37372 11892
rect 37424 11880 37430 11892
rect 38289 11883 38347 11889
rect 38289 11880 38301 11883
rect 37424 11852 38301 11880
rect 37424 11840 37430 11852
rect 38289 11849 38301 11852
rect 38335 11849 38347 11883
rect 38289 11843 38347 11849
rect 39390 11840 39396 11892
rect 39448 11880 39454 11892
rect 40497 11883 40555 11889
rect 40497 11880 40509 11883
rect 39448 11852 40509 11880
rect 39448 11840 39454 11852
rect 40497 11849 40509 11852
rect 40543 11849 40555 11883
rect 40497 11843 40555 11849
rect 40862 11840 40868 11892
rect 40920 11840 40926 11892
rect 42058 11840 42064 11892
rect 42116 11840 42122 11892
rect 42610 11840 42616 11892
rect 42668 11840 42674 11892
rect 43070 11840 43076 11892
rect 43128 11840 43134 11892
rect 33873 11815 33931 11821
rect 33873 11781 33885 11815
rect 33919 11812 33931 11815
rect 34701 11815 34759 11821
rect 34701 11812 34713 11815
rect 33919 11784 34713 11812
rect 33919 11781 33931 11784
rect 33873 11775 33931 11781
rect 34701 11781 34713 11784
rect 34747 11812 34759 11815
rect 34747 11784 35848 11812
rect 34747 11781 34759 11784
rect 34701 11775 34759 11781
rect 32861 11747 32919 11753
rect 32861 11713 32873 11747
rect 32907 11713 32919 11747
rect 32861 11707 32919 11713
rect 32953 11747 33011 11753
rect 32953 11713 32965 11747
rect 32999 11713 33011 11747
rect 32953 11707 33011 11713
rect 33137 11747 33195 11753
rect 33137 11713 33149 11747
rect 33183 11713 33195 11747
rect 33137 11707 33195 11713
rect 33965 11747 34023 11753
rect 33965 11713 33977 11747
rect 34011 11744 34023 11747
rect 34054 11744 34060 11756
rect 34011 11716 34060 11744
rect 34011 11713 34023 11716
rect 33965 11707 34023 11713
rect 29178 11568 29184 11620
rect 29236 11608 29242 11620
rect 29380 11608 29408 11704
rect 29641 11679 29699 11685
rect 29641 11645 29653 11679
rect 29687 11676 29699 11679
rect 30006 11676 30012 11688
rect 29687 11648 30012 11676
rect 29687 11645 29699 11648
rect 29641 11639 29699 11645
rect 30006 11636 30012 11648
rect 30064 11636 30070 11688
rect 30558 11636 30564 11688
rect 30616 11676 30622 11688
rect 30926 11676 30932 11688
rect 30616 11648 30932 11676
rect 30616 11636 30622 11648
rect 30926 11636 30932 11648
rect 30984 11636 30990 11688
rect 31018 11636 31024 11688
rect 31076 11676 31082 11688
rect 32876 11676 32904 11707
rect 31076 11648 32904 11676
rect 32968 11676 32996 11707
rect 34054 11704 34060 11716
rect 34112 11704 34118 11756
rect 34609 11747 34667 11753
rect 34609 11713 34621 11747
rect 34655 11713 34667 11747
rect 34609 11707 34667 11713
rect 33318 11676 33324 11688
rect 32968 11648 33324 11676
rect 31076 11636 31082 11648
rect 31573 11611 31631 11617
rect 31573 11608 31585 11611
rect 29236 11580 31585 11608
rect 29236 11568 29242 11580
rect 31573 11577 31585 11580
rect 31619 11577 31631 11611
rect 32876 11608 32904 11648
rect 33318 11636 33324 11648
rect 33376 11676 33382 11688
rect 34624 11676 34652 11707
rect 34790 11704 34796 11756
rect 34848 11704 34854 11756
rect 34974 11704 34980 11756
rect 35032 11704 35038 11756
rect 35820 11753 35848 11784
rect 37274 11772 37280 11824
rect 37332 11812 37338 11824
rect 39408 11812 39436 11840
rect 37332 11784 37780 11812
rect 37332 11772 37338 11784
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11713 35679 11747
rect 35621 11707 35679 11713
rect 35805 11747 35863 11753
rect 35805 11713 35817 11747
rect 35851 11713 35863 11747
rect 35805 11707 35863 11713
rect 35897 11747 35955 11753
rect 35897 11713 35909 11747
rect 35943 11744 35955 11747
rect 36170 11744 36176 11756
rect 35943 11716 36176 11744
rect 35943 11713 35955 11716
rect 35897 11707 35955 11713
rect 35636 11676 35664 11707
rect 36170 11704 36176 11716
rect 36228 11744 36234 11756
rect 36633 11747 36691 11753
rect 36633 11744 36645 11747
rect 36228 11716 36645 11744
rect 36228 11704 36234 11716
rect 36633 11713 36645 11716
rect 36679 11713 36691 11747
rect 36633 11707 36691 11713
rect 36817 11747 36875 11753
rect 36817 11713 36829 11747
rect 36863 11744 36875 11747
rect 37461 11747 37519 11753
rect 37461 11744 37473 11747
rect 36863 11716 37473 11744
rect 36863 11713 36875 11716
rect 36817 11707 36875 11713
rect 37461 11713 37473 11716
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 37642 11704 37648 11756
rect 37700 11704 37706 11756
rect 37752 11753 37780 11784
rect 38488 11784 39436 11812
rect 38488 11753 38516 11784
rect 39666 11772 39672 11824
rect 39724 11812 39730 11824
rect 40034 11812 40040 11824
rect 39724 11784 40040 11812
rect 39724 11772 39730 11784
rect 40034 11772 40040 11784
rect 40092 11772 40098 11824
rect 37737 11747 37795 11753
rect 37737 11713 37749 11747
rect 37783 11713 37795 11747
rect 37737 11707 37795 11713
rect 38473 11747 38531 11753
rect 38473 11713 38485 11747
rect 38519 11713 38531 11747
rect 38473 11707 38531 11713
rect 38654 11704 38660 11756
rect 38712 11704 38718 11756
rect 39761 11747 39819 11753
rect 39761 11713 39773 11747
rect 39807 11744 39819 11747
rect 40126 11744 40132 11756
rect 39807 11716 40132 11744
rect 39807 11713 39819 11716
rect 39761 11707 39819 11713
rect 40126 11704 40132 11716
rect 40184 11704 40190 11756
rect 40957 11747 41015 11753
rect 40957 11713 40969 11747
rect 41003 11744 41015 11747
rect 41138 11744 41144 11756
rect 41003 11716 41144 11744
rect 41003 11713 41015 11716
rect 40957 11707 41015 11713
rect 41138 11704 41144 11716
rect 41196 11704 41202 11756
rect 41877 11747 41935 11753
rect 41877 11713 41889 11747
rect 41923 11744 41935 11747
rect 42334 11744 42340 11756
rect 41923 11716 42340 11744
rect 41923 11713 41935 11716
rect 41877 11707 41935 11713
rect 42334 11704 42340 11716
rect 42392 11704 42398 11756
rect 42978 11704 42984 11756
rect 43036 11704 43042 11756
rect 33376 11648 35664 11676
rect 39945 11679 40003 11685
rect 33376 11636 33382 11648
rect 39945 11645 39957 11679
rect 39991 11676 40003 11679
rect 41046 11676 41052 11688
rect 39991 11648 41052 11676
rect 39991 11645 40003 11648
rect 39945 11639 40003 11645
rect 41046 11636 41052 11648
rect 41104 11636 41110 11688
rect 43162 11636 43168 11688
rect 43220 11636 43226 11688
rect 34974 11608 34980 11620
rect 32876 11580 34980 11608
rect 31573 11571 31631 11577
rect 34974 11568 34980 11580
rect 35032 11568 35038 11620
rect 28994 11500 29000 11552
rect 29052 11500 29058 11552
rect 30374 11500 30380 11552
rect 30432 11500 30438 11552
rect 34422 11500 34428 11552
rect 34480 11500 34486 11552
rect 35434 11500 35440 11552
rect 35492 11500 35498 11552
rect 38378 11500 38384 11552
rect 38436 11540 38442 11552
rect 39301 11543 39359 11549
rect 39301 11540 39313 11543
rect 38436 11512 39313 11540
rect 38436 11500 38442 11512
rect 39301 11509 39313 11512
rect 39347 11509 39359 11543
rect 39301 11503 39359 11509
rect 1104 11450 43884 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 43884 11450
rect 1104 11376 43884 11398
rect 25590 11296 25596 11348
rect 25648 11296 25654 11348
rect 29178 11296 29184 11348
rect 29236 11296 29242 11348
rect 30650 11296 30656 11348
rect 30708 11296 30714 11348
rect 31018 11296 31024 11348
rect 31076 11336 31082 11348
rect 31113 11339 31171 11345
rect 31113 11336 31125 11339
rect 31076 11308 31125 11336
rect 31076 11296 31082 11308
rect 31113 11305 31125 11308
rect 31159 11336 31171 11339
rect 31938 11336 31944 11348
rect 31159 11308 31944 11336
rect 31159 11305 31171 11308
rect 31113 11299 31171 11305
rect 31938 11296 31944 11308
rect 31996 11296 32002 11348
rect 32214 11296 32220 11348
rect 32272 11296 32278 11348
rect 37001 11339 37059 11345
rect 37001 11336 37013 11339
rect 32692 11308 37013 11336
rect 27522 11268 27528 11280
rect 26068 11240 27528 11268
rect 26068 11209 26096 11240
rect 27522 11228 27528 11240
rect 27580 11228 27586 11280
rect 30668 11268 30696 11296
rect 32692 11268 32720 11308
rect 37001 11305 37013 11308
rect 37047 11305 37059 11339
rect 41046 11336 41052 11348
rect 37001 11299 37059 11305
rect 38948 11308 41052 11336
rect 30668 11240 32720 11268
rect 36541 11271 36599 11277
rect 36541 11237 36553 11271
rect 36587 11268 36599 11271
rect 36906 11268 36912 11280
rect 36587 11240 36912 11268
rect 36587 11237 36599 11240
rect 36541 11231 36599 11237
rect 36906 11228 36912 11240
rect 36964 11228 36970 11280
rect 26053 11203 26111 11209
rect 26053 11169 26065 11203
rect 26099 11169 26111 11203
rect 26053 11163 26111 11169
rect 26237 11203 26295 11209
rect 26237 11169 26249 11203
rect 26283 11200 26295 11203
rect 26418 11200 26424 11212
rect 26283 11172 26424 11200
rect 26283 11169 26295 11172
rect 26237 11163 26295 11169
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 27154 11160 27160 11212
rect 27212 11200 27218 11212
rect 27801 11203 27859 11209
rect 27801 11200 27813 11203
rect 27212 11172 27813 11200
rect 27212 11160 27218 11172
rect 27801 11169 27813 11172
rect 27847 11169 27859 11203
rect 27801 11163 27859 11169
rect 33594 11160 33600 11212
rect 33652 11200 33658 11212
rect 35161 11203 35219 11209
rect 35161 11200 35173 11203
rect 33652 11172 35173 11200
rect 33652 11160 33658 11172
rect 35161 11169 35173 11172
rect 35207 11169 35219 11203
rect 37642 11200 37648 11212
rect 35161 11163 35219 11169
rect 37016 11172 37648 11200
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11132 29791 11135
rect 29822 11132 29828 11144
rect 29779 11104 29828 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 29822 11092 29828 11104
rect 29880 11092 29886 11144
rect 34146 11092 34152 11144
rect 34204 11092 34210 11144
rect 37016 11141 37044 11172
rect 37642 11160 37648 11172
rect 37700 11160 37706 11212
rect 38378 11200 38384 11212
rect 38120 11172 38384 11200
rect 37001 11135 37059 11141
rect 34256 11104 35572 11132
rect 25961 11067 26019 11073
rect 25961 11033 25973 11067
rect 26007 11064 26019 11067
rect 26142 11064 26148 11076
rect 26007 11036 26148 11064
rect 26007 11033 26019 11036
rect 25961 11027 26019 11033
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 28068 11067 28126 11073
rect 28068 11033 28080 11067
rect 28114 11064 28126 11067
rect 28350 11064 28356 11076
rect 28114 11036 28356 11064
rect 28114 11033 28126 11036
rect 28068 11027 28126 11033
rect 28350 11024 28356 11036
rect 28408 11024 28414 11076
rect 30000 11067 30058 11073
rect 30000 11033 30012 11067
rect 30046 11064 30058 11067
rect 30558 11064 30564 11076
rect 30046 11036 30564 11064
rect 30046 11033 30058 11036
rect 30000 11027 30058 11033
rect 30558 11024 30564 11036
rect 30616 11024 30622 11076
rect 33134 11024 33140 11076
rect 33192 11064 33198 11076
rect 33330 11067 33388 11073
rect 33330 11064 33342 11067
rect 33192 11036 33342 11064
rect 33192 11024 33198 11036
rect 33330 11033 33342 11036
rect 33376 11033 33388 11067
rect 33330 11027 33388 11033
rect 33686 11024 33692 11076
rect 33744 11064 33750 11076
rect 34256 11064 34284 11104
rect 35406 11067 35464 11073
rect 35406 11064 35418 11067
rect 33744 11036 34284 11064
rect 34348 11036 35418 11064
rect 33744 11024 33750 11036
rect 34348 11005 34376 11036
rect 35406 11033 35418 11036
rect 35452 11033 35464 11067
rect 35544 11064 35572 11104
rect 37001 11101 37013 11135
rect 37047 11101 37059 11135
rect 37001 11095 37059 11101
rect 37185 11135 37243 11141
rect 37185 11101 37197 11135
rect 37231 11132 37243 11135
rect 37274 11132 37280 11144
rect 37231 11104 37280 11132
rect 37231 11101 37243 11104
rect 37185 11095 37243 11101
rect 37274 11092 37280 11104
rect 37332 11092 37338 11144
rect 38120 11141 38148 11172
rect 38378 11160 38384 11172
rect 38436 11160 38442 11212
rect 38948 11209 38976 11308
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 41138 11296 41144 11348
rect 41196 11336 41202 11348
rect 41785 11339 41843 11345
rect 41785 11336 41797 11339
rect 41196 11308 41797 11336
rect 41196 11296 41202 11308
rect 41785 11305 41797 11308
rect 41831 11305 41843 11339
rect 41785 11299 41843 11305
rect 42334 11296 42340 11348
rect 42392 11296 42398 11348
rect 42978 11336 42984 11348
rect 42720 11308 42984 11336
rect 38933 11203 38991 11209
rect 38933 11169 38945 11203
rect 38979 11169 38991 11203
rect 38933 11163 38991 11169
rect 38105 11135 38163 11141
rect 38105 11101 38117 11135
rect 38151 11101 38163 11135
rect 38105 11095 38163 11101
rect 38286 11092 38292 11144
rect 38344 11092 38350 11144
rect 38396 11104 40264 11132
rect 38396 11064 38424 11104
rect 35544 11036 38424 11064
rect 39025 11067 39083 11073
rect 35406 11027 35464 11033
rect 39025 11033 39037 11067
rect 39071 11064 39083 11067
rect 40126 11064 40132 11076
rect 39071 11036 40132 11064
rect 39071 11033 39083 11036
rect 39025 11027 39083 11033
rect 40126 11024 40132 11036
rect 40184 11024 40190 11076
rect 40236 11064 40264 11104
rect 40402 11092 40408 11144
rect 40460 11092 40466 11144
rect 42720 11141 42748 11308
rect 42978 11296 42984 11308
rect 43036 11296 43042 11348
rect 43070 11268 43076 11280
rect 42812 11240 43076 11268
rect 42812 11209 42840 11240
rect 43070 11228 43076 11240
rect 43128 11228 43134 11280
rect 42797 11203 42855 11209
rect 42797 11169 42809 11203
rect 42843 11169 42855 11203
rect 42797 11163 42855 11169
rect 42886 11160 42892 11212
rect 42944 11160 42950 11212
rect 42705 11135 42763 11141
rect 42705 11132 42717 11135
rect 40880 11104 42717 11132
rect 40678 11073 40684 11076
rect 40236 11036 40632 11064
rect 34333 10999 34391 11005
rect 34333 10965 34345 10999
rect 34379 10965 34391 10999
rect 34333 10959 34391 10965
rect 37918 10956 37924 11008
rect 37976 10956 37982 11008
rect 39114 10956 39120 11008
rect 39172 10956 39178 11008
rect 39390 10956 39396 11008
rect 39448 10996 39454 11008
rect 39485 10999 39543 11005
rect 39485 10996 39497 10999
rect 39448 10968 39497 10996
rect 39448 10956 39454 10968
rect 39485 10965 39497 10968
rect 39531 10965 39543 10999
rect 40604 10996 40632 11036
rect 40672 11027 40684 11073
rect 40678 11024 40684 11027
rect 40736 11024 40742 11076
rect 40880 10996 40908 11104
rect 42705 11101 42717 11104
rect 42751 11101 42763 11135
rect 42705 11095 42763 11101
rect 41046 11024 41052 11076
rect 41104 11064 41110 11076
rect 42904 11064 42932 11160
rect 41104 11036 42932 11064
rect 41104 11024 41110 11036
rect 40604 10968 40908 10996
rect 39485 10959 39543 10965
rect 1104 10906 43884 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 43884 10906
rect 1104 10832 43884 10854
rect 28350 10752 28356 10804
rect 28408 10752 28414 10804
rect 29917 10795 29975 10801
rect 29917 10761 29929 10795
rect 29963 10761 29975 10795
rect 29917 10755 29975 10761
rect 29932 10724 29960 10755
rect 30006 10752 30012 10804
rect 30064 10792 30070 10804
rect 30064 10764 30788 10792
rect 30064 10752 30070 10764
rect 30622 10727 30680 10733
rect 30622 10724 30634 10727
rect 29932 10696 30634 10724
rect 30622 10693 30634 10696
rect 30668 10693 30680 10727
rect 30760 10724 30788 10764
rect 31754 10752 31760 10804
rect 31812 10752 31818 10804
rect 32401 10795 32459 10801
rect 32401 10761 32413 10795
rect 32447 10792 32459 10795
rect 33134 10792 33140 10804
rect 32447 10764 33140 10792
rect 32447 10761 32459 10764
rect 32401 10755 32459 10761
rect 33134 10752 33140 10764
rect 33192 10752 33198 10804
rect 34146 10752 34152 10804
rect 34204 10792 34210 10804
rect 34425 10795 34483 10801
rect 34425 10792 34437 10795
rect 34204 10764 34437 10792
rect 34204 10752 34210 10764
rect 34425 10761 34437 10764
rect 34471 10761 34483 10795
rect 34425 10755 34483 10761
rect 34885 10795 34943 10801
rect 34885 10761 34897 10795
rect 34931 10792 34943 10795
rect 35434 10792 35440 10804
rect 34931 10764 35440 10792
rect 34931 10761 34943 10764
rect 34885 10755 34943 10761
rect 35434 10752 35440 10764
rect 35492 10752 35498 10804
rect 35713 10795 35771 10801
rect 35713 10761 35725 10795
rect 35759 10792 35771 10795
rect 36906 10792 36912 10804
rect 35759 10764 36912 10792
rect 35759 10761 35771 10764
rect 35713 10755 35771 10761
rect 33965 10727 34023 10733
rect 33965 10724 33977 10727
rect 30760 10696 33977 10724
rect 30622 10687 30680 10693
rect 33965 10693 33977 10696
rect 34011 10724 34023 10727
rect 34011 10696 35020 10724
rect 34011 10693 34023 10696
rect 33965 10687 34023 10693
rect 28537 10659 28595 10665
rect 28537 10625 28549 10659
rect 28583 10656 28595 10659
rect 28994 10656 29000 10668
rect 28583 10628 29000 10656
rect 28583 10625 28595 10628
rect 28537 10619 28595 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 29733 10659 29791 10665
rect 29733 10625 29745 10659
rect 29779 10625 29791 10659
rect 29733 10619 29791 10625
rect 29748 10588 29776 10619
rect 29822 10616 29828 10668
rect 29880 10656 29886 10668
rect 30377 10659 30435 10665
rect 30377 10656 30389 10659
rect 29880 10628 30389 10656
rect 29880 10616 29886 10628
rect 30377 10625 30389 10628
rect 30423 10625 30435 10659
rect 30377 10619 30435 10625
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 30984 10628 31754 10656
rect 30984 10616 30990 10628
rect 31726 10588 31754 10628
rect 32582 10616 32588 10668
rect 32640 10616 32646 10668
rect 33045 10659 33103 10665
rect 33045 10656 33057 10659
rect 32692 10628 33057 10656
rect 32692 10588 32720 10628
rect 33045 10625 33057 10628
rect 33091 10625 33103 10659
rect 33045 10619 33103 10625
rect 34793 10659 34851 10665
rect 34793 10625 34805 10659
rect 34839 10625 34851 10659
rect 34793 10619 34851 10625
rect 29748 10560 30420 10588
rect 31726 10560 32720 10588
rect 32769 10591 32827 10597
rect 30392 10532 30420 10560
rect 32769 10557 32781 10591
rect 32815 10557 32827 10591
rect 32769 10551 32827 10557
rect 30374 10480 30380 10532
rect 30432 10480 30438 10532
rect 31846 10480 31852 10532
rect 31904 10520 31910 10532
rect 32677 10523 32735 10529
rect 32677 10520 32689 10523
rect 31904 10492 32689 10520
rect 31904 10480 31910 10492
rect 32677 10489 32689 10492
rect 32723 10489 32735 10523
rect 32784 10520 32812 10551
rect 32858 10548 32864 10600
rect 32916 10548 32922 10600
rect 34422 10520 34428 10532
rect 32784 10492 34428 10520
rect 32677 10483 32735 10489
rect 34422 10480 34428 10492
rect 34480 10480 34486 10532
rect 34808 10520 34836 10619
rect 34992 10597 35020 10696
rect 34977 10591 35035 10597
rect 34977 10557 34989 10591
rect 35023 10557 35035 10591
rect 34977 10551 35035 10557
rect 35728 10520 35756 10755
rect 36906 10752 36912 10764
rect 36964 10752 36970 10804
rect 40126 10752 40132 10804
rect 40184 10752 40190 10804
rect 40862 10752 40868 10804
rect 40920 10792 40926 10804
rect 41049 10795 41107 10801
rect 41049 10792 41061 10795
rect 40920 10764 41061 10792
rect 40920 10752 40926 10764
rect 41049 10761 41061 10764
rect 41095 10761 41107 10795
rect 41049 10755 41107 10761
rect 37274 10684 37280 10736
rect 37332 10724 37338 10736
rect 37829 10727 37887 10733
rect 37829 10724 37841 10727
rect 37332 10696 37841 10724
rect 37332 10684 37338 10696
rect 37829 10693 37841 10696
rect 37875 10693 37887 10727
rect 37829 10687 37887 10693
rect 37918 10684 37924 10736
rect 37976 10724 37982 10736
rect 38013 10727 38071 10733
rect 38013 10724 38025 10727
rect 37976 10696 38025 10724
rect 37976 10684 37982 10696
rect 38013 10693 38025 10696
rect 38059 10693 38071 10727
rect 40402 10724 40408 10736
rect 38013 10687 38071 10693
rect 38764 10696 40408 10724
rect 38764 10665 38792 10696
rect 40402 10684 40408 10696
rect 40460 10684 40466 10736
rect 41064 10724 41092 10755
rect 41138 10752 41144 10804
rect 41196 10752 41202 10804
rect 42242 10752 42248 10804
rect 42300 10792 42306 10804
rect 42613 10795 42671 10801
rect 42613 10792 42625 10795
rect 42300 10764 42625 10792
rect 42300 10752 42306 10764
rect 42613 10761 42625 10764
rect 42659 10761 42671 10795
rect 42613 10755 42671 10761
rect 43349 10795 43407 10801
rect 43349 10761 43361 10795
rect 43395 10792 43407 10795
rect 43530 10792 43536 10804
rect 43395 10764 43536 10792
rect 43395 10761 43407 10764
rect 43349 10755 43407 10761
rect 43530 10752 43536 10764
rect 43588 10752 43594 10804
rect 41414 10724 41420 10736
rect 41064 10696 41420 10724
rect 41414 10684 41420 10696
rect 41472 10684 41478 10736
rect 39022 10665 39028 10668
rect 38749 10659 38807 10665
rect 38749 10625 38761 10659
rect 38795 10625 38807 10659
rect 38749 10619 38807 10625
rect 39016 10619 39028 10665
rect 39022 10616 39028 10619
rect 39080 10616 39086 10668
rect 41046 10548 41052 10600
rect 41104 10588 41110 10600
rect 41233 10591 41291 10597
rect 41233 10588 41245 10591
rect 41104 10560 41245 10588
rect 41104 10548 41110 10560
rect 41233 10557 41245 10560
rect 41279 10557 41291 10591
rect 41233 10551 41291 10557
rect 34808 10492 35756 10520
rect 40681 10455 40739 10461
rect 40681 10421 40693 10455
rect 40727 10452 40739 10455
rect 40862 10452 40868 10464
rect 40727 10424 40868 10452
rect 40727 10421 40739 10424
rect 40681 10415 40739 10421
rect 40862 10412 40868 10424
rect 40920 10412 40926 10464
rect 41690 10412 41696 10464
rect 41748 10452 41754 10464
rect 41969 10455 42027 10461
rect 41969 10452 41981 10455
rect 41748 10424 41981 10452
rect 41748 10412 41754 10424
rect 41969 10421 41981 10424
rect 42015 10452 42027 10455
rect 42058 10452 42064 10464
rect 42015 10424 42064 10452
rect 42015 10421 42027 10424
rect 41969 10415 42027 10421
rect 42058 10412 42064 10424
rect 42116 10412 42122 10464
rect 1104 10362 43884 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 43884 10362
rect 1104 10288 43884 10310
rect 30558 10208 30564 10260
rect 30616 10208 30622 10260
rect 30926 10208 30932 10260
rect 30984 10208 30990 10260
rect 37829 10251 37887 10257
rect 37829 10217 37841 10251
rect 37875 10248 37887 10251
rect 38286 10248 38292 10260
rect 37875 10220 38292 10248
rect 37875 10217 37887 10220
rect 37829 10211 37887 10217
rect 38286 10208 38292 10220
rect 38344 10208 38350 10260
rect 39022 10208 39028 10260
rect 39080 10248 39086 10260
rect 39209 10251 39267 10257
rect 39209 10248 39221 10251
rect 39080 10220 39221 10248
rect 39080 10208 39086 10220
rect 39209 10217 39221 10220
rect 39255 10217 39267 10251
rect 39209 10211 39267 10217
rect 40034 10208 40040 10260
rect 40092 10208 40098 10260
rect 40678 10208 40684 10260
rect 40736 10208 40742 10260
rect 42058 10208 42064 10260
rect 42116 10208 42122 10260
rect 31018 10072 31024 10124
rect 31076 10072 31082 10124
rect 42978 10072 42984 10124
rect 43036 10112 43042 10124
rect 43073 10115 43131 10121
rect 43073 10112 43085 10115
rect 43036 10084 43085 10112
rect 43036 10072 43042 10084
rect 43073 10081 43085 10084
rect 43119 10081 43131 10115
rect 43073 10075 43131 10081
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 39390 10004 39396 10056
rect 39448 10004 39454 10056
rect 40862 10004 40868 10056
rect 40920 10004 40926 10056
rect 43349 10047 43407 10053
rect 43349 10013 43361 10047
rect 43395 10044 43407 10047
rect 43990 10044 43996 10056
rect 43395 10016 43996 10044
rect 43395 10013 43407 10016
rect 43349 10007 43407 10013
rect 43990 10004 43996 10016
rect 44048 10004 44054 10056
rect 41417 9911 41475 9917
rect 41417 9877 41429 9911
rect 41463 9908 41475 9911
rect 43254 9908 43260 9920
rect 41463 9880 43260 9908
rect 41463 9877 41475 9880
rect 41417 9871 41475 9877
rect 43254 9868 43260 9880
rect 43312 9868 43318 9920
rect 1104 9818 43884 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 43884 9818
rect 1104 9744 43884 9766
rect 40034 9664 40040 9716
rect 40092 9704 40098 9716
rect 40129 9707 40187 9713
rect 40129 9704 40141 9707
rect 40092 9676 40141 9704
rect 40092 9664 40098 9676
rect 40129 9673 40141 9676
rect 40175 9673 40187 9707
rect 40129 9667 40187 9673
rect 43254 9664 43260 9716
rect 43312 9664 43318 9716
rect 40865 9639 40923 9645
rect 40865 9605 40877 9639
rect 40911 9636 40923 9639
rect 41322 9636 41328 9648
rect 40911 9608 41328 9636
rect 40911 9605 40923 9608
rect 40865 9599 40923 9605
rect 41322 9596 41328 9608
rect 41380 9636 41386 9648
rect 41601 9639 41659 9645
rect 41601 9636 41613 9639
rect 41380 9608 41613 9636
rect 41380 9596 41386 9608
rect 41601 9605 41613 9608
rect 41647 9605 41659 9639
rect 41601 9599 41659 9605
rect 42794 9596 42800 9648
rect 42852 9596 42858 9648
rect 40034 9324 40040 9376
rect 40092 9364 40098 9376
rect 42978 9364 42984 9376
rect 40092 9336 42984 9364
rect 40092 9324 40098 9336
rect 42978 9324 42984 9336
rect 43036 9324 43042 9376
rect 1104 9274 43884 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 43884 9274
rect 1104 9200 43884 9222
rect 41414 9120 41420 9172
rect 41472 9160 41478 9172
rect 41877 9163 41935 9169
rect 41877 9160 41889 9163
rect 41472 9132 41889 9160
rect 41472 9120 41478 9132
rect 41877 9129 41889 9132
rect 41923 9160 41935 9163
rect 43070 9160 43076 9172
rect 41923 9132 43076 9160
rect 41923 9129 41935 9132
rect 41877 9123 41935 9129
rect 43070 9120 43076 9132
rect 43128 9120 43134 9172
rect 43346 9120 43352 9172
rect 43404 9120 43410 9172
rect 42797 9095 42855 9101
rect 42797 9061 42809 9095
rect 42843 9092 42855 9095
rect 43364 9092 43392 9120
rect 42843 9064 43392 9092
rect 42843 9061 42855 9064
rect 42797 9055 42855 9061
rect 1104 8730 43884 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 43884 8730
rect 1104 8656 43884 8678
rect 42797 8619 42855 8625
rect 42797 8585 42809 8619
rect 42843 8616 42855 8619
rect 42886 8616 42892 8628
rect 42843 8588 42892 8616
rect 42843 8585 42855 8588
rect 42797 8579 42855 8585
rect 42886 8576 42892 8588
rect 42944 8616 42950 8628
rect 43257 8619 43315 8625
rect 43257 8616 43269 8619
rect 42944 8588 43269 8616
rect 42944 8576 42950 8588
rect 43257 8585 43269 8588
rect 43303 8585 43315 8619
rect 43257 8579 43315 8585
rect 1104 8186 43884 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 43884 8186
rect 1104 8112 43884 8134
rect 43349 8075 43407 8081
rect 43349 8041 43361 8075
rect 43395 8072 43407 8075
rect 43990 8072 43996 8084
rect 43395 8044 43996 8072
rect 43395 8041 43407 8044
rect 43349 8035 43407 8041
rect 43990 8032 43996 8044
rect 44048 8032 44054 8084
rect 1104 7642 43884 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 43884 7642
rect 1104 7568 43884 7590
rect 1104 7098 43884 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 43884 7098
rect 1104 7024 43884 7046
rect 1104 6554 43884 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 43884 6554
rect 1104 6480 43884 6502
rect 43070 6332 43076 6384
rect 43128 6332 43134 6384
rect 43346 6264 43352 6316
rect 43404 6264 43410 6316
rect 1104 6010 43884 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 43884 6010
rect 1104 5936 43884 5958
rect 43346 5856 43352 5908
rect 43404 5856 43410 5908
rect 1104 5466 43884 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 43884 5466
rect 1104 5392 43884 5414
rect 1104 4922 43884 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 43884 4922
rect 1104 4848 43884 4870
rect 1104 4378 43884 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 43884 4378
rect 1104 4304 43884 4326
rect 1104 3834 43884 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 43884 3834
rect 1104 3760 43884 3782
rect 1104 3290 43884 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 43884 3290
rect 1104 3216 43884 3238
rect 43346 2796 43352 2848
rect 43404 2796 43410 2848
rect 1104 2746 43884 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 43884 2746
rect 1104 2672 43884 2694
rect 42978 2456 42984 2508
rect 43036 2496 43042 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 43036 2468 43085 2496
rect 43036 2456 43042 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 43346 2388 43352 2440
rect 43404 2428 43410 2440
rect 43990 2428 43996 2440
rect 43404 2400 43996 2428
rect 43404 2388 43410 2400
rect 43990 2388 43996 2400
rect 44048 2388 44054 2440
rect 1104 2202 43884 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 43884 2202
rect 1104 2128 43884 2150
<< via1 >>
rect 29460 44072 29512 44124
rect 31760 44072 31812 44124
rect 34152 44072 34204 44124
rect 34612 44072 34664 44124
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 27068 42304 27120 42356
rect 27528 42236 27580 42288
rect 37924 42304 37976 42356
rect 13820 42168 13872 42220
rect 15384 42168 15436 42220
rect 20720 42168 20772 42220
rect 22744 42211 22796 42220
rect 22744 42177 22753 42211
rect 22753 42177 22787 42211
rect 22787 42177 22796 42211
rect 22744 42168 22796 42177
rect 25412 42211 25464 42220
rect 25412 42177 25421 42211
rect 25421 42177 25455 42211
rect 25455 42177 25464 42211
rect 25412 42168 25464 42177
rect 27344 42211 27396 42220
rect 27344 42177 27353 42211
rect 27353 42177 27387 42211
rect 27387 42177 27396 42211
rect 27344 42168 27396 42177
rect 27436 42168 27488 42220
rect 30656 42211 30708 42220
rect 30656 42177 30665 42211
rect 30665 42177 30699 42211
rect 30699 42177 30708 42211
rect 30656 42168 30708 42177
rect 32312 42211 32364 42220
rect 32312 42177 32321 42211
rect 32321 42177 32355 42211
rect 32355 42177 32364 42211
rect 32312 42168 32364 42177
rect 34796 42168 34848 42220
rect 37556 42236 37608 42288
rect 38384 42168 38436 42220
rect 21456 42075 21508 42084
rect 21456 42041 21465 42075
rect 21465 42041 21499 42075
rect 21499 42041 21508 42075
rect 21456 42032 21508 42041
rect 29644 42032 29696 42084
rect 31576 42032 31628 42084
rect 34336 42100 34388 42152
rect 38200 42100 38252 42152
rect 43996 42168 44048 42220
rect 42800 42100 42852 42152
rect 39304 42032 39356 42084
rect 20444 42007 20496 42016
rect 20444 41973 20453 42007
rect 20453 41973 20487 42007
rect 20487 41973 20496 42007
rect 20444 41964 20496 41973
rect 22100 42007 22152 42016
rect 22100 41973 22109 42007
rect 22109 41973 22143 42007
rect 22143 41973 22152 42007
rect 22100 41964 22152 41973
rect 22560 42007 22612 42016
rect 22560 41973 22569 42007
rect 22569 41973 22603 42007
rect 22603 41973 22612 42007
rect 22560 41964 22612 41973
rect 23388 42007 23440 42016
rect 23388 41973 23397 42007
rect 23397 41973 23431 42007
rect 23431 41973 23440 42007
rect 23388 41964 23440 41973
rect 25044 41964 25096 42016
rect 25228 42007 25280 42016
rect 25228 41973 25237 42007
rect 25237 41973 25271 42007
rect 25271 41973 25280 42007
rect 25228 41964 25280 41973
rect 26608 41964 26660 42016
rect 27068 41964 27120 42016
rect 27160 42007 27212 42016
rect 27160 41973 27169 42007
rect 27169 41973 27203 42007
rect 27203 41973 27212 42007
rect 27160 41964 27212 41973
rect 29000 41964 29052 42016
rect 30840 42007 30892 42016
rect 30840 41973 30849 42007
rect 30849 41973 30883 42007
rect 30883 41973 30892 42007
rect 30840 41964 30892 41973
rect 32588 41964 32640 42016
rect 33600 41964 33652 42016
rect 34244 42007 34296 42016
rect 34244 41973 34253 42007
rect 34253 41973 34287 42007
rect 34287 41973 34296 42007
rect 34244 41964 34296 41973
rect 35440 41964 35492 42016
rect 36084 42007 36136 42016
rect 36084 41973 36093 42007
rect 36093 41973 36127 42007
rect 36127 41973 36136 42007
rect 36084 41964 36136 41973
rect 36176 41964 36228 42016
rect 38384 41964 38436 42016
rect 38936 41964 38988 42016
rect 40500 41964 40552 42016
rect 40592 42007 40644 42016
rect 40592 41973 40601 42007
rect 40601 41973 40635 42007
rect 40635 41973 40644 42007
rect 40592 41964 40644 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 31484 41760 31536 41812
rect 37556 41760 37608 41812
rect 41972 41760 42024 41812
rect 39396 41692 39448 41744
rect 29644 41624 29696 41676
rect 31576 41667 31628 41676
rect 31576 41633 31585 41667
rect 31585 41633 31619 41667
rect 31619 41633 31628 41667
rect 31576 41624 31628 41633
rect 40132 41667 40184 41676
rect 40132 41633 40141 41667
rect 40141 41633 40175 41667
rect 40175 41633 40184 41667
rect 40132 41624 40184 41633
rect 20076 41556 20128 41608
rect 22560 41599 22612 41608
rect 22560 41565 22594 41599
rect 22594 41565 22612 41599
rect 22560 41556 22612 41565
rect 24952 41556 25004 41608
rect 26884 41599 26936 41608
rect 20444 41488 20496 41540
rect 21364 41463 21416 41472
rect 21364 41429 21373 41463
rect 21373 41429 21407 41463
rect 21407 41429 21416 41463
rect 21364 41420 21416 41429
rect 24124 41420 24176 41472
rect 25228 41488 25280 41540
rect 26884 41565 26893 41599
rect 26893 41565 26927 41599
rect 26927 41565 26936 41599
rect 26884 41556 26936 41565
rect 27160 41599 27212 41608
rect 27160 41565 27194 41599
rect 27194 41565 27212 41599
rect 27160 41556 27212 41565
rect 29092 41556 29144 41608
rect 30840 41556 30892 41608
rect 35440 41556 35492 41608
rect 36728 41556 36780 41608
rect 36912 41599 36964 41608
rect 36912 41565 36921 41599
rect 36921 41565 36955 41599
rect 36955 41565 36964 41599
rect 36912 41556 36964 41565
rect 37464 41599 37516 41608
rect 37464 41565 37473 41599
rect 37473 41565 37507 41599
rect 37507 41565 37516 41599
rect 37464 41556 37516 41565
rect 38660 41599 38712 41608
rect 38660 41565 38669 41599
rect 38669 41565 38703 41599
rect 38703 41565 38712 41599
rect 38660 41556 38712 41565
rect 42156 41599 42208 41608
rect 42156 41565 42165 41599
rect 42165 41565 42199 41599
rect 42199 41565 42208 41599
rect 42156 41556 42208 41565
rect 43536 41556 43588 41608
rect 26700 41420 26752 41472
rect 28264 41463 28316 41472
rect 28264 41429 28273 41463
rect 28273 41429 28307 41463
rect 28307 41429 28316 41463
rect 28264 41420 28316 41429
rect 33508 41531 33560 41540
rect 33508 41497 33517 41531
rect 33517 41497 33551 41531
rect 33551 41497 33560 41531
rect 33508 41488 33560 41497
rect 33876 41531 33928 41540
rect 33876 41497 33885 41531
rect 33885 41497 33919 41531
rect 33919 41497 33928 41531
rect 33876 41488 33928 41497
rect 40592 41488 40644 41540
rect 43076 41488 43128 41540
rect 30932 41420 30984 41472
rect 31852 41420 31904 41472
rect 32496 41420 32548 41472
rect 34704 41420 34756 41472
rect 36268 41420 36320 41472
rect 37740 41420 37792 41472
rect 38384 41420 38436 41472
rect 39304 41463 39356 41472
rect 39304 41429 39313 41463
rect 39313 41429 39347 41463
rect 39347 41429 39356 41463
rect 39304 41420 39356 41429
rect 39672 41420 39724 41472
rect 40316 41463 40368 41472
rect 40316 41429 40325 41463
rect 40325 41429 40359 41463
rect 40359 41429 40368 41463
rect 40316 41420 40368 41429
rect 40408 41463 40460 41472
rect 40408 41429 40417 41463
rect 40417 41429 40451 41463
rect 40451 41429 40460 41463
rect 40408 41420 40460 41429
rect 41144 41420 41196 41472
rect 41236 41463 41288 41472
rect 41236 41429 41245 41463
rect 41245 41429 41279 41463
rect 41279 41429 41288 41463
rect 41236 41420 41288 41429
rect 42616 41463 42668 41472
rect 42616 41429 42625 41463
rect 42625 41429 42659 41463
rect 42659 41429 42668 41463
rect 42616 41420 42668 41429
rect 42892 41420 42944 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 21456 41216 21508 41268
rect 22744 41216 22796 41268
rect 25412 41216 25464 41268
rect 27344 41216 27396 41268
rect 28264 41216 28316 41268
rect 29092 41259 29144 41268
rect 29092 41225 29101 41259
rect 29101 41225 29135 41259
rect 29135 41225 29144 41259
rect 29092 41216 29144 41225
rect 30656 41259 30708 41268
rect 30656 41225 30665 41259
rect 30665 41225 30699 41259
rect 30699 41225 30708 41259
rect 30656 41216 30708 41225
rect 32864 41216 32916 41268
rect 34796 41216 34848 41268
rect 39948 41216 40000 41268
rect 42892 41216 42944 41268
rect 43076 41216 43128 41268
rect 21364 41148 21416 41200
rect 21548 41148 21600 41200
rect 31852 41148 31904 41200
rect 21640 41080 21692 41132
rect 21824 41080 21876 41132
rect 24124 41080 24176 41132
rect 26700 41080 26752 41132
rect 27896 41080 27948 41132
rect 30472 41080 30524 41132
rect 30932 41080 30984 41132
rect 31668 41080 31720 41132
rect 39304 41148 39356 41200
rect 39396 41148 39448 41200
rect 32588 41123 32640 41132
rect 32588 41089 32622 41123
rect 32622 41089 32640 41123
rect 32588 41080 32640 41089
rect 34704 41123 34756 41132
rect 34704 41089 34713 41123
rect 34713 41089 34747 41123
rect 34747 41089 34756 41123
rect 34704 41080 34756 41089
rect 36268 41080 36320 41132
rect 37740 41123 37792 41132
rect 37740 41089 37774 41123
rect 37774 41089 37792 41123
rect 37740 41080 37792 41089
rect 41144 41123 41196 41132
rect 41144 41089 41153 41123
rect 41153 41089 41187 41123
rect 41187 41089 41196 41123
rect 41144 41080 41196 41089
rect 18880 41012 18932 41064
rect 23296 41055 23348 41064
rect 23296 41021 23305 41055
rect 23305 41021 23339 41055
rect 23339 41021 23348 41055
rect 23296 41012 23348 41021
rect 23388 41012 23440 41064
rect 20720 40987 20772 40996
rect 20720 40953 20729 40987
rect 20729 40953 20763 40987
rect 20763 40953 20772 40987
rect 20720 40944 20772 40953
rect 22100 40944 22152 40996
rect 24860 41012 24912 41064
rect 25780 41055 25832 41064
rect 25780 41021 25789 41055
rect 25789 41021 25823 41055
rect 25823 41021 25832 41055
rect 25780 41012 25832 41021
rect 26332 41012 26384 41064
rect 27620 41055 27672 41064
rect 27620 41021 27629 41055
rect 27629 41021 27663 41055
rect 27663 41021 27672 41055
rect 27620 41012 27672 41021
rect 28540 41012 28592 41064
rect 30288 41012 30340 41064
rect 31116 41055 31168 41064
rect 31116 41021 31125 41055
rect 31125 41021 31159 41055
rect 31159 41021 31168 41055
rect 31116 41012 31168 41021
rect 33508 41012 33560 41064
rect 34428 41055 34480 41064
rect 34428 41021 34437 41055
rect 34437 41021 34471 41055
rect 34471 41021 34480 41055
rect 34428 41012 34480 41021
rect 34612 41055 34664 41064
rect 34612 41021 34621 41055
rect 34621 41021 34655 41055
rect 34655 41021 34664 41055
rect 34612 41012 34664 41021
rect 34796 41012 34848 41064
rect 22652 40876 22704 40928
rect 25228 40876 25280 40928
rect 26608 40919 26660 40928
rect 26608 40885 26617 40919
rect 26617 40885 26651 40919
rect 26651 40885 26660 40919
rect 26608 40876 26660 40885
rect 26976 40876 27028 40928
rect 30104 40919 30156 40928
rect 30104 40885 30113 40919
rect 30113 40885 30147 40919
rect 30147 40885 30156 40919
rect 30104 40876 30156 40885
rect 31576 40876 31628 40928
rect 33876 40944 33928 40996
rect 34060 40944 34112 40996
rect 37004 40876 37056 40928
rect 38844 41012 38896 41064
rect 38752 40876 38804 40928
rect 41420 40944 41472 40996
rect 41328 40919 41380 40928
rect 41328 40885 41337 40919
rect 41337 40885 41371 40919
rect 41371 40885 41380 40919
rect 41328 40876 41380 40885
rect 41788 40919 41840 40928
rect 41788 40885 41797 40919
rect 41797 40885 41831 40919
rect 41831 40885 41840 40919
rect 41788 40876 41840 40885
rect 42616 40919 42668 40928
rect 42616 40885 42625 40919
rect 42625 40885 42659 40919
rect 42659 40885 42668 40919
rect 42616 40876 42668 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 24308 40672 24360 40724
rect 32312 40672 32364 40724
rect 30288 40604 30340 40656
rect 34244 40672 34296 40724
rect 34428 40672 34480 40724
rect 22928 40536 22980 40588
rect 24952 40536 25004 40588
rect 31576 40579 31628 40588
rect 31576 40545 31585 40579
rect 31585 40545 31619 40579
rect 31619 40545 31628 40579
rect 31576 40536 31628 40545
rect 36912 40715 36964 40724
rect 36912 40681 36921 40715
rect 36921 40681 36955 40715
rect 36955 40681 36964 40715
rect 36912 40672 36964 40681
rect 37464 40672 37516 40724
rect 38660 40672 38712 40724
rect 38384 40604 38436 40656
rect 40408 40672 40460 40724
rect 40132 40536 40184 40588
rect 20628 40511 20680 40520
rect 20628 40477 20637 40511
rect 20637 40477 20671 40511
rect 20671 40477 20680 40511
rect 20628 40468 20680 40477
rect 25044 40511 25096 40520
rect 25044 40477 25053 40511
rect 25053 40477 25087 40511
rect 25087 40477 25096 40511
rect 25044 40468 25096 40477
rect 27712 40468 27764 40520
rect 31484 40468 31536 40520
rect 32864 40468 32916 40520
rect 34060 40511 34112 40520
rect 34060 40477 34069 40511
rect 34069 40477 34103 40511
rect 34103 40477 34112 40511
rect 34060 40468 34112 40477
rect 35716 40511 35768 40520
rect 35716 40477 35725 40511
rect 35725 40477 35759 40511
rect 35759 40477 35768 40511
rect 35716 40468 35768 40477
rect 37004 40468 37056 40520
rect 37740 40468 37792 40520
rect 37924 40468 37976 40520
rect 23572 40400 23624 40452
rect 24860 40400 24912 40452
rect 25964 40400 26016 40452
rect 26240 40400 26292 40452
rect 28356 40400 28408 40452
rect 28908 40443 28960 40452
rect 28908 40409 28917 40443
rect 28917 40409 28951 40443
rect 28951 40409 28960 40443
rect 28908 40400 28960 40409
rect 30656 40400 30708 40452
rect 31760 40443 31812 40452
rect 31760 40409 31769 40443
rect 31769 40409 31803 40443
rect 31803 40409 31812 40443
rect 31760 40400 31812 40409
rect 32772 40400 32824 40452
rect 33140 40400 33192 40452
rect 18788 40375 18840 40384
rect 18788 40341 18797 40375
rect 18797 40341 18831 40375
rect 18831 40341 18840 40375
rect 18788 40332 18840 40341
rect 21088 40332 21140 40384
rect 21272 40332 21324 40384
rect 22560 40332 22612 40384
rect 22744 40332 22796 40384
rect 26332 40332 26384 40384
rect 27896 40332 27948 40384
rect 29828 40375 29880 40384
rect 29828 40341 29837 40375
rect 29837 40341 29871 40375
rect 29871 40341 29880 40375
rect 29828 40332 29880 40341
rect 30380 40375 30432 40384
rect 30380 40341 30389 40375
rect 30389 40341 30423 40375
rect 30423 40341 30432 40375
rect 30380 40332 30432 40341
rect 33232 40332 33284 40384
rect 33968 40400 34020 40452
rect 34336 40400 34388 40452
rect 37188 40400 37240 40452
rect 37464 40400 37516 40452
rect 39948 40400 40000 40452
rect 35900 40332 35952 40384
rect 36452 40375 36504 40384
rect 36452 40341 36461 40375
rect 36461 40341 36495 40375
rect 36495 40341 36504 40375
rect 36452 40332 36504 40341
rect 38752 40332 38804 40384
rect 38936 40375 38988 40384
rect 38936 40341 38945 40375
rect 38945 40341 38979 40375
rect 38979 40341 38988 40375
rect 38936 40332 38988 40341
rect 39028 40375 39080 40384
rect 39028 40341 39037 40375
rect 39037 40341 39071 40375
rect 39071 40341 39080 40375
rect 39028 40332 39080 40341
rect 39488 40332 39540 40384
rect 41328 40468 41380 40520
rect 41420 40511 41472 40520
rect 41420 40477 41429 40511
rect 41429 40477 41463 40511
rect 41463 40477 41472 40511
rect 41420 40468 41472 40477
rect 41880 40468 41932 40520
rect 42616 40400 42668 40452
rect 41604 40332 41656 40384
rect 42340 40332 42392 40384
rect 42892 40332 42944 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 9128 40060 9180 40112
rect 9680 40060 9732 40112
rect 16948 40060 17000 40112
rect 19156 40060 19208 40112
rect 18328 39992 18380 40044
rect 20628 40060 20680 40112
rect 19892 39992 19944 40044
rect 22376 40128 22428 40180
rect 22652 39992 22704 40044
rect 23112 40128 23164 40180
rect 25044 40060 25096 40112
rect 29184 40128 29236 40180
rect 30104 40128 30156 40180
rect 20076 39967 20128 39976
rect 20076 39933 20085 39967
rect 20085 39933 20119 39967
rect 20119 39933 20128 39967
rect 20076 39924 20128 39933
rect 21180 39856 21232 39908
rect 23572 39924 23624 39976
rect 23756 39967 23808 39976
rect 23756 39933 23765 39967
rect 23765 39933 23799 39967
rect 23799 39933 23808 39967
rect 23756 39924 23808 39933
rect 24584 39967 24636 39976
rect 24584 39933 24593 39967
rect 24593 39933 24627 39967
rect 24627 39933 24636 39967
rect 24584 39924 24636 39933
rect 20720 39788 20772 39840
rect 22652 39788 22704 39840
rect 24216 39856 24268 39908
rect 24860 39967 24912 39976
rect 24860 39933 24869 39967
rect 24869 39933 24903 39967
rect 24903 39933 24912 39967
rect 24860 39924 24912 39933
rect 27804 39992 27856 40044
rect 28724 40035 28776 40044
rect 28724 40001 28758 40035
rect 28758 40001 28776 40035
rect 28724 39992 28776 40001
rect 30196 40060 30248 40112
rect 31852 40060 31904 40112
rect 33968 40128 34020 40180
rect 34152 40128 34204 40180
rect 37096 40128 37148 40180
rect 37924 40128 37976 40180
rect 41328 40171 41380 40180
rect 41328 40137 41337 40171
rect 41337 40137 41371 40171
rect 41371 40137 41380 40171
rect 41328 40128 41380 40137
rect 30380 39992 30432 40044
rect 26884 39924 26936 39976
rect 27160 39924 27212 39976
rect 31024 39992 31076 40044
rect 31760 40035 31812 40044
rect 31760 40001 31769 40035
rect 31769 40001 31803 40035
rect 31803 40001 31812 40035
rect 31760 39992 31812 40001
rect 32680 39992 32732 40044
rect 33232 40035 33284 40044
rect 33232 40001 33241 40035
rect 33241 40001 33275 40035
rect 33275 40001 33284 40035
rect 33232 39992 33284 40001
rect 33784 39992 33836 40044
rect 35440 39992 35492 40044
rect 36636 39992 36688 40044
rect 38476 39992 38528 40044
rect 31392 39924 31444 39976
rect 33508 39924 33560 39976
rect 36728 39967 36780 39976
rect 36728 39933 36737 39967
rect 36737 39933 36771 39967
rect 36771 39933 36780 39967
rect 36728 39924 36780 39933
rect 38844 39924 38896 39976
rect 32404 39899 32456 39908
rect 32404 39865 32413 39899
rect 32413 39865 32447 39899
rect 32447 39865 32456 39899
rect 41236 39924 41288 39976
rect 32404 39856 32456 39865
rect 25044 39788 25096 39840
rect 27068 39788 27120 39840
rect 27528 39788 27580 39840
rect 27712 39831 27764 39840
rect 27712 39797 27721 39831
rect 27721 39797 27755 39831
rect 27755 39797 27764 39831
rect 27712 39788 27764 39797
rect 29092 39788 29144 39840
rect 30840 39788 30892 39840
rect 31576 39831 31628 39840
rect 31576 39797 31585 39831
rect 31585 39797 31619 39831
rect 31619 39797 31628 39831
rect 31576 39788 31628 39797
rect 34612 39788 34664 39840
rect 37556 39831 37608 39840
rect 37556 39797 37565 39831
rect 37565 39797 37599 39831
rect 37599 39797 37608 39831
rect 37556 39788 37608 39797
rect 38108 39788 38160 39840
rect 42708 39856 42760 39908
rect 39304 39788 39356 39840
rect 39396 39788 39448 39840
rect 42616 39831 42668 39840
rect 42616 39797 42625 39831
rect 42625 39797 42659 39831
rect 42659 39797 42668 39831
rect 42616 39788 42668 39797
rect 43444 39788 43496 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 16120 39584 16172 39636
rect 18328 39627 18380 39636
rect 18328 39593 18337 39627
rect 18337 39593 18371 39627
rect 18371 39593 18380 39627
rect 18328 39584 18380 39593
rect 18880 39627 18932 39636
rect 18880 39593 18889 39627
rect 18889 39593 18923 39627
rect 18923 39593 18932 39627
rect 18880 39584 18932 39593
rect 20628 39584 20680 39636
rect 23112 39627 23164 39636
rect 23112 39593 23121 39627
rect 23121 39593 23155 39627
rect 23155 39593 23164 39627
rect 23112 39584 23164 39593
rect 20812 39516 20864 39568
rect 22192 39516 22244 39568
rect 28724 39584 28776 39636
rect 36084 39627 36136 39636
rect 36084 39593 36118 39627
rect 36118 39593 36136 39627
rect 36084 39584 36136 39593
rect 29736 39516 29788 39568
rect 33692 39516 33744 39568
rect 35440 39559 35492 39568
rect 35440 39525 35449 39559
rect 35449 39525 35483 39559
rect 35483 39525 35492 39559
rect 35440 39516 35492 39525
rect 36912 39516 36964 39568
rect 37188 39516 37240 39568
rect 41328 39584 41380 39636
rect 18788 39380 18840 39432
rect 19432 39380 19484 39432
rect 20720 39380 20772 39432
rect 21088 39380 21140 39432
rect 22928 39380 22980 39432
rect 24952 39448 25004 39500
rect 26516 39491 26568 39500
rect 26516 39457 26525 39491
rect 26525 39457 26559 39491
rect 26559 39457 26568 39491
rect 26516 39448 26568 39457
rect 26792 39491 26844 39500
rect 26792 39457 26801 39491
rect 26801 39457 26835 39491
rect 26835 39457 26844 39491
rect 26792 39448 26844 39457
rect 28356 39491 28408 39500
rect 28356 39457 28365 39491
rect 28365 39457 28399 39491
rect 28399 39457 28408 39491
rect 28356 39448 28408 39457
rect 30288 39448 30340 39500
rect 31760 39448 31812 39500
rect 23664 39423 23716 39432
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 24584 39380 24636 39432
rect 25044 39423 25096 39432
rect 25044 39389 25053 39423
rect 25053 39389 25087 39423
rect 25087 39389 25096 39423
rect 25044 39380 25096 39389
rect 28908 39380 28960 39432
rect 31576 39380 31628 39432
rect 31668 39423 31720 39432
rect 31668 39389 31677 39423
rect 31677 39389 31711 39423
rect 31711 39389 31720 39423
rect 31668 39380 31720 39389
rect 32864 39423 32916 39432
rect 32864 39389 32873 39423
rect 32873 39389 32907 39423
rect 32907 39389 32916 39423
rect 32864 39380 32916 39389
rect 34520 39380 34572 39432
rect 35348 39448 35400 39500
rect 36084 39448 36136 39500
rect 40040 39516 40092 39568
rect 18880 39244 18932 39296
rect 20536 39355 20588 39364
rect 20536 39321 20545 39355
rect 20545 39321 20579 39355
rect 20579 39321 20588 39355
rect 20536 39312 20588 39321
rect 22192 39312 22244 39364
rect 22928 39244 22980 39296
rect 25044 39244 25096 39296
rect 26516 39312 26568 39364
rect 29644 39312 29696 39364
rect 32588 39312 32640 39364
rect 38016 39423 38068 39432
rect 38016 39389 38025 39423
rect 38025 39389 38059 39423
rect 38059 39389 38068 39423
rect 38016 39380 38068 39389
rect 39120 39423 39172 39432
rect 29000 39244 29052 39296
rect 29460 39244 29512 39296
rect 30196 39244 30248 39296
rect 33232 39244 33284 39296
rect 33324 39244 33376 39296
rect 33600 39244 33652 39296
rect 33876 39244 33928 39296
rect 35992 39244 36044 39296
rect 36084 39287 36136 39296
rect 36084 39253 36109 39287
rect 36109 39253 36136 39287
rect 39120 39389 39129 39423
rect 39129 39389 39163 39423
rect 39163 39389 39172 39423
rect 39120 39380 39172 39389
rect 36084 39244 36136 39253
rect 36268 39287 36320 39296
rect 36268 39253 36277 39287
rect 36277 39253 36311 39287
rect 36311 39253 36320 39287
rect 38844 39312 38896 39364
rect 41880 39423 41932 39432
rect 41880 39389 41889 39423
rect 41889 39389 41923 39423
rect 41923 39389 41932 39423
rect 41880 39380 41932 39389
rect 40408 39312 40460 39364
rect 41144 39312 41196 39364
rect 36268 39244 36320 39253
rect 38568 39244 38620 39296
rect 39304 39244 39356 39296
rect 40316 39244 40368 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 19984 39040 20036 39092
rect 23664 39040 23716 39092
rect 18880 38972 18932 39024
rect 20812 39015 20864 39024
rect 20812 38981 20821 39015
rect 20821 38981 20855 39015
rect 20855 38981 20864 39015
rect 20812 38972 20864 38981
rect 22468 38972 22520 39024
rect 22744 38972 22796 39024
rect 24492 39040 24544 39092
rect 24584 39040 24636 39092
rect 29644 39040 29696 39092
rect 31024 39083 31076 39092
rect 31024 39049 31033 39083
rect 31033 39049 31067 39083
rect 31067 39049 31076 39083
rect 31024 39040 31076 39049
rect 31760 39040 31812 39092
rect 32588 39040 32640 39092
rect 16580 38904 16632 38956
rect 21180 38904 21232 38956
rect 22100 38904 22152 38956
rect 22560 38947 22612 38956
rect 18052 38836 18104 38888
rect 22560 38913 22568 38947
rect 22568 38913 22602 38947
rect 22602 38913 22612 38947
rect 22560 38904 22612 38913
rect 22652 38947 22704 38956
rect 22652 38913 22661 38947
rect 22661 38913 22695 38947
rect 22695 38913 22704 38947
rect 22652 38904 22704 38913
rect 24400 38947 24452 38956
rect 24400 38913 24409 38947
rect 24409 38913 24443 38947
rect 24443 38913 24452 38947
rect 24400 38904 24452 38913
rect 16948 38811 17000 38820
rect 16948 38777 16957 38811
rect 16957 38777 16991 38811
rect 16991 38777 17000 38811
rect 16948 38768 17000 38777
rect 19800 38768 19852 38820
rect 20536 38811 20588 38820
rect 20536 38777 20545 38811
rect 20545 38777 20579 38811
rect 20579 38777 20588 38811
rect 20536 38768 20588 38777
rect 20996 38768 21048 38820
rect 24216 38768 24268 38820
rect 24860 38768 24912 38820
rect 26792 38972 26844 39024
rect 27528 38972 27580 39024
rect 29828 38972 29880 39024
rect 30564 38972 30616 39024
rect 25136 38947 25188 38956
rect 25136 38913 25145 38947
rect 25145 38913 25179 38947
rect 25179 38913 25188 38947
rect 25136 38904 25188 38913
rect 28632 38904 28684 38956
rect 29092 38904 29144 38956
rect 26792 38836 26844 38888
rect 27160 38879 27212 38888
rect 27160 38845 27169 38879
rect 27169 38845 27203 38879
rect 27203 38845 27212 38879
rect 27160 38836 27212 38845
rect 30656 38947 30708 38956
rect 30656 38913 30665 38947
rect 30665 38913 30699 38947
rect 30699 38913 30708 38947
rect 30656 38904 30708 38913
rect 30840 38947 30892 38956
rect 30840 38913 30849 38947
rect 30849 38913 30883 38947
rect 30883 38913 30892 38947
rect 30840 38904 30892 38913
rect 32680 38972 32732 39024
rect 33600 38947 33652 38956
rect 33600 38913 33609 38947
rect 33609 38913 33643 38947
rect 33643 38913 33652 38947
rect 33600 38904 33652 38913
rect 33232 38836 33284 38888
rect 25320 38768 25372 38820
rect 26332 38768 26384 38820
rect 28356 38768 28408 38820
rect 29276 38768 29328 38820
rect 31392 38768 31444 38820
rect 31760 38768 31812 38820
rect 20260 38700 20312 38752
rect 21364 38743 21416 38752
rect 21364 38709 21373 38743
rect 21373 38709 21407 38743
rect 21407 38709 21416 38743
rect 21364 38700 21416 38709
rect 23388 38700 23440 38752
rect 25596 38743 25648 38752
rect 25596 38709 25605 38743
rect 25605 38709 25639 38743
rect 25639 38709 25648 38743
rect 25596 38700 25648 38709
rect 26424 38743 26476 38752
rect 26424 38709 26433 38743
rect 26433 38709 26467 38743
rect 26467 38709 26476 38743
rect 26424 38700 26476 38709
rect 28448 38700 28500 38752
rect 28908 38700 28960 38752
rect 32864 38768 32916 38820
rect 33140 38768 33192 38820
rect 34796 39015 34848 39024
rect 34796 38981 34805 39015
rect 34805 38981 34839 39015
rect 34839 38981 34848 39015
rect 34796 38972 34848 38981
rect 34244 38947 34296 38956
rect 34244 38913 34253 38947
rect 34253 38913 34287 38947
rect 34287 38913 34296 38947
rect 34244 38904 34296 38913
rect 34428 38904 34480 38956
rect 35532 38947 35584 38956
rect 35532 38913 35541 38947
rect 35541 38913 35575 38947
rect 35575 38913 35584 38947
rect 35532 38904 35584 38913
rect 35624 38947 35676 38956
rect 35624 38913 35633 38947
rect 35633 38913 35667 38947
rect 35667 38913 35676 38947
rect 35624 38904 35676 38913
rect 37648 39040 37700 39092
rect 39304 39083 39356 39092
rect 39304 39049 39313 39083
rect 39313 39049 39347 39083
rect 39347 39049 39356 39083
rect 39304 39040 39356 39049
rect 41144 39083 41196 39092
rect 41144 39049 41153 39083
rect 41153 39049 41187 39083
rect 41187 39049 41196 39083
rect 41144 39040 41196 39049
rect 42616 39040 42668 39092
rect 35992 38972 36044 39024
rect 34704 38836 34756 38888
rect 35440 38836 35492 38888
rect 39120 38972 39172 39024
rect 40132 38972 40184 39024
rect 40684 38972 40736 39024
rect 36268 38904 36320 38956
rect 36912 38947 36964 38956
rect 36912 38913 36921 38947
rect 36921 38913 36955 38947
rect 36955 38913 36964 38947
rect 36912 38904 36964 38913
rect 40868 38904 40920 38956
rect 41052 38947 41104 38956
rect 41052 38913 41061 38947
rect 41061 38913 41095 38947
rect 41095 38913 41104 38947
rect 41052 38904 41104 38913
rect 38844 38879 38896 38888
rect 38844 38845 38853 38879
rect 38853 38845 38887 38879
rect 38887 38845 38896 38879
rect 38844 38836 38896 38845
rect 33784 38700 33836 38752
rect 34244 38700 34296 38752
rect 37280 38700 37332 38752
rect 40316 38768 40368 38820
rect 41144 38836 41196 38888
rect 40868 38768 40920 38820
rect 40040 38700 40092 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 18788 38496 18840 38548
rect 19432 38539 19484 38548
rect 19432 38505 19441 38539
rect 19441 38505 19475 38539
rect 19475 38505 19484 38539
rect 19432 38496 19484 38505
rect 21456 38496 21508 38548
rect 21640 38496 21692 38548
rect 22100 38496 22152 38548
rect 22468 38496 22520 38548
rect 23112 38496 23164 38548
rect 24400 38496 24452 38548
rect 24676 38496 24728 38548
rect 18972 38360 19024 38412
rect 19432 38360 19484 38412
rect 17500 38335 17552 38344
rect 17500 38301 17509 38335
rect 17509 38301 17543 38335
rect 17543 38301 17552 38335
rect 17500 38292 17552 38301
rect 18052 38292 18104 38344
rect 19800 38335 19852 38344
rect 19800 38301 19809 38335
rect 19809 38301 19843 38335
rect 19843 38301 19852 38335
rect 19800 38292 19852 38301
rect 20168 38292 20220 38344
rect 18236 38224 18288 38276
rect 14464 38156 14516 38208
rect 19248 38156 19300 38208
rect 20812 38335 20864 38344
rect 20812 38301 20822 38335
rect 20822 38301 20856 38335
rect 20856 38301 20864 38335
rect 22652 38428 22704 38480
rect 26792 38496 26844 38548
rect 21548 38360 21600 38412
rect 20812 38292 20864 38301
rect 21640 38292 21692 38344
rect 21456 38224 21508 38276
rect 22744 38403 22796 38412
rect 22744 38369 22753 38403
rect 22753 38369 22787 38403
rect 22787 38369 22796 38403
rect 22744 38360 22796 38369
rect 24584 38360 24636 38412
rect 28356 38428 28408 38480
rect 28632 38539 28684 38548
rect 28632 38505 28641 38539
rect 28641 38505 28675 38539
rect 28675 38505 28684 38539
rect 28632 38496 28684 38505
rect 29184 38539 29236 38548
rect 29184 38505 29193 38539
rect 29193 38505 29227 38539
rect 29227 38505 29236 38539
rect 29184 38496 29236 38505
rect 29552 38496 29604 38548
rect 29736 38539 29788 38548
rect 29736 38505 29745 38539
rect 29745 38505 29779 38539
rect 29779 38505 29788 38539
rect 29736 38496 29788 38505
rect 30564 38539 30616 38548
rect 30564 38505 30573 38539
rect 30573 38505 30607 38539
rect 30607 38505 30616 38539
rect 30564 38496 30616 38505
rect 31116 38496 31168 38548
rect 32772 38539 32824 38548
rect 32772 38505 32781 38539
rect 32781 38505 32815 38539
rect 32815 38505 32824 38539
rect 32772 38496 32824 38505
rect 35624 38496 35676 38548
rect 36452 38496 36504 38548
rect 39212 38496 39264 38548
rect 41052 38496 41104 38548
rect 29276 38428 29328 38480
rect 33232 38428 33284 38480
rect 34888 38428 34940 38480
rect 40500 38428 40552 38480
rect 21824 38335 21876 38344
rect 21824 38301 21833 38335
rect 21833 38301 21867 38335
rect 21867 38301 21876 38335
rect 21824 38292 21876 38301
rect 22468 38335 22520 38344
rect 22468 38301 22477 38335
rect 22477 38301 22511 38335
rect 22511 38301 22520 38335
rect 22468 38292 22520 38301
rect 22744 38224 22796 38276
rect 22008 38156 22060 38208
rect 23204 38156 23256 38208
rect 24768 38335 24820 38344
rect 24768 38301 24772 38335
rect 24772 38301 24806 38335
rect 24806 38301 24820 38335
rect 24768 38292 24820 38301
rect 23756 38224 23808 38276
rect 23572 38156 23624 38208
rect 25872 38292 25924 38344
rect 26240 38292 26292 38344
rect 29644 38360 29696 38412
rect 26700 38335 26752 38344
rect 26700 38301 26745 38335
rect 26745 38301 26752 38335
rect 26700 38292 26752 38301
rect 26976 38292 27028 38344
rect 27988 38335 28040 38344
rect 27988 38301 27997 38335
rect 27997 38301 28031 38335
rect 28031 38301 28040 38335
rect 27988 38292 28040 38301
rect 28172 38335 28224 38344
rect 28172 38301 28179 38335
rect 28179 38301 28224 38335
rect 28172 38292 28224 38301
rect 28356 38335 28408 38344
rect 28356 38301 28365 38335
rect 28365 38301 28399 38335
rect 28399 38301 28408 38335
rect 28356 38292 28408 38301
rect 28632 38292 28684 38344
rect 30840 38292 30892 38344
rect 25688 38199 25740 38208
rect 25688 38165 25697 38199
rect 25697 38165 25731 38199
rect 25731 38165 25740 38199
rect 25688 38156 25740 38165
rect 26332 38156 26384 38208
rect 26608 38267 26660 38276
rect 26608 38233 26617 38267
rect 26617 38233 26651 38267
rect 26651 38233 26660 38267
rect 26608 38224 26660 38233
rect 26884 38156 26936 38208
rect 27896 38156 27948 38208
rect 28172 38156 28224 38208
rect 29920 38267 29972 38276
rect 29920 38233 29929 38267
rect 29929 38233 29963 38267
rect 29963 38233 29972 38267
rect 29920 38224 29972 38233
rect 30196 38224 30248 38276
rect 30012 38156 30064 38208
rect 32312 38360 32364 38412
rect 32772 38360 32824 38412
rect 31024 38292 31076 38344
rect 31576 38224 31628 38276
rect 33324 38335 33376 38344
rect 33324 38301 33333 38335
rect 33333 38301 33367 38335
rect 33367 38301 33376 38335
rect 33324 38292 33376 38301
rect 33416 38335 33468 38344
rect 33416 38301 33425 38335
rect 33425 38301 33459 38335
rect 33459 38301 33468 38335
rect 33416 38292 33468 38301
rect 34152 38360 34204 38412
rect 32220 38224 32272 38276
rect 33048 38224 33100 38276
rect 33232 38224 33284 38276
rect 34428 38292 34480 38344
rect 34888 38335 34940 38344
rect 34888 38301 34897 38335
rect 34897 38301 34931 38335
rect 34931 38301 34940 38335
rect 34888 38292 34940 38301
rect 34520 38224 34572 38276
rect 36820 38292 36872 38344
rect 39396 38360 39448 38412
rect 41052 38403 41104 38412
rect 41052 38369 41061 38403
rect 41061 38369 41095 38403
rect 41095 38369 41104 38403
rect 41052 38360 41104 38369
rect 37096 38335 37148 38344
rect 37096 38301 37105 38335
rect 37105 38301 37139 38335
rect 37139 38301 37148 38335
rect 37096 38292 37148 38301
rect 37372 38335 37424 38344
rect 37372 38301 37381 38335
rect 37381 38301 37415 38335
rect 37415 38301 37424 38335
rect 37372 38292 37424 38301
rect 37648 38335 37700 38344
rect 37648 38301 37657 38335
rect 37657 38301 37691 38335
rect 37691 38301 37700 38335
rect 37648 38292 37700 38301
rect 37832 38335 37884 38344
rect 37832 38301 37841 38335
rect 37841 38301 37875 38335
rect 37875 38301 37884 38335
rect 37832 38292 37884 38301
rect 40040 38335 40092 38344
rect 40040 38301 40049 38335
rect 40049 38301 40083 38335
rect 40083 38301 40092 38335
rect 40040 38292 40092 38301
rect 40132 38335 40184 38344
rect 40132 38301 40141 38335
rect 40141 38301 40175 38335
rect 40175 38301 40184 38335
rect 40132 38292 40184 38301
rect 41144 38335 41196 38344
rect 41144 38301 41153 38335
rect 41153 38301 41187 38335
rect 41187 38301 41196 38335
rect 41144 38292 41196 38301
rect 41880 38292 41932 38344
rect 35072 38267 35124 38276
rect 35072 38233 35081 38267
rect 35081 38233 35115 38267
rect 35115 38233 35124 38267
rect 35072 38224 35124 38233
rect 35164 38267 35216 38276
rect 35164 38233 35173 38267
rect 35173 38233 35207 38267
rect 35207 38233 35216 38267
rect 35164 38224 35216 38233
rect 35992 38199 36044 38208
rect 35992 38165 36001 38199
rect 36001 38165 36035 38199
rect 36035 38165 36044 38199
rect 35992 38156 36044 38165
rect 36636 38156 36688 38208
rect 37004 38156 37056 38208
rect 37924 38224 37976 38276
rect 40684 38224 40736 38276
rect 38476 38156 38528 38208
rect 39856 38156 39908 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 18236 37995 18288 38004
rect 18236 37961 18245 37995
rect 18245 37961 18279 37995
rect 18279 37961 18288 37995
rect 18236 37952 18288 37961
rect 15200 37927 15252 37936
rect 15200 37893 15209 37927
rect 15209 37893 15243 37927
rect 15243 37893 15252 37927
rect 15200 37884 15252 37893
rect 19248 37995 19300 38004
rect 19248 37961 19257 37995
rect 19257 37961 19291 37995
rect 19291 37961 19300 37995
rect 19248 37952 19300 37961
rect 23940 37952 23992 38004
rect 24676 37952 24728 38004
rect 25136 37952 25188 38004
rect 20168 37884 20220 37936
rect 20812 37884 20864 37936
rect 21088 37884 21140 37936
rect 22284 37927 22336 37936
rect 22284 37893 22293 37927
rect 22293 37893 22327 37927
rect 22327 37893 22336 37927
rect 22284 37884 22336 37893
rect 23112 37884 23164 37936
rect 20904 37859 20956 37868
rect 20904 37825 20913 37859
rect 20913 37825 20947 37859
rect 20947 37825 20956 37859
rect 20904 37816 20956 37825
rect 21272 37859 21324 37868
rect 21272 37825 21281 37859
rect 21281 37825 21315 37859
rect 21315 37825 21324 37859
rect 21272 37816 21324 37825
rect 21456 37859 21508 37868
rect 21456 37825 21465 37859
rect 21465 37825 21499 37859
rect 21499 37825 21508 37859
rect 21456 37816 21508 37825
rect 22100 37816 22152 37868
rect 18512 37748 18564 37800
rect 19248 37748 19300 37800
rect 19432 37791 19484 37800
rect 19432 37757 19441 37791
rect 19441 37757 19475 37791
rect 19475 37757 19484 37791
rect 19432 37748 19484 37757
rect 20996 37791 21048 37800
rect 20996 37757 21005 37791
rect 21005 37757 21039 37791
rect 21039 37757 21048 37791
rect 20996 37748 21048 37757
rect 22652 37859 22704 37868
rect 22652 37825 22661 37859
rect 22661 37825 22695 37859
rect 22695 37825 22704 37859
rect 22652 37816 22704 37825
rect 23296 37884 23348 37936
rect 24216 37859 24268 37868
rect 24216 37825 24225 37859
rect 24225 37825 24259 37859
rect 24259 37825 24268 37859
rect 24216 37816 24268 37825
rect 24676 37816 24728 37868
rect 24768 37859 24820 37868
rect 24768 37825 24777 37859
rect 24777 37825 24811 37859
rect 24811 37825 24820 37859
rect 24768 37816 24820 37825
rect 23296 37748 23348 37800
rect 23572 37748 23624 37800
rect 24032 37791 24084 37800
rect 24032 37757 24041 37791
rect 24041 37757 24075 37791
rect 24075 37757 24084 37791
rect 24032 37748 24084 37757
rect 17224 37680 17276 37732
rect 21364 37680 21416 37732
rect 26608 37952 26660 38004
rect 26332 37927 26384 37936
rect 26332 37893 26341 37927
rect 26341 37893 26375 37927
rect 26375 37893 26384 37927
rect 26332 37884 26384 37893
rect 25228 37816 25280 37868
rect 25688 37859 25740 37868
rect 25688 37825 25733 37859
rect 25733 37825 25740 37859
rect 25688 37816 25740 37825
rect 25872 37859 25924 37868
rect 25872 37825 25881 37859
rect 25881 37825 25915 37859
rect 25915 37825 25924 37859
rect 25872 37816 25924 37825
rect 26148 37816 26200 37868
rect 26240 37748 26292 37800
rect 26792 37816 26844 37868
rect 27896 37884 27948 37936
rect 27436 37859 27488 37868
rect 27436 37825 27443 37859
rect 27443 37825 27488 37859
rect 27436 37816 27488 37825
rect 27528 37859 27580 37868
rect 27528 37825 27537 37859
rect 27537 37825 27571 37859
rect 27571 37825 27580 37859
rect 27528 37816 27580 37825
rect 28632 37927 28684 37936
rect 28632 37893 28641 37927
rect 28641 37893 28675 37927
rect 28675 37893 28684 37927
rect 28632 37884 28684 37893
rect 30380 37884 30432 37936
rect 30564 37952 30616 38004
rect 30748 37952 30800 38004
rect 31760 37995 31812 38004
rect 31760 37961 31769 37995
rect 31769 37961 31803 37995
rect 31803 37961 31812 37995
rect 31760 37952 31812 37961
rect 32312 37995 32364 38004
rect 32312 37961 32321 37995
rect 32321 37961 32355 37995
rect 32355 37961 32364 37995
rect 32312 37952 32364 37961
rect 26516 37680 26568 37732
rect 27252 37680 27304 37732
rect 27344 37680 27396 37732
rect 28448 37859 28500 37868
rect 28448 37825 28485 37859
rect 28485 37825 28500 37859
rect 28448 37816 28500 37825
rect 28816 37859 28868 37868
rect 28816 37825 28830 37859
rect 28830 37825 28864 37859
rect 28864 37825 28868 37859
rect 28816 37816 28868 37825
rect 27988 37748 28040 37800
rect 29184 37748 29236 37800
rect 16212 37655 16264 37664
rect 16212 37621 16221 37655
rect 16221 37621 16255 37655
rect 16255 37621 16264 37655
rect 16212 37612 16264 37621
rect 17132 37655 17184 37664
rect 17132 37621 17141 37655
rect 17141 37621 17175 37655
rect 17175 37621 17184 37655
rect 17132 37612 17184 37621
rect 21916 37612 21968 37664
rect 22560 37612 22612 37664
rect 26884 37612 26936 37664
rect 27712 37612 27764 37664
rect 27896 37655 27948 37664
rect 27896 37621 27905 37655
rect 27905 37621 27939 37655
rect 27939 37621 27948 37655
rect 27896 37612 27948 37621
rect 28172 37680 28224 37732
rect 30472 37859 30524 37868
rect 30472 37825 30481 37859
rect 30481 37825 30515 37859
rect 30515 37825 30524 37859
rect 30472 37816 30524 37825
rect 30656 37816 30708 37868
rect 29736 37791 29788 37800
rect 29736 37757 29745 37791
rect 29745 37757 29779 37791
rect 29779 37757 29788 37791
rect 29736 37748 29788 37757
rect 30196 37748 30248 37800
rect 28816 37612 28868 37664
rect 29000 37655 29052 37664
rect 29000 37621 29009 37655
rect 29009 37621 29043 37655
rect 29043 37621 29052 37655
rect 29000 37612 29052 37621
rect 29920 37680 29972 37732
rect 31484 37859 31536 37868
rect 31484 37825 31493 37859
rect 31493 37825 31527 37859
rect 31527 37825 31536 37859
rect 31484 37816 31536 37825
rect 32404 37884 32456 37936
rect 34704 37884 34756 37936
rect 32588 37859 32640 37868
rect 32588 37825 32597 37859
rect 32597 37825 32631 37859
rect 32631 37825 32640 37859
rect 32588 37816 32640 37825
rect 32772 37859 32824 37868
rect 32772 37825 32781 37859
rect 32781 37825 32815 37859
rect 32815 37825 32824 37859
rect 32772 37816 32824 37825
rect 32864 37859 32916 37868
rect 32864 37825 32873 37859
rect 32873 37825 32907 37859
rect 32907 37825 32916 37859
rect 32864 37816 32916 37825
rect 33600 37816 33652 37868
rect 33968 37859 34020 37868
rect 33968 37825 33978 37859
rect 33978 37825 34012 37859
rect 34012 37825 34020 37859
rect 33968 37816 34020 37825
rect 34152 37859 34204 37868
rect 34152 37825 34161 37859
rect 34161 37825 34195 37859
rect 34195 37825 34204 37859
rect 34152 37816 34204 37825
rect 34428 37816 34480 37868
rect 35256 37952 35308 38004
rect 36084 37952 36136 38004
rect 37372 37952 37424 38004
rect 35532 37859 35584 37868
rect 35532 37825 35541 37859
rect 35541 37825 35575 37859
rect 35575 37825 35584 37859
rect 35532 37816 35584 37825
rect 35900 37816 35952 37868
rect 35808 37748 35860 37800
rect 36452 37859 36504 37868
rect 36452 37825 36461 37859
rect 36461 37825 36495 37859
rect 36495 37825 36504 37859
rect 36452 37816 36504 37825
rect 36544 37859 36596 37868
rect 36544 37825 36553 37859
rect 36553 37825 36587 37859
rect 36587 37825 36596 37859
rect 36544 37816 36596 37825
rect 36820 37816 36872 37868
rect 37004 37816 37056 37868
rect 39028 37952 39080 38004
rect 39488 37995 39540 38004
rect 39488 37961 39497 37995
rect 39497 37961 39531 37995
rect 39531 37961 39540 37995
rect 39488 37952 39540 37961
rect 40040 37952 40092 38004
rect 40960 37884 41012 37936
rect 41144 37927 41196 37936
rect 41144 37893 41153 37927
rect 41153 37893 41187 37927
rect 41187 37893 41196 37927
rect 41144 37884 41196 37893
rect 41328 37927 41380 37936
rect 41328 37893 41353 37927
rect 41353 37893 41380 37927
rect 41328 37884 41380 37893
rect 38476 37859 38528 37868
rect 38476 37825 38485 37859
rect 38485 37825 38519 37859
rect 38519 37825 38528 37859
rect 38476 37816 38528 37825
rect 36728 37748 36780 37800
rect 36912 37748 36964 37800
rect 39028 37859 39080 37868
rect 39028 37825 39037 37859
rect 39037 37825 39071 37859
rect 39071 37825 39080 37859
rect 39028 37816 39080 37825
rect 39396 37816 39448 37868
rect 40040 37859 40092 37868
rect 40040 37825 40049 37859
rect 40049 37825 40083 37859
rect 40083 37825 40092 37859
rect 40040 37816 40092 37825
rect 40316 37859 40368 37868
rect 40316 37825 40325 37859
rect 40325 37825 40359 37859
rect 40359 37825 40368 37859
rect 40316 37816 40368 37825
rect 40592 37816 40644 37868
rect 40408 37748 40460 37800
rect 40776 37748 40828 37800
rect 32220 37680 32272 37732
rect 29828 37612 29880 37664
rect 30012 37655 30064 37664
rect 30012 37621 30021 37655
rect 30021 37621 30055 37655
rect 30055 37621 30064 37655
rect 30012 37612 30064 37621
rect 31208 37612 31260 37664
rect 34796 37680 34848 37732
rect 35072 37680 35124 37732
rect 36452 37680 36504 37732
rect 33508 37612 33560 37664
rect 34520 37612 34572 37664
rect 34704 37612 34756 37664
rect 38200 37680 38252 37732
rect 36636 37612 36688 37664
rect 39212 37612 39264 37664
rect 41144 37612 41196 37664
rect 41512 37655 41564 37664
rect 41512 37621 41521 37655
rect 41521 37621 41555 37655
rect 41555 37621 41564 37655
rect 41512 37612 41564 37621
rect 42064 37612 42116 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 14464 37451 14516 37460
rect 14464 37417 14473 37451
rect 14473 37417 14507 37451
rect 14507 37417 14516 37451
rect 14464 37408 14516 37417
rect 15568 37451 15620 37460
rect 15568 37417 15577 37451
rect 15577 37417 15611 37451
rect 15611 37417 15620 37451
rect 15568 37408 15620 37417
rect 16120 37451 16172 37460
rect 16120 37417 16129 37451
rect 16129 37417 16163 37451
rect 16163 37417 16172 37451
rect 16120 37408 16172 37417
rect 16672 37451 16724 37460
rect 16672 37417 16681 37451
rect 16681 37417 16715 37451
rect 16715 37417 16724 37451
rect 16672 37408 16724 37417
rect 17224 37451 17276 37460
rect 17224 37417 17233 37451
rect 17233 37417 17267 37451
rect 17267 37417 17276 37451
rect 17224 37408 17276 37417
rect 17776 37451 17828 37460
rect 17776 37417 17785 37451
rect 17785 37417 17819 37451
rect 17819 37417 17828 37451
rect 17776 37408 17828 37417
rect 23940 37408 23992 37460
rect 16580 37340 16632 37392
rect 19432 37340 19484 37392
rect 20076 37340 20128 37392
rect 21272 37340 21324 37392
rect 16212 37272 16264 37324
rect 19340 37204 19392 37256
rect 21916 37315 21968 37324
rect 21916 37281 21925 37315
rect 21925 37281 21959 37315
rect 21959 37281 21968 37315
rect 21916 37272 21968 37281
rect 19248 37136 19300 37188
rect 22192 37204 22244 37256
rect 22652 37340 22704 37392
rect 24124 37408 24176 37460
rect 25688 37408 25740 37460
rect 25872 37408 25924 37460
rect 27528 37408 27580 37460
rect 28632 37408 28684 37460
rect 24032 37272 24084 37324
rect 24308 37272 24360 37324
rect 24584 37315 24636 37324
rect 24584 37281 24593 37315
rect 24593 37281 24627 37315
rect 24627 37281 24636 37315
rect 24584 37272 24636 37281
rect 19432 37111 19484 37120
rect 19432 37077 19441 37111
rect 19441 37077 19475 37111
rect 19475 37077 19484 37111
rect 19432 37068 19484 37077
rect 20260 37111 20312 37120
rect 20260 37077 20269 37111
rect 20269 37077 20303 37111
rect 20303 37077 20312 37111
rect 20260 37068 20312 37077
rect 22376 37068 22428 37120
rect 23112 37204 23164 37256
rect 23204 37204 23256 37256
rect 23480 37247 23532 37256
rect 23480 37213 23490 37247
rect 23490 37213 23524 37247
rect 23524 37213 23532 37247
rect 23480 37204 23532 37213
rect 23848 37247 23900 37256
rect 23848 37213 23862 37247
rect 23862 37213 23896 37247
rect 23896 37213 23900 37247
rect 26332 37340 26384 37392
rect 27252 37340 27304 37392
rect 28172 37340 28224 37392
rect 25228 37315 25280 37324
rect 25228 37281 25237 37315
rect 25237 37281 25271 37315
rect 25271 37281 25280 37315
rect 25228 37272 25280 37281
rect 27896 37272 27948 37324
rect 28448 37272 28500 37324
rect 29092 37272 29144 37324
rect 23848 37204 23900 37213
rect 24860 37247 24912 37256
rect 24860 37213 24869 37247
rect 24869 37213 24903 37247
rect 24903 37213 24912 37247
rect 24860 37204 24912 37213
rect 26056 37204 26108 37256
rect 26424 37247 26476 37256
rect 26424 37213 26433 37247
rect 26433 37213 26467 37247
rect 26467 37213 26476 37247
rect 26424 37204 26476 37213
rect 26792 37204 26844 37256
rect 23572 37136 23624 37188
rect 24124 37136 24176 37188
rect 24952 37136 25004 37188
rect 25780 37136 25832 37188
rect 27252 37204 27304 37256
rect 27620 37247 27672 37256
rect 27620 37213 27629 37247
rect 27629 37213 27663 37247
rect 27663 37213 27672 37247
rect 27620 37204 27672 37213
rect 28264 37247 28316 37256
rect 28264 37213 28273 37247
rect 28273 37213 28307 37247
rect 28307 37213 28316 37247
rect 28264 37204 28316 37213
rect 31024 37408 31076 37460
rect 31484 37408 31536 37460
rect 32220 37408 32272 37460
rect 31760 37340 31812 37392
rect 32588 37340 32640 37392
rect 31024 37272 31076 37324
rect 36360 37408 36412 37460
rect 36912 37451 36964 37460
rect 36912 37417 36921 37451
rect 36921 37417 36955 37451
rect 36955 37417 36964 37451
rect 36912 37408 36964 37417
rect 37464 37451 37516 37460
rect 37464 37417 37473 37451
rect 37473 37417 37507 37451
rect 37507 37417 37516 37451
rect 37464 37408 37516 37417
rect 34152 37340 34204 37392
rect 34796 37340 34848 37392
rect 33048 37272 33100 37324
rect 29276 37204 29328 37256
rect 29920 37247 29972 37256
rect 29920 37213 29929 37247
rect 29929 37213 29963 37247
rect 29963 37213 29972 37247
rect 29920 37204 29972 37213
rect 30012 37204 30064 37256
rect 30932 37204 30984 37256
rect 32036 37247 32088 37256
rect 32036 37213 32045 37247
rect 32045 37213 32079 37247
rect 32079 37213 32088 37247
rect 32036 37204 32088 37213
rect 22652 37068 22704 37120
rect 24676 37068 24728 37120
rect 29368 37136 29420 37188
rect 30288 37136 30340 37188
rect 30380 37136 30432 37188
rect 27712 37068 27764 37120
rect 30564 37068 30616 37120
rect 31852 37068 31904 37120
rect 32128 37179 32180 37188
rect 32128 37145 32137 37179
rect 32137 37145 32171 37179
rect 32171 37145 32180 37179
rect 32128 37136 32180 37145
rect 32588 37204 32640 37256
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 33232 37136 33284 37188
rect 33968 37272 34020 37324
rect 34152 37204 34204 37256
rect 34520 37204 34572 37256
rect 34796 37204 34848 37256
rect 35072 37247 35124 37256
rect 35072 37213 35079 37247
rect 35079 37213 35124 37247
rect 32404 37068 32456 37120
rect 33508 37068 33560 37120
rect 33600 37068 33652 37120
rect 34428 37136 34480 37188
rect 35072 37204 35124 37213
rect 35164 37247 35216 37256
rect 35164 37213 35173 37247
rect 35173 37213 35207 37247
rect 35207 37213 35216 37247
rect 35164 37204 35216 37213
rect 37096 37340 37148 37392
rect 39856 37408 39908 37460
rect 40684 37451 40736 37460
rect 40684 37417 40693 37451
rect 40693 37417 40727 37451
rect 40727 37417 40736 37451
rect 40684 37408 40736 37417
rect 35624 37204 35676 37256
rect 36636 37272 36688 37324
rect 36452 37204 36504 37256
rect 36820 37204 36872 37256
rect 39396 37340 39448 37392
rect 39580 37340 39632 37392
rect 40776 37340 40828 37392
rect 41420 37383 41472 37392
rect 41420 37349 41429 37383
rect 41429 37349 41463 37383
rect 41463 37349 41472 37383
rect 41420 37340 41472 37349
rect 39304 37315 39356 37324
rect 39304 37281 39313 37315
rect 39313 37281 39347 37315
rect 39347 37281 39356 37315
rect 39304 37272 39356 37281
rect 38108 37247 38160 37256
rect 38108 37213 38117 37247
rect 38117 37213 38151 37247
rect 38151 37213 38160 37247
rect 38108 37204 38160 37213
rect 38200 37247 38252 37256
rect 38200 37213 38209 37247
rect 38209 37213 38243 37247
rect 38243 37213 38252 37247
rect 38200 37204 38252 37213
rect 38292 37204 38344 37256
rect 38476 37247 38528 37256
rect 38476 37213 38485 37247
rect 38485 37213 38519 37247
rect 38519 37213 38528 37247
rect 38476 37204 38528 37213
rect 38660 37247 38712 37256
rect 38660 37213 38669 37247
rect 38669 37213 38703 37247
rect 38703 37213 38712 37247
rect 38660 37204 38712 37213
rect 34244 37111 34296 37120
rect 34244 37077 34253 37111
rect 34253 37077 34287 37111
rect 34287 37077 34296 37111
rect 34244 37068 34296 37077
rect 34612 37068 34664 37120
rect 36176 37136 36228 37188
rect 36544 37179 36596 37188
rect 36544 37145 36553 37179
rect 36553 37145 36587 37179
rect 36587 37145 36596 37179
rect 36544 37136 36596 37145
rect 37188 37136 37240 37188
rect 35072 37068 35124 37120
rect 35440 37068 35492 37120
rect 40224 37247 40276 37256
rect 40224 37213 40231 37247
rect 40231 37213 40276 37247
rect 40224 37204 40276 37213
rect 40592 37204 40644 37256
rect 41144 37247 41196 37256
rect 41144 37213 41153 37247
rect 41153 37213 41187 37247
rect 41187 37213 41196 37247
rect 41144 37204 41196 37213
rect 41236 37247 41288 37256
rect 41236 37213 41245 37247
rect 41245 37213 41279 37247
rect 41279 37213 41288 37247
rect 41236 37204 41288 37213
rect 41880 37247 41932 37256
rect 41880 37213 41889 37247
rect 41889 37213 41923 37247
rect 41923 37213 41932 37247
rect 41880 37204 41932 37213
rect 40316 37179 40368 37188
rect 40316 37145 40325 37179
rect 40325 37145 40359 37179
rect 40359 37145 40368 37179
rect 40316 37136 40368 37145
rect 40776 37136 40828 37188
rect 41328 37136 41380 37188
rect 41972 37136 42024 37188
rect 40224 37068 40276 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 16212 36864 16264 36916
rect 22376 36864 22428 36916
rect 22468 36864 22520 36916
rect 23664 36864 23716 36916
rect 25872 36864 25924 36916
rect 16120 36796 16172 36848
rect 17500 36796 17552 36848
rect 16856 36771 16908 36780
rect 16856 36737 16865 36771
rect 16865 36737 16899 36771
rect 16899 36737 16908 36771
rect 16856 36728 16908 36737
rect 20720 36796 20772 36848
rect 23112 36796 23164 36848
rect 24400 36796 24452 36848
rect 16212 36660 16264 36712
rect 19432 36728 19484 36780
rect 20260 36728 20312 36780
rect 22652 36728 22704 36780
rect 24124 36771 24176 36780
rect 24124 36737 24128 36771
rect 24128 36737 24162 36771
rect 24162 36737 24176 36771
rect 24124 36728 24176 36737
rect 24308 36771 24360 36780
rect 24308 36737 24317 36771
rect 24317 36737 24351 36771
rect 24351 36737 24360 36771
rect 24308 36728 24360 36737
rect 24768 36796 24820 36848
rect 26424 36907 26476 36916
rect 26424 36873 26433 36907
rect 26433 36873 26467 36907
rect 26467 36873 26476 36907
rect 26424 36864 26476 36873
rect 27344 36864 27396 36916
rect 28540 36907 28592 36916
rect 28540 36873 28549 36907
rect 28549 36873 28583 36907
rect 28583 36873 28592 36907
rect 28540 36864 28592 36873
rect 30472 36907 30524 36916
rect 30472 36873 30481 36907
rect 30481 36873 30515 36907
rect 30515 36873 30524 36907
rect 30472 36864 30524 36873
rect 30564 36864 30616 36916
rect 32128 36864 32180 36916
rect 32864 36864 32916 36916
rect 33232 36864 33284 36916
rect 33784 36864 33836 36916
rect 26700 36796 26752 36848
rect 24676 36728 24728 36780
rect 25044 36771 25096 36780
rect 25044 36737 25053 36771
rect 25053 36737 25087 36771
rect 25087 36737 25096 36771
rect 25044 36728 25096 36737
rect 25412 36728 25464 36780
rect 25780 36771 25832 36780
rect 25780 36737 25789 36771
rect 25789 36737 25823 36771
rect 25823 36737 25832 36771
rect 25780 36728 25832 36737
rect 25872 36771 25924 36780
rect 25872 36737 25882 36771
rect 25882 36737 25916 36771
rect 25916 36737 25924 36771
rect 25872 36728 25924 36737
rect 26332 36728 26384 36780
rect 35348 36864 35400 36916
rect 38200 36864 38252 36916
rect 39120 36864 39172 36916
rect 33968 36839 34020 36848
rect 33968 36805 33977 36839
rect 33977 36805 34011 36839
rect 34011 36805 34020 36839
rect 33968 36796 34020 36805
rect 34336 36796 34388 36848
rect 14096 36635 14148 36644
rect 14096 36601 14105 36635
rect 14105 36601 14139 36635
rect 14139 36601 14148 36635
rect 14096 36592 14148 36601
rect 19984 36524 20036 36576
rect 20168 36567 20220 36576
rect 20168 36533 20177 36567
rect 20177 36533 20211 36567
rect 20211 36533 20220 36567
rect 20168 36524 20220 36533
rect 21548 36592 21600 36644
rect 22284 36660 22336 36712
rect 22560 36703 22612 36712
rect 22560 36669 22569 36703
rect 22569 36669 22603 36703
rect 22603 36669 22612 36703
rect 22560 36660 22612 36669
rect 23388 36660 23440 36712
rect 26148 36660 26200 36712
rect 26516 36660 26568 36712
rect 27068 36660 27120 36712
rect 27528 36771 27580 36780
rect 27528 36737 27537 36771
rect 27537 36737 27571 36771
rect 27571 36737 27580 36771
rect 27528 36728 27580 36737
rect 28080 36728 28132 36780
rect 29092 36728 29144 36780
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 29460 36771 29512 36780
rect 29460 36737 29469 36771
rect 29469 36737 29503 36771
rect 29503 36737 29512 36771
rect 29460 36728 29512 36737
rect 27436 36660 27488 36712
rect 29000 36660 29052 36712
rect 30104 36771 30156 36780
rect 30104 36737 30113 36771
rect 30113 36737 30147 36771
rect 30147 36737 30156 36771
rect 30104 36728 30156 36737
rect 30196 36771 30248 36780
rect 30196 36737 30205 36771
rect 30205 36737 30239 36771
rect 30239 36737 30248 36771
rect 30196 36728 30248 36737
rect 30288 36771 30340 36780
rect 30288 36737 30297 36771
rect 30297 36737 30331 36771
rect 30331 36737 30340 36771
rect 30288 36728 30340 36737
rect 30932 36728 30984 36780
rect 31208 36728 31260 36780
rect 31576 36728 31628 36780
rect 32496 36771 32548 36780
rect 32496 36737 32505 36771
rect 32505 36737 32539 36771
rect 32539 36737 32548 36771
rect 32496 36728 32548 36737
rect 32680 36771 32732 36780
rect 32680 36737 32689 36771
rect 32689 36737 32723 36771
rect 32723 36737 32732 36771
rect 32680 36728 32732 36737
rect 32772 36771 32824 36780
rect 32772 36737 32781 36771
rect 32781 36737 32815 36771
rect 32815 36737 32824 36771
rect 32772 36728 32824 36737
rect 33508 36728 33560 36780
rect 33600 36728 33652 36780
rect 22836 36592 22888 36644
rect 30564 36660 30616 36712
rect 32312 36660 32364 36712
rect 33140 36660 33192 36712
rect 33876 36728 33928 36780
rect 34152 36771 34204 36780
rect 35808 36796 35860 36848
rect 36176 36796 36228 36848
rect 38292 36796 38344 36848
rect 34152 36737 34166 36771
rect 34166 36737 34200 36771
rect 34200 36737 34204 36771
rect 34152 36728 34204 36737
rect 33600 36592 33652 36644
rect 34152 36592 34204 36644
rect 35164 36728 35216 36780
rect 35900 36728 35952 36780
rect 36360 36771 36412 36780
rect 36360 36737 36369 36771
rect 36369 36737 36403 36771
rect 36403 36737 36412 36771
rect 36360 36728 36412 36737
rect 36636 36771 36688 36780
rect 36636 36737 36645 36771
rect 36645 36737 36679 36771
rect 36679 36737 36688 36771
rect 36636 36728 36688 36737
rect 36820 36728 36872 36780
rect 37648 36728 37700 36780
rect 38384 36771 38436 36780
rect 38384 36737 38393 36771
rect 38393 36737 38427 36771
rect 38427 36737 38436 36771
rect 38384 36728 38436 36737
rect 39672 36839 39724 36848
rect 39672 36805 39681 36839
rect 39681 36805 39715 36839
rect 39715 36805 39724 36839
rect 39672 36796 39724 36805
rect 39948 36796 40000 36848
rect 40776 36907 40828 36916
rect 40776 36873 40785 36907
rect 40785 36873 40819 36907
rect 40819 36873 40828 36907
rect 40776 36864 40828 36873
rect 41420 36864 41472 36916
rect 41972 36907 42024 36916
rect 41972 36873 41981 36907
rect 41981 36873 42015 36907
rect 42015 36873 42024 36907
rect 41972 36864 42024 36873
rect 35900 36592 35952 36644
rect 37004 36592 37056 36644
rect 37924 36592 37976 36644
rect 38016 36592 38068 36644
rect 38660 36592 38712 36644
rect 39396 36728 39448 36780
rect 40132 36771 40184 36780
rect 40132 36737 40141 36771
rect 40141 36737 40175 36771
rect 40175 36737 40184 36771
rect 40132 36728 40184 36737
rect 40224 36771 40276 36780
rect 40224 36737 40234 36771
rect 40234 36737 40268 36771
rect 40268 36737 40276 36771
rect 40224 36728 40276 36737
rect 40316 36728 40368 36780
rect 40592 36771 40644 36780
rect 40592 36737 40606 36771
rect 40606 36737 40640 36771
rect 40640 36737 40644 36771
rect 40592 36728 40644 36737
rect 39488 36660 39540 36712
rect 38936 36592 38988 36644
rect 22376 36524 22428 36576
rect 23204 36524 23256 36576
rect 23388 36524 23440 36576
rect 23664 36524 23716 36576
rect 25136 36567 25188 36576
rect 25136 36533 25145 36567
rect 25145 36533 25179 36567
rect 25179 36533 25188 36567
rect 25136 36524 25188 36533
rect 26332 36524 26384 36576
rect 27620 36524 27672 36576
rect 30380 36524 30432 36576
rect 31208 36524 31260 36576
rect 33692 36524 33744 36576
rect 33876 36524 33928 36576
rect 36360 36524 36412 36576
rect 37740 36524 37792 36576
rect 38108 36524 38160 36576
rect 41236 36771 41288 36780
rect 41236 36737 41245 36771
rect 41245 36737 41279 36771
rect 41279 36737 41288 36771
rect 41236 36728 41288 36737
rect 41512 36728 41564 36780
rect 43352 36771 43404 36780
rect 43352 36737 43361 36771
rect 43361 36737 43395 36771
rect 43395 36737 43404 36771
rect 43352 36728 43404 36737
rect 43996 36728 44048 36780
rect 41052 36660 41104 36712
rect 42524 36660 42576 36712
rect 41788 36592 41840 36644
rect 41328 36567 41380 36576
rect 41328 36533 41337 36567
rect 41337 36533 41371 36567
rect 41371 36533 41380 36567
rect 41328 36524 41380 36533
rect 42248 36524 42300 36576
rect 42984 36524 43036 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 9680 36363 9732 36372
rect 9680 36329 9689 36363
rect 9689 36329 9723 36363
rect 9723 36329 9732 36363
rect 9680 36320 9732 36329
rect 17776 36363 17828 36372
rect 17776 36329 17785 36363
rect 17785 36329 17819 36363
rect 17819 36329 17828 36363
rect 17776 36320 17828 36329
rect 19340 36320 19392 36372
rect 21548 36320 21600 36372
rect 22928 36320 22980 36372
rect 24952 36320 25004 36372
rect 26608 36320 26660 36372
rect 26792 36320 26844 36372
rect 28908 36320 28960 36372
rect 30472 36320 30524 36372
rect 30840 36320 30892 36372
rect 31392 36320 31444 36372
rect 32680 36363 32732 36372
rect 32680 36329 32689 36363
rect 32689 36329 32723 36363
rect 32723 36329 32732 36363
rect 32680 36320 32732 36329
rect 33692 36363 33744 36372
rect 33692 36329 33701 36363
rect 33701 36329 33735 36363
rect 33735 36329 33744 36363
rect 33692 36320 33744 36329
rect 16856 36184 16908 36236
rect 19156 36184 19208 36236
rect 20076 36227 20128 36236
rect 20076 36193 20085 36227
rect 20085 36193 20119 36227
rect 20119 36193 20128 36227
rect 20076 36184 20128 36193
rect 23572 36252 23624 36304
rect 16488 36159 16540 36168
rect 16488 36125 16497 36159
rect 16497 36125 16531 36159
rect 16531 36125 16540 36159
rect 16488 36116 16540 36125
rect 20168 36116 20220 36168
rect 12624 36048 12676 36100
rect 10416 36023 10468 36032
rect 10416 35989 10425 36023
rect 10425 35989 10459 36023
rect 10459 35989 10468 36023
rect 10416 35980 10468 35989
rect 17132 35980 17184 36032
rect 20076 36048 20128 36100
rect 22468 36159 22520 36168
rect 22468 36125 22477 36159
rect 22477 36125 22511 36159
rect 22511 36125 22520 36159
rect 22468 36116 22520 36125
rect 22836 36159 22888 36168
rect 22836 36125 22845 36159
rect 22845 36125 22879 36159
rect 22879 36125 22888 36159
rect 22836 36116 22888 36125
rect 22928 36116 22980 36168
rect 23848 36184 23900 36236
rect 23664 36159 23716 36168
rect 23664 36125 23673 36159
rect 23673 36125 23707 36159
rect 23707 36125 23716 36159
rect 23664 36116 23716 36125
rect 18788 36023 18840 36032
rect 18788 35989 18797 36023
rect 18797 35989 18831 36023
rect 18831 35989 18840 36023
rect 18788 35980 18840 35989
rect 24032 36252 24084 36304
rect 24492 36252 24544 36304
rect 26056 36295 26108 36304
rect 26056 36261 26065 36295
rect 26065 36261 26099 36295
rect 26099 36261 26108 36295
rect 26056 36252 26108 36261
rect 29276 36252 29328 36304
rect 24584 36116 24636 36168
rect 23940 35980 23992 36032
rect 24768 35980 24820 36032
rect 25504 36116 25556 36168
rect 26240 36159 26292 36168
rect 26240 36125 26249 36159
rect 26249 36125 26283 36159
rect 26283 36125 26292 36159
rect 26240 36116 26292 36125
rect 26424 36159 26476 36168
rect 26424 36125 26433 36159
rect 26433 36125 26467 36159
rect 26467 36125 26476 36159
rect 26424 36116 26476 36125
rect 26608 36159 26660 36168
rect 26608 36125 26617 36159
rect 26617 36125 26651 36159
rect 26651 36125 26660 36159
rect 26608 36116 26660 36125
rect 26700 36116 26752 36168
rect 27068 36116 27120 36168
rect 25320 36091 25372 36100
rect 25320 36057 25329 36091
rect 25329 36057 25363 36091
rect 25363 36057 25372 36091
rect 25320 36048 25372 36057
rect 26056 36048 26108 36100
rect 26516 36048 26568 36100
rect 27804 36116 27856 36168
rect 29184 36116 29236 36168
rect 26148 35980 26200 36032
rect 27344 36091 27396 36100
rect 27344 36057 27353 36091
rect 27353 36057 27387 36091
rect 27387 36057 27396 36091
rect 27344 36048 27396 36057
rect 27528 36048 27580 36100
rect 28172 36091 28224 36100
rect 28172 36057 28181 36091
rect 28181 36057 28215 36091
rect 28215 36057 28224 36091
rect 28172 36048 28224 36057
rect 28816 36048 28868 36100
rect 33600 36184 33652 36236
rect 33876 36320 33928 36372
rect 34428 36320 34480 36372
rect 36728 36320 36780 36372
rect 36820 36320 36872 36372
rect 38752 36320 38804 36372
rect 38936 36363 38988 36372
rect 38936 36329 38945 36363
rect 38945 36329 38979 36363
rect 38979 36329 38988 36363
rect 38936 36320 38988 36329
rect 41144 36320 41196 36372
rect 34888 36252 34940 36304
rect 35624 36252 35676 36304
rect 37280 36252 37332 36304
rect 35348 36184 35400 36236
rect 36268 36184 36320 36236
rect 37740 36252 37792 36304
rect 38200 36252 38252 36304
rect 40132 36252 40184 36304
rect 42340 36320 42392 36372
rect 42616 36320 42668 36372
rect 30472 36159 30524 36168
rect 30472 36125 30481 36159
rect 30481 36125 30515 36159
rect 30515 36125 30524 36159
rect 30472 36116 30524 36125
rect 31484 36116 31536 36168
rect 30656 36091 30708 36100
rect 26700 35980 26752 36032
rect 29644 35980 29696 36032
rect 30656 36057 30665 36091
rect 30665 36057 30699 36091
rect 30699 36057 30708 36091
rect 30656 36048 30708 36057
rect 30840 36048 30892 36100
rect 34244 36116 34296 36168
rect 35900 36159 35952 36168
rect 35900 36125 35909 36159
rect 35909 36125 35943 36159
rect 35943 36125 35952 36159
rect 35900 36116 35952 36125
rect 36728 36159 36780 36168
rect 36728 36125 36737 36159
rect 36737 36125 36771 36159
rect 36771 36125 36780 36159
rect 36728 36116 36780 36125
rect 36820 36159 36872 36168
rect 36820 36125 36830 36159
rect 36830 36125 36864 36159
rect 36864 36125 36872 36159
rect 36820 36116 36872 36125
rect 37280 36116 37332 36168
rect 30288 35980 30340 36032
rect 30380 35980 30432 36032
rect 31116 35980 31168 36032
rect 34980 36048 35032 36100
rect 35164 36048 35216 36100
rect 36084 36048 36136 36100
rect 37740 36116 37792 36168
rect 38016 36159 38068 36168
rect 38016 36125 38023 36159
rect 38023 36125 38068 36159
rect 38016 36116 38068 36125
rect 38200 36159 38252 36168
rect 38200 36125 38209 36159
rect 38209 36125 38243 36159
rect 38243 36125 38252 36159
rect 38200 36116 38252 36125
rect 38292 36159 38344 36168
rect 38292 36125 38306 36159
rect 38306 36125 38340 36159
rect 38340 36125 38344 36159
rect 38292 36116 38344 36125
rect 38752 36116 38804 36168
rect 39396 36116 39448 36168
rect 35256 35980 35308 36032
rect 35532 35980 35584 36032
rect 39212 36091 39264 36100
rect 39212 36057 39221 36091
rect 39221 36057 39255 36091
rect 39255 36057 39264 36091
rect 39212 36048 39264 36057
rect 39304 36091 39356 36100
rect 39304 36057 39313 36091
rect 39313 36057 39347 36091
rect 39347 36057 39356 36091
rect 39304 36048 39356 36057
rect 37464 35980 37516 36032
rect 38476 35980 38528 36032
rect 39856 36048 39908 36100
rect 40224 36116 40276 36168
rect 41696 36184 41748 36236
rect 40500 36159 40552 36168
rect 40500 36125 40514 36159
rect 40514 36125 40548 36159
rect 40548 36125 40552 36159
rect 40500 36116 40552 36125
rect 41236 36116 41288 36168
rect 41420 36116 41472 36168
rect 41512 36116 41564 36168
rect 41880 36116 41932 36168
rect 40316 36091 40368 36100
rect 40316 36057 40325 36091
rect 40325 36057 40359 36091
rect 40359 36057 40368 36091
rect 40316 36048 40368 36057
rect 42616 36048 42668 36100
rect 41052 35980 41104 36032
rect 41788 35980 41840 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1308 35776 1360 35828
rect 15568 35776 15620 35828
rect 16120 35819 16172 35828
rect 16120 35785 16129 35819
rect 16129 35785 16163 35819
rect 16163 35785 16172 35819
rect 16120 35776 16172 35785
rect 16488 35776 16540 35828
rect 14004 35640 14056 35692
rect 15476 35640 15528 35692
rect 17960 35708 18012 35760
rect 17132 35683 17184 35692
rect 17132 35649 17141 35683
rect 17141 35649 17175 35683
rect 17175 35649 17184 35683
rect 17132 35640 17184 35649
rect 16672 35572 16724 35624
rect 16212 35504 16264 35556
rect 18420 35615 18472 35624
rect 18420 35581 18429 35615
rect 18429 35581 18463 35615
rect 18463 35581 18472 35615
rect 18420 35572 18472 35581
rect 16948 35436 17000 35488
rect 17224 35436 17276 35488
rect 18788 35436 18840 35488
rect 19984 35819 20036 35828
rect 19984 35785 19993 35819
rect 19993 35785 20027 35819
rect 20027 35785 20036 35819
rect 19984 35776 20036 35785
rect 21548 35776 21600 35828
rect 22468 35776 22520 35828
rect 22008 35751 22060 35760
rect 22008 35717 22017 35751
rect 22017 35717 22051 35751
rect 22051 35717 22060 35751
rect 22008 35708 22060 35717
rect 22100 35708 22152 35760
rect 22928 35708 22980 35760
rect 22836 35640 22888 35692
rect 23664 35708 23716 35760
rect 23940 35640 23992 35692
rect 29000 35776 29052 35828
rect 29092 35776 29144 35828
rect 29276 35776 29328 35828
rect 29736 35776 29788 35828
rect 30840 35819 30892 35828
rect 30840 35785 30849 35819
rect 30849 35785 30883 35819
rect 30883 35785 30892 35819
rect 30840 35776 30892 35785
rect 31668 35776 31720 35828
rect 32128 35776 32180 35828
rect 35624 35776 35676 35828
rect 35808 35776 35860 35828
rect 24584 35751 24636 35760
rect 24584 35717 24593 35751
rect 24593 35717 24627 35751
rect 24627 35717 24636 35751
rect 24584 35708 24636 35717
rect 27160 35708 27212 35760
rect 27528 35708 27580 35760
rect 27712 35708 27764 35760
rect 30104 35708 30156 35760
rect 24400 35640 24452 35692
rect 23296 35572 23348 35624
rect 23572 35572 23624 35624
rect 24308 35572 24360 35624
rect 25320 35572 25372 35624
rect 25780 35572 25832 35624
rect 26240 35640 26292 35692
rect 26608 35640 26660 35692
rect 28908 35683 28960 35692
rect 28908 35649 28917 35683
rect 28917 35649 28951 35683
rect 28951 35649 28960 35683
rect 28908 35640 28960 35649
rect 29276 35640 29328 35692
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 29920 35640 29972 35649
rect 30196 35683 30248 35692
rect 30196 35649 30204 35683
rect 30204 35649 30238 35683
rect 30238 35649 30248 35683
rect 30196 35640 30248 35649
rect 33140 35708 33192 35760
rect 30380 35640 30432 35692
rect 31760 35640 31812 35692
rect 32128 35640 32180 35692
rect 32956 35640 33008 35692
rect 27528 35572 27580 35624
rect 27620 35572 27672 35624
rect 28540 35615 28592 35624
rect 28540 35581 28549 35615
rect 28549 35581 28583 35615
rect 28583 35581 28592 35615
rect 28540 35572 28592 35581
rect 28632 35615 28684 35624
rect 28632 35581 28641 35615
rect 28641 35581 28675 35615
rect 28675 35581 28684 35615
rect 28632 35572 28684 35581
rect 29000 35615 29052 35624
rect 29000 35581 29009 35615
rect 29009 35581 29043 35615
rect 29043 35581 29052 35615
rect 29000 35572 29052 35581
rect 29092 35572 29144 35624
rect 26608 35547 26660 35556
rect 26608 35513 26617 35547
rect 26617 35513 26651 35547
rect 26651 35513 26660 35547
rect 26608 35504 26660 35513
rect 31208 35504 31260 35556
rect 24584 35436 24636 35488
rect 26884 35436 26936 35488
rect 29368 35436 29420 35488
rect 30012 35436 30064 35488
rect 31024 35436 31076 35488
rect 31944 35572 31996 35624
rect 32404 35572 32456 35624
rect 34152 35640 34204 35692
rect 35072 35708 35124 35760
rect 35256 35708 35308 35760
rect 37188 35708 37240 35760
rect 34888 35683 34940 35692
rect 34888 35649 34897 35683
rect 34897 35649 34931 35683
rect 34931 35649 34940 35683
rect 34888 35640 34940 35649
rect 35164 35683 35216 35692
rect 35164 35649 35173 35683
rect 35173 35649 35207 35683
rect 35207 35649 35216 35683
rect 35164 35640 35216 35649
rect 33324 35572 33376 35624
rect 34980 35615 35032 35624
rect 34980 35581 34989 35615
rect 34989 35581 35023 35615
rect 35023 35581 35032 35615
rect 34980 35572 35032 35581
rect 31484 35504 31536 35556
rect 35256 35504 35308 35556
rect 35992 35683 36044 35692
rect 35992 35649 36001 35683
rect 36001 35649 36035 35683
rect 36035 35649 36044 35683
rect 35992 35640 36044 35649
rect 36728 35640 36780 35692
rect 37648 35683 37700 35692
rect 37648 35649 37655 35683
rect 37655 35649 37700 35683
rect 37648 35640 37700 35649
rect 38476 35708 38528 35760
rect 39028 35708 39080 35760
rect 40316 35776 40368 35828
rect 41236 35776 41288 35828
rect 42616 35819 42668 35828
rect 42616 35785 42625 35819
rect 42625 35785 42659 35819
rect 42659 35785 42668 35819
rect 42616 35776 42668 35785
rect 42708 35776 42760 35828
rect 36820 35572 36872 35624
rect 35808 35504 35860 35556
rect 36176 35504 36228 35556
rect 37832 35504 37884 35556
rect 32404 35436 32456 35488
rect 32496 35479 32548 35488
rect 32496 35445 32505 35479
rect 32505 35445 32539 35479
rect 32539 35445 32548 35479
rect 32496 35436 32548 35445
rect 33876 35436 33928 35488
rect 34428 35479 34480 35488
rect 34428 35445 34437 35479
rect 34437 35445 34471 35479
rect 34471 35445 34480 35479
rect 34428 35436 34480 35445
rect 34612 35436 34664 35488
rect 35072 35436 35124 35488
rect 36636 35479 36688 35488
rect 36636 35445 36645 35479
rect 36645 35445 36679 35479
rect 36679 35445 36688 35479
rect 36636 35436 36688 35445
rect 37280 35436 37332 35488
rect 39488 35683 39540 35692
rect 39488 35649 39498 35683
rect 39498 35649 39532 35683
rect 39532 35649 39540 35683
rect 39488 35640 39540 35649
rect 39764 35683 39816 35692
rect 39764 35649 39773 35683
rect 39773 35649 39807 35683
rect 39807 35649 39816 35683
rect 39764 35640 39816 35649
rect 40408 35640 40460 35692
rect 40500 35683 40552 35692
rect 40500 35649 40509 35683
rect 40509 35649 40543 35683
rect 40543 35649 40552 35683
rect 40500 35640 40552 35649
rect 40592 35640 40644 35692
rect 40316 35572 40368 35624
rect 40868 35683 40920 35692
rect 40868 35649 40877 35683
rect 40877 35649 40911 35683
rect 40911 35649 40920 35683
rect 40868 35640 40920 35649
rect 40408 35504 40460 35556
rect 41788 35683 41840 35692
rect 41788 35649 41797 35683
rect 41797 35649 41831 35683
rect 41831 35649 41840 35683
rect 41788 35640 41840 35649
rect 41328 35572 41380 35624
rect 38200 35436 38252 35488
rect 40592 35436 40644 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6000 35232 6052 35284
rect 15384 35232 15436 35284
rect 15476 35275 15528 35284
rect 15476 35241 15485 35275
rect 15485 35241 15519 35275
rect 15519 35241 15528 35275
rect 15476 35232 15528 35241
rect 16212 35275 16264 35284
rect 16212 35241 16221 35275
rect 16221 35241 16255 35275
rect 16255 35241 16264 35275
rect 16212 35232 16264 35241
rect 20812 35232 20864 35284
rect 20904 35232 20956 35284
rect 23664 35275 23716 35284
rect 23664 35241 23673 35275
rect 23673 35241 23707 35275
rect 23707 35241 23716 35275
rect 23664 35232 23716 35241
rect 4620 35164 4672 35216
rect 2872 35096 2924 35148
rect 15016 35096 15068 35148
rect 24768 35164 24820 35216
rect 24860 35164 24912 35216
rect 26608 35232 26660 35284
rect 27712 35232 27764 35284
rect 28540 35232 28592 35284
rect 29552 35232 29604 35284
rect 30748 35232 30800 35284
rect 33416 35232 33468 35284
rect 33600 35232 33652 35284
rect 33784 35232 33836 35284
rect 33876 35232 33928 35284
rect 35808 35232 35860 35284
rect 36268 35275 36320 35284
rect 36268 35241 36277 35275
rect 36277 35241 36311 35275
rect 36311 35241 36320 35275
rect 36268 35232 36320 35241
rect 37004 35232 37056 35284
rect 28172 35164 28224 35216
rect 30104 35164 30156 35216
rect 31852 35164 31904 35216
rect 32128 35164 32180 35216
rect 32404 35164 32456 35216
rect 33968 35164 34020 35216
rect 34888 35207 34940 35216
rect 34888 35173 34897 35207
rect 34897 35173 34931 35207
rect 34931 35173 34940 35207
rect 34888 35164 34940 35173
rect 16120 35139 16172 35148
rect 16120 35105 16129 35139
rect 16129 35105 16163 35139
rect 16163 35105 16172 35139
rect 16120 35096 16172 35105
rect 14556 35028 14608 35080
rect 15108 35071 15160 35080
rect 15108 35037 15117 35071
rect 15117 35037 15151 35071
rect 15151 35037 15160 35071
rect 15108 35028 15160 35037
rect 14464 35003 14516 35012
rect 14464 34969 14473 35003
rect 14473 34969 14507 35003
rect 14507 34969 14516 35003
rect 14464 34960 14516 34969
rect 15200 34960 15252 35012
rect 13728 34935 13780 34944
rect 13728 34901 13737 34935
rect 13737 34901 13771 34935
rect 13771 34901 13780 34935
rect 13728 34892 13780 34901
rect 16304 35028 16356 35080
rect 18788 35096 18840 35148
rect 16856 35028 16908 35080
rect 17132 35028 17184 35080
rect 17960 35071 18012 35080
rect 17960 35037 17969 35071
rect 17969 35037 18003 35071
rect 18003 35037 18012 35071
rect 17960 35028 18012 35037
rect 18052 35071 18104 35080
rect 18052 35037 18061 35071
rect 18061 35037 18095 35071
rect 18095 35037 18104 35071
rect 18052 35028 18104 35037
rect 18144 35028 18196 35080
rect 18328 35071 18380 35080
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 22560 35096 22612 35148
rect 23112 35096 23164 35148
rect 23848 35096 23900 35148
rect 24584 35139 24636 35148
rect 24584 35105 24593 35139
rect 24593 35105 24627 35139
rect 24627 35105 24636 35139
rect 24584 35096 24636 35105
rect 22008 35028 22060 35080
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 22652 35028 22704 35080
rect 16028 34960 16080 35012
rect 15384 34892 15436 34944
rect 22468 35003 22520 35012
rect 22468 34969 22477 35003
rect 22477 34969 22511 35003
rect 22511 34969 22520 35003
rect 22468 34960 22520 34969
rect 22836 34960 22888 35012
rect 17132 34892 17184 34944
rect 17224 34892 17276 34944
rect 17408 34892 17460 34944
rect 18512 34892 18564 34944
rect 22100 34892 22152 34944
rect 22744 34892 22796 34944
rect 23204 35028 23256 35080
rect 23940 35028 23992 35080
rect 24860 35028 24912 35080
rect 26332 35096 26384 35148
rect 25412 35028 25464 35080
rect 25872 35028 25924 35080
rect 26056 35028 26108 35080
rect 26608 35028 26660 35080
rect 23296 34960 23348 35012
rect 24400 34960 24452 35012
rect 23572 34892 23624 34944
rect 26792 35003 26844 35012
rect 26792 34969 26801 35003
rect 26801 34969 26835 35003
rect 26835 34969 26844 35003
rect 26792 34960 26844 34969
rect 27896 35096 27948 35148
rect 33140 35096 33192 35148
rect 36176 35164 36228 35216
rect 37188 35164 37240 35216
rect 40500 35232 40552 35284
rect 36820 35096 36872 35148
rect 36912 35096 36964 35148
rect 27068 35071 27120 35080
rect 27068 35037 27076 35071
rect 27076 35037 27110 35071
rect 27110 35037 27120 35071
rect 27068 35028 27120 35037
rect 27804 35028 27856 35080
rect 28356 35071 28408 35080
rect 28356 35037 28365 35071
rect 28365 35037 28399 35071
rect 28399 35037 28408 35071
rect 28356 35028 28408 35037
rect 29276 35028 29328 35080
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30104 35071 30156 35080
rect 30104 35037 30113 35071
rect 30113 35037 30147 35071
rect 30147 35037 30156 35071
rect 30104 35028 30156 35037
rect 30288 35071 30340 35080
rect 30288 35037 30297 35071
rect 30297 35037 30331 35071
rect 30331 35037 30340 35071
rect 30288 35028 30340 35037
rect 31392 35028 31444 35080
rect 31668 35028 31720 35080
rect 32588 35028 32640 35080
rect 32680 35071 32732 35080
rect 32680 35037 32689 35071
rect 32689 35037 32723 35071
rect 32723 35037 32732 35071
rect 32680 35028 32732 35037
rect 33324 35028 33376 35080
rect 33508 35071 33560 35080
rect 33508 35037 33517 35071
rect 33517 35037 33551 35071
rect 33551 35037 33560 35071
rect 33508 35028 33560 35037
rect 33600 35071 33652 35080
rect 33600 35037 33609 35071
rect 33609 35037 33643 35071
rect 33643 35037 33652 35071
rect 33600 35028 33652 35037
rect 33784 35071 33836 35080
rect 33784 35037 33793 35071
rect 33793 35037 33827 35071
rect 33827 35037 33836 35071
rect 33784 35028 33836 35037
rect 33968 35028 34020 35080
rect 28632 35003 28684 35012
rect 28632 34969 28641 35003
rect 28641 34969 28675 35003
rect 28675 34969 28684 35003
rect 28632 34960 28684 34969
rect 29460 34960 29512 35012
rect 29828 34960 29880 35012
rect 31208 34960 31260 35012
rect 32772 34960 32824 35012
rect 33416 34960 33468 35012
rect 34520 34960 34572 35012
rect 34612 34960 34664 35012
rect 35348 35028 35400 35080
rect 35532 35071 35584 35080
rect 35532 35037 35541 35071
rect 35541 35037 35575 35071
rect 35575 35037 35584 35071
rect 35532 35028 35584 35037
rect 36728 35028 36780 35080
rect 38292 35139 38344 35148
rect 38292 35105 38301 35139
rect 38301 35105 38335 35139
rect 38335 35105 38344 35139
rect 38292 35096 38344 35105
rect 39488 35164 39540 35216
rect 40408 35096 40460 35148
rect 40592 35139 40644 35148
rect 40592 35105 40601 35139
rect 40601 35105 40635 35139
rect 40635 35105 40644 35139
rect 40592 35096 40644 35105
rect 41512 35139 41564 35148
rect 41512 35105 41521 35139
rect 41521 35105 41555 35139
rect 41555 35105 41564 35139
rect 41512 35096 41564 35105
rect 38200 35028 38252 35080
rect 38476 35028 38528 35080
rect 40132 35028 40184 35080
rect 41328 35028 41380 35080
rect 35624 34960 35676 35012
rect 36176 35003 36228 35012
rect 36176 34969 36185 35003
rect 36185 34969 36219 35003
rect 36219 34969 36228 35003
rect 36176 34960 36228 34969
rect 36360 34960 36412 35012
rect 37832 34960 37884 35012
rect 39304 34960 39356 35012
rect 39672 34960 39724 35012
rect 40960 34960 41012 35012
rect 27988 34892 28040 34944
rect 28172 34892 28224 34944
rect 34704 34892 34756 34944
rect 35808 34892 35860 34944
rect 40500 34892 40552 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 14004 34731 14056 34740
rect 14004 34697 14013 34731
rect 14013 34697 14047 34731
rect 14047 34697 14056 34731
rect 14004 34688 14056 34697
rect 16304 34731 16356 34740
rect 16304 34697 16313 34731
rect 16313 34697 16347 34731
rect 16347 34697 16356 34731
rect 16304 34688 16356 34697
rect 15016 34620 15068 34672
rect 23296 34688 23348 34740
rect 27804 34688 27856 34740
rect 29000 34731 29052 34740
rect 29000 34697 29009 34731
rect 29009 34697 29043 34731
rect 29043 34697 29052 34731
rect 29000 34688 29052 34697
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 14464 34595 14516 34604
rect 14464 34561 14473 34595
rect 14473 34561 14507 34595
rect 14507 34561 14516 34595
rect 14464 34552 14516 34561
rect 14648 34552 14700 34604
rect 15200 34552 15252 34604
rect 15568 34552 15620 34604
rect 15108 34484 15160 34536
rect 15936 34595 15988 34604
rect 15936 34561 15945 34595
rect 15945 34561 15979 34595
rect 15979 34561 15988 34595
rect 15936 34552 15988 34561
rect 16580 34552 16632 34604
rect 17132 34595 17184 34604
rect 17132 34561 17141 34595
rect 17141 34561 17175 34595
rect 17175 34561 17184 34595
rect 17132 34552 17184 34561
rect 17316 34595 17368 34604
rect 17316 34561 17325 34595
rect 17325 34561 17359 34595
rect 17359 34561 17368 34595
rect 17316 34552 17368 34561
rect 17408 34595 17460 34604
rect 17408 34561 17417 34595
rect 17417 34561 17451 34595
rect 17451 34561 17460 34595
rect 17408 34552 17460 34561
rect 17592 34552 17644 34604
rect 18420 34552 18472 34604
rect 18512 34552 18564 34604
rect 20076 34552 20128 34604
rect 22928 34620 22980 34672
rect 26240 34620 26292 34672
rect 27344 34663 27396 34672
rect 27344 34629 27353 34663
rect 27353 34629 27387 34663
rect 27387 34629 27396 34663
rect 27344 34620 27396 34629
rect 29092 34620 29144 34672
rect 16764 34484 16816 34536
rect 22284 34595 22336 34604
rect 22284 34561 22293 34595
rect 22293 34561 22327 34595
rect 22327 34561 22336 34595
rect 22284 34552 22336 34561
rect 23572 34552 23624 34604
rect 24768 34552 24820 34604
rect 25136 34552 25188 34604
rect 25596 34595 25648 34604
rect 25596 34561 25605 34595
rect 25605 34561 25639 34595
rect 25639 34561 25648 34595
rect 25596 34552 25648 34561
rect 25688 34595 25740 34604
rect 25688 34561 25697 34595
rect 25697 34561 25731 34595
rect 25731 34561 25740 34595
rect 25688 34552 25740 34561
rect 25872 34595 25924 34604
rect 25872 34561 25881 34595
rect 25881 34561 25915 34595
rect 25915 34561 25924 34595
rect 25872 34552 25924 34561
rect 27988 34595 28040 34604
rect 27988 34561 27997 34595
rect 27997 34561 28031 34595
rect 28031 34561 28040 34595
rect 27988 34552 28040 34561
rect 28172 34552 28224 34604
rect 28356 34595 28408 34604
rect 28356 34561 28365 34595
rect 28365 34561 28399 34595
rect 28399 34561 28408 34595
rect 28356 34552 28408 34561
rect 31668 34688 31720 34740
rect 31760 34731 31812 34740
rect 31760 34697 31769 34731
rect 31769 34697 31803 34731
rect 31803 34697 31812 34731
rect 31760 34688 31812 34697
rect 30840 34620 30892 34672
rect 20628 34484 20680 34536
rect 20812 34484 20864 34536
rect 23296 34484 23348 34536
rect 20536 34459 20588 34468
rect 20536 34425 20545 34459
rect 20545 34425 20579 34459
rect 20579 34425 20588 34459
rect 20536 34416 20588 34425
rect 20720 34416 20772 34468
rect 23664 34484 23716 34536
rect 24124 34484 24176 34536
rect 25228 34484 25280 34536
rect 25504 34484 25556 34536
rect 26056 34484 26108 34536
rect 27436 34484 27488 34536
rect 29368 34595 29420 34604
rect 29368 34561 29377 34595
rect 29377 34561 29411 34595
rect 29411 34561 29420 34595
rect 29368 34552 29420 34561
rect 30012 34552 30064 34604
rect 29276 34527 29328 34536
rect 29276 34493 29285 34527
rect 29285 34493 29319 34527
rect 29319 34493 29328 34527
rect 29276 34484 29328 34493
rect 29736 34484 29788 34536
rect 33508 34688 33560 34740
rect 33968 34688 34020 34740
rect 34060 34620 34112 34672
rect 35348 34688 35400 34740
rect 38568 34688 38620 34740
rect 42708 34688 42760 34740
rect 32772 34552 32824 34604
rect 38108 34620 38160 34672
rect 40316 34663 40368 34672
rect 40316 34629 40325 34663
rect 40325 34629 40359 34663
rect 40359 34629 40368 34663
rect 40316 34620 40368 34629
rect 40500 34620 40552 34672
rect 13728 34348 13780 34400
rect 20812 34348 20864 34400
rect 22560 34391 22612 34400
rect 22560 34357 22569 34391
rect 22569 34357 22603 34391
rect 22603 34357 22612 34391
rect 22560 34348 22612 34357
rect 23296 34348 23348 34400
rect 28540 34416 28592 34468
rect 26516 34391 26568 34400
rect 26516 34357 26525 34391
rect 26525 34357 26559 34391
rect 26559 34357 26568 34391
rect 26516 34348 26568 34357
rect 32220 34484 32272 34536
rect 32680 34416 32732 34468
rect 33048 34527 33100 34536
rect 33048 34493 33057 34527
rect 33057 34493 33091 34527
rect 33091 34493 33100 34527
rect 33048 34484 33100 34493
rect 34244 34484 34296 34536
rect 36176 34552 36228 34604
rect 36452 34595 36504 34604
rect 36452 34561 36461 34595
rect 36461 34561 36495 34595
rect 36495 34561 36504 34595
rect 36452 34552 36504 34561
rect 36084 34484 36136 34536
rect 36728 34552 36780 34604
rect 36820 34595 36872 34604
rect 36820 34561 36829 34595
rect 36829 34561 36863 34595
rect 36863 34561 36872 34595
rect 36820 34552 36872 34561
rect 37556 34552 37608 34604
rect 37648 34595 37700 34604
rect 37648 34561 37657 34595
rect 37657 34561 37691 34595
rect 37691 34561 37700 34595
rect 37648 34552 37700 34561
rect 37740 34595 37792 34604
rect 37740 34561 37749 34595
rect 37749 34561 37783 34595
rect 37783 34561 37792 34595
rect 37740 34552 37792 34561
rect 37924 34552 37976 34604
rect 39028 34552 39080 34604
rect 40224 34552 40276 34604
rect 42800 34595 42852 34604
rect 42800 34561 42809 34595
rect 42809 34561 42843 34595
rect 42843 34561 42852 34595
rect 42800 34552 42852 34561
rect 38292 34484 38344 34536
rect 30840 34348 30892 34400
rect 33692 34348 33744 34400
rect 38844 34416 38896 34468
rect 37188 34348 37240 34400
rect 37280 34348 37332 34400
rect 37556 34348 37608 34400
rect 38476 34391 38528 34400
rect 38476 34357 38485 34391
rect 38485 34357 38519 34391
rect 38519 34357 38528 34391
rect 38476 34348 38528 34357
rect 40132 34484 40184 34536
rect 42708 34527 42760 34536
rect 42708 34493 42717 34527
rect 42717 34493 42751 34527
rect 42751 34493 42760 34527
rect 42708 34484 42760 34493
rect 43076 34416 43128 34468
rect 40960 34348 41012 34400
rect 42156 34348 42208 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 13820 34144 13872 34196
rect 14464 34187 14516 34196
rect 14464 34153 14473 34187
rect 14473 34153 14507 34187
rect 14507 34153 14516 34187
rect 14464 34144 14516 34153
rect 16856 34187 16908 34196
rect 16856 34153 16865 34187
rect 16865 34153 16899 34187
rect 16899 34153 16908 34187
rect 16856 34144 16908 34153
rect 17316 34144 17368 34196
rect 22192 34187 22244 34196
rect 22192 34153 22201 34187
rect 22201 34153 22235 34187
rect 22235 34153 22244 34187
rect 22192 34144 22244 34153
rect 24216 34144 24268 34196
rect 26792 34144 26844 34196
rect 27068 34144 27120 34196
rect 29092 34187 29144 34196
rect 29092 34153 29101 34187
rect 29101 34153 29135 34187
rect 29135 34153 29144 34187
rect 29092 34144 29144 34153
rect 29276 34144 29328 34196
rect 30748 34144 30800 34196
rect 32220 34144 32272 34196
rect 32496 34144 32548 34196
rect 32864 34144 32916 34196
rect 35992 34144 36044 34196
rect 39028 34144 39080 34196
rect 13268 34076 13320 34128
rect 20536 34119 20588 34128
rect 20536 34085 20545 34119
rect 20545 34085 20579 34119
rect 20579 34085 20588 34119
rect 20536 34076 20588 34085
rect 22008 34076 22060 34128
rect 17040 34008 17092 34060
rect 18144 34008 18196 34060
rect 21088 34008 21140 34060
rect 13176 33983 13228 33992
rect 13176 33949 13185 33983
rect 13185 33949 13219 33983
rect 13219 33949 13228 33983
rect 13176 33940 13228 33949
rect 13268 33983 13320 33992
rect 13268 33949 13277 33983
rect 13277 33949 13311 33983
rect 13311 33949 13320 33983
rect 13268 33940 13320 33949
rect 13544 33983 13596 33992
rect 13544 33949 13553 33983
rect 13553 33949 13587 33983
rect 13587 33949 13596 33983
rect 13544 33940 13596 33949
rect 14280 33983 14332 33992
rect 14280 33949 14289 33983
rect 14289 33949 14323 33983
rect 14323 33949 14332 33983
rect 14280 33940 14332 33949
rect 14648 33983 14700 33992
rect 14648 33949 14657 33983
rect 14657 33949 14691 33983
rect 14691 33949 14700 33983
rect 14648 33940 14700 33949
rect 15936 33940 15988 33992
rect 16672 33983 16724 33992
rect 16672 33949 16681 33983
rect 16681 33949 16715 33983
rect 16715 33949 16724 33983
rect 16672 33940 16724 33949
rect 16764 33983 16816 33992
rect 16764 33949 16773 33983
rect 16773 33949 16807 33983
rect 16807 33949 16816 33983
rect 16764 33940 16816 33949
rect 17960 33983 18012 33992
rect 17960 33949 17969 33983
rect 17969 33949 18003 33983
rect 18003 33949 18012 33983
rect 17960 33940 18012 33949
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 18236 33983 18288 33992
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 18788 33940 18840 33992
rect 22928 34051 22980 34060
rect 22928 34017 22937 34051
rect 22937 34017 22971 34051
rect 22971 34017 22980 34051
rect 22928 34008 22980 34017
rect 23388 34008 23440 34060
rect 26516 34076 26568 34128
rect 28172 34076 28224 34128
rect 25504 34008 25556 34060
rect 13820 33804 13872 33856
rect 15108 33872 15160 33924
rect 15752 33804 15804 33856
rect 16396 33872 16448 33924
rect 16580 33872 16632 33924
rect 19340 33872 19392 33924
rect 20904 33915 20956 33924
rect 20904 33881 20913 33915
rect 20913 33881 20947 33915
rect 20947 33881 20956 33915
rect 20904 33872 20956 33881
rect 16856 33804 16908 33856
rect 19984 33847 20036 33856
rect 19984 33813 19993 33847
rect 19993 33813 20027 33847
rect 20027 33813 20036 33847
rect 19984 33804 20036 33813
rect 20444 33847 20496 33856
rect 20444 33813 20453 33847
rect 20453 33813 20487 33847
rect 20487 33813 20496 33847
rect 20444 33804 20496 33813
rect 22192 33872 22244 33924
rect 22560 33872 22612 33924
rect 23204 33872 23256 33924
rect 23296 33872 23348 33924
rect 23572 33872 23624 33924
rect 24400 33940 24452 33992
rect 25320 33983 25372 33992
rect 25320 33949 25324 33983
rect 25324 33949 25358 33983
rect 25358 33949 25372 33983
rect 25320 33940 25372 33949
rect 23848 33872 23900 33924
rect 24400 33804 24452 33856
rect 25228 33872 25280 33924
rect 26700 34008 26752 34060
rect 25872 33940 25924 33992
rect 27804 34008 27856 34060
rect 27068 33983 27120 33992
rect 27068 33949 27077 33983
rect 27077 33949 27111 33983
rect 27111 33949 27120 33983
rect 27068 33940 27120 33949
rect 27712 33983 27764 33992
rect 27712 33949 27730 33983
rect 27730 33949 27764 33983
rect 27712 33940 27764 33949
rect 27896 33983 27948 33992
rect 27896 33949 27905 33983
rect 27905 33949 27939 33983
rect 27939 33949 27948 33983
rect 27896 33940 27948 33949
rect 27988 33983 28040 33992
rect 27988 33949 28033 33983
rect 28033 33949 28040 33983
rect 27988 33940 28040 33949
rect 28816 34008 28868 34060
rect 29092 34008 29144 34060
rect 30104 34076 30156 34128
rect 29460 33940 29512 33992
rect 29552 33940 29604 33992
rect 30104 33940 30156 33992
rect 31484 33940 31536 33992
rect 31852 33940 31904 33992
rect 32588 33940 32640 33992
rect 32864 33940 32916 33992
rect 34428 33940 34480 33992
rect 34520 33940 34572 33992
rect 35808 33940 35860 33992
rect 26056 33872 26108 33924
rect 28724 33872 28776 33924
rect 28816 33915 28868 33924
rect 28816 33881 28825 33915
rect 28825 33881 28859 33915
rect 28859 33881 28868 33915
rect 28816 33872 28868 33881
rect 28908 33872 28960 33924
rect 32956 33872 33008 33924
rect 33600 33872 33652 33924
rect 26424 33847 26476 33856
rect 26424 33813 26433 33847
rect 26433 33813 26467 33847
rect 26467 33813 26476 33847
rect 26424 33804 26476 33813
rect 26516 33804 26568 33856
rect 27620 33804 27672 33856
rect 30012 33804 30064 33856
rect 30472 33847 30524 33856
rect 30472 33813 30481 33847
rect 30481 33813 30515 33847
rect 30515 33813 30524 33847
rect 30472 33804 30524 33813
rect 30932 33804 30984 33856
rect 33508 33804 33560 33856
rect 35348 33872 35400 33924
rect 37188 34076 37240 34128
rect 38016 34076 38068 34128
rect 40960 34144 41012 34196
rect 41052 34144 41104 34196
rect 41420 34119 41472 34128
rect 41420 34085 41429 34119
rect 41429 34085 41463 34119
rect 41463 34085 41472 34119
rect 41420 34076 41472 34085
rect 36912 33940 36964 33992
rect 37648 33940 37700 33992
rect 38384 33940 38436 33992
rect 39120 33983 39172 33992
rect 39120 33949 39129 33983
rect 39129 33949 39163 33983
rect 39163 33949 39172 33983
rect 39120 33940 39172 33949
rect 39764 33940 39816 33992
rect 40040 33983 40092 33992
rect 40040 33949 40049 33983
rect 40049 33949 40083 33983
rect 40083 33949 40092 33983
rect 40040 33940 40092 33949
rect 41328 33940 41380 33992
rect 43168 33940 43220 33992
rect 37096 33872 37148 33924
rect 36452 33804 36504 33856
rect 37188 33804 37240 33856
rect 38016 33872 38068 33924
rect 37924 33847 37976 33856
rect 37924 33813 37933 33847
rect 37933 33813 37967 33847
rect 37967 33813 37976 33847
rect 37924 33804 37976 33813
rect 38108 33804 38160 33856
rect 38936 33872 38988 33924
rect 38384 33804 38436 33856
rect 38476 33804 38528 33856
rect 39396 33804 39448 33856
rect 42156 33872 42208 33924
rect 42800 33872 42852 33924
rect 42984 33915 43036 33924
rect 42984 33881 43002 33915
rect 43002 33881 43036 33915
rect 42984 33872 43036 33881
rect 41880 33847 41932 33856
rect 41880 33813 41889 33847
rect 41889 33813 41923 33847
rect 41923 33813 41932 33847
rect 41880 33804 41932 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 13544 33600 13596 33652
rect 13820 33600 13872 33652
rect 15108 33643 15160 33652
rect 15108 33609 15117 33643
rect 15117 33609 15151 33643
rect 15151 33609 15160 33643
rect 15108 33600 15160 33609
rect 15568 33643 15620 33652
rect 15568 33609 15577 33643
rect 15577 33609 15611 33643
rect 15611 33609 15620 33643
rect 15568 33600 15620 33609
rect 15936 33600 15988 33652
rect 16580 33600 16632 33652
rect 19984 33600 20036 33652
rect 23572 33600 23624 33652
rect 24216 33600 24268 33652
rect 24860 33600 24912 33652
rect 25688 33600 25740 33652
rect 28264 33600 28316 33652
rect 28540 33600 28592 33652
rect 31208 33600 31260 33652
rect 31300 33600 31352 33652
rect 15752 33507 15804 33516
rect 15752 33473 15761 33507
rect 15761 33473 15795 33507
rect 15795 33473 15804 33507
rect 15752 33464 15804 33473
rect 16948 33464 17000 33516
rect 18052 33507 18104 33516
rect 18052 33473 18061 33507
rect 18061 33473 18095 33507
rect 18095 33473 18104 33507
rect 18052 33464 18104 33473
rect 20168 33464 20220 33516
rect 24768 33532 24820 33584
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 22560 33507 22612 33516
rect 22560 33473 22569 33507
rect 22569 33473 22603 33507
rect 22603 33473 22612 33507
rect 22560 33464 22612 33473
rect 23572 33507 23624 33516
rect 23572 33473 23581 33507
rect 23581 33473 23615 33507
rect 23615 33473 23624 33507
rect 23572 33464 23624 33473
rect 24308 33507 24360 33516
rect 24308 33473 24317 33507
rect 24317 33473 24351 33507
rect 24351 33473 24360 33507
rect 24308 33464 24360 33473
rect 25872 33532 25924 33584
rect 27528 33532 27580 33584
rect 29552 33532 29604 33584
rect 30748 33532 30800 33584
rect 31024 33532 31076 33584
rect 31760 33532 31812 33584
rect 32404 33643 32456 33652
rect 32404 33609 32413 33643
rect 32413 33609 32447 33643
rect 32447 33609 32456 33643
rect 32404 33600 32456 33609
rect 33692 33600 33744 33652
rect 33784 33600 33836 33652
rect 37740 33600 37792 33652
rect 38936 33643 38988 33652
rect 38936 33609 38945 33643
rect 38945 33609 38979 33643
rect 38979 33609 38988 33643
rect 38936 33600 38988 33609
rect 39028 33600 39080 33652
rect 41604 33600 41656 33652
rect 43076 33600 43128 33652
rect 25136 33507 25188 33516
rect 25136 33473 25145 33507
rect 25145 33473 25179 33507
rect 25179 33473 25188 33507
rect 25136 33464 25188 33473
rect 16488 33396 16540 33448
rect 17684 33396 17736 33448
rect 18696 33396 18748 33448
rect 19248 33439 19300 33448
rect 19248 33405 19257 33439
rect 19257 33405 19291 33439
rect 19291 33405 19300 33439
rect 19248 33396 19300 33405
rect 19616 33439 19668 33448
rect 19616 33405 19625 33439
rect 19625 33405 19659 33439
rect 19659 33405 19668 33439
rect 19616 33396 19668 33405
rect 20260 33439 20312 33448
rect 20260 33405 20269 33439
rect 20269 33405 20303 33439
rect 20303 33405 20312 33439
rect 20260 33396 20312 33405
rect 14372 33260 14424 33312
rect 17224 33303 17276 33312
rect 17224 33269 17233 33303
rect 17233 33269 17267 33303
rect 17267 33269 17276 33303
rect 17224 33260 17276 33269
rect 19156 33260 19208 33312
rect 19340 33260 19392 33312
rect 20352 33260 20404 33312
rect 20720 33328 20772 33380
rect 23756 33396 23808 33448
rect 24584 33396 24636 33448
rect 24952 33396 25004 33448
rect 25320 33507 25372 33516
rect 25320 33473 25329 33507
rect 25329 33473 25363 33507
rect 25363 33473 25372 33507
rect 25320 33464 25372 33473
rect 22652 33328 22704 33380
rect 23480 33328 23532 33380
rect 21272 33260 21324 33312
rect 22468 33303 22520 33312
rect 22468 33269 22477 33303
rect 22477 33269 22511 33303
rect 22511 33269 22520 33303
rect 22468 33260 22520 33269
rect 23388 33260 23440 33312
rect 24492 33328 24544 33380
rect 25044 33328 25096 33380
rect 26516 33464 26568 33516
rect 27712 33396 27764 33448
rect 27988 33396 28040 33448
rect 28908 33464 28960 33516
rect 29644 33507 29696 33516
rect 29644 33473 29648 33507
rect 29648 33473 29682 33507
rect 29682 33473 29696 33507
rect 29644 33464 29696 33473
rect 30012 33507 30064 33516
rect 28264 33439 28316 33448
rect 28264 33405 28273 33439
rect 28273 33405 28307 33439
rect 28307 33405 28316 33439
rect 28264 33396 28316 33405
rect 29736 33396 29788 33448
rect 30012 33473 30020 33507
rect 30020 33473 30054 33507
rect 30054 33473 30064 33507
rect 30012 33464 30064 33473
rect 30104 33507 30156 33516
rect 30104 33473 30113 33507
rect 30113 33473 30147 33507
rect 30147 33473 30156 33507
rect 30104 33464 30156 33473
rect 30288 33464 30340 33516
rect 37648 33532 37700 33584
rect 38568 33532 38620 33584
rect 41052 33532 41104 33584
rect 31208 33396 31260 33448
rect 32772 33507 32824 33516
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 33876 33464 33928 33516
rect 34060 33507 34112 33516
rect 34060 33473 34069 33507
rect 34069 33473 34103 33507
rect 34103 33473 34112 33507
rect 34060 33464 34112 33473
rect 32588 33396 32640 33448
rect 32864 33396 32916 33448
rect 33600 33396 33652 33448
rect 34704 33464 34756 33516
rect 35256 33439 35308 33448
rect 35256 33405 35265 33439
rect 35265 33405 35299 33439
rect 35299 33405 35308 33439
rect 35256 33396 35308 33405
rect 31024 33328 31076 33380
rect 25412 33260 25464 33312
rect 26332 33260 26384 33312
rect 27344 33260 27396 33312
rect 27712 33260 27764 33312
rect 28540 33260 28592 33312
rect 29000 33303 29052 33312
rect 29000 33269 29009 33303
rect 29009 33269 29043 33303
rect 29043 33269 29052 33303
rect 29000 33260 29052 33269
rect 29460 33303 29512 33312
rect 29460 33269 29469 33303
rect 29469 33269 29503 33303
rect 29503 33269 29512 33303
rect 29460 33260 29512 33269
rect 29736 33260 29788 33312
rect 30932 33260 30984 33312
rect 31116 33303 31168 33312
rect 31116 33269 31125 33303
rect 31125 33269 31159 33303
rect 31159 33269 31168 33303
rect 31116 33260 31168 33269
rect 31484 33260 31536 33312
rect 32680 33260 32732 33312
rect 32956 33260 33008 33312
rect 33140 33260 33192 33312
rect 33968 33260 34020 33312
rect 36636 33464 36688 33516
rect 37004 33464 37056 33516
rect 37556 33464 37608 33516
rect 38292 33464 38344 33516
rect 35900 33396 35952 33448
rect 39396 33507 39448 33516
rect 39396 33473 39405 33507
rect 39405 33473 39439 33507
rect 39439 33473 39448 33507
rect 39396 33464 39448 33473
rect 39948 33464 40000 33516
rect 40776 33464 40828 33516
rect 40868 33507 40920 33516
rect 40868 33473 40877 33507
rect 40877 33473 40911 33507
rect 40911 33473 40920 33507
rect 40868 33464 40920 33473
rect 41420 33464 41472 33516
rect 42984 33532 43036 33584
rect 42800 33507 42852 33516
rect 42800 33473 42809 33507
rect 42809 33473 42843 33507
rect 42843 33473 42852 33507
rect 42800 33464 42852 33473
rect 36084 33328 36136 33380
rect 37464 33328 37516 33380
rect 37740 33328 37792 33380
rect 39488 33396 39540 33448
rect 37648 33260 37700 33312
rect 38476 33260 38528 33312
rect 38752 33303 38804 33312
rect 38752 33269 38761 33303
rect 38761 33269 38795 33303
rect 38795 33269 38804 33303
rect 38752 33260 38804 33269
rect 39028 33260 39080 33312
rect 41604 33328 41656 33380
rect 41880 33303 41932 33312
rect 41880 33269 41889 33303
rect 41889 33269 41923 33303
rect 41923 33269 41932 33303
rect 41880 33260 41932 33269
rect 42432 33260 42484 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 12624 33099 12676 33108
rect 12624 33065 12633 33099
rect 12633 33065 12667 33099
rect 12667 33065 12676 33099
rect 12624 33056 12676 33065
rect 13268 33056 13320 33108
rect 14372 33099 14424 33108
rect 14372 33065 14381 33099
rect 14381 33065 14415 33099
rect 14415 33065 14424 33099
rect 14372 33056 14424 33065
rect 16488 33099 16540 33108
rect 16488 33065 16497 33099
rect 16497 33065 16531 33099
rect 16531 33065 16540 33099
rect 16488 33056 16540 33065
rect 16672 33056 16724 33108
rect 18052 33056 18104 33108
rect 18328 33056 18380 33108
rect 18696 33031 18748 33040
rect 18696 32997 18705 33031
rect 18705 32997 18739 33031
rect 18739 32997 18748 33031
rect 18696 32988 18748 32997
rect 20260 33056 20312 33108
rect 24124 33056 24176 33108
rect 24308 33056 24360 33108
rect 25228 33056 25280 33108
rect 27068 33099 27120 33108
rect 27068 33065 27077 33099
rect 27077 33065 27111 33099
rect 27111 33065 27120 33099
rect 27068 33056 27120 33065
rect 28816 33099 28868 33108
rect 28816 33065 28825 33099
rect 28825 33065 28859 33099
rect 28859 33065 28868 33099
rect 28816 33056 28868 33065
rect 30380 33056 30432 33108
rect 30932 33056 30984 33108
rect 34336 33056 34388 33108
rect 35716 33056 35768 33108
rect 16212 32920 16264 32972
rect 16304 32920 16356 32972
rect 19616 32920 19668 32972
rect 20444 32963 20496 32972
rect 20444 32929 20453 32963
rect 20453 32929 20487 32963
rect 20487 32929 20496 32963
rect 20444 32920 20496 32929
rect 12624 32895 12676 32904
rect 12624 32861 12633 32895
rect 12633 32861 12667 32895
rect 12667 32861 12676 32895
rect 12624 32852 12676 32861
rect 13360 32895 13412 32904
rect 13360 32861 13369 32895
rect 13369 32861 13403 32895
rect 13403 32861 13412 32895
rect 13360 32852 13412 32861
rect 13912 32852 13964 32904
rect 13084 32827 13136 32836
rect 13084 32793 13093 32827
rect 13093 32793 13127 32827
rect 13127 32793 13136 32827
rect 13084 32784 13136 32793
rect 14556 32827 14608 32836
rect 14556 32793 14565 32827
rect 14565 32793 14599 32827
rect 14599 32793 14608 32827
rect 14556 32784 14608 32793
rect 16396 32895 16448 32904
rect 16396 32861 16405 32895
rect 16405 32861 16439 32895
rect 16439 32861 16448 32895
rect 16396 32852 16448 32861
rect 17224 32852 17276 32904
rect 20720 32852 20772 32904
rect 13268 32759 13320 32768
rect 13268 32725 13277 32759
rect 13277 32725 13311 32759
rect 13311 32725 13320 32759
rect 13268 32716 13320 32725
rect 14096 32716 14148 32768
rect 15384 32716 15436 32768
rect 15936 32716 15988 32768
rect 17684 32827 17736 32836
rect 17684 32793 17693 32827
rect 17693 32793 17727 32827
rect 17727 32793 17736 32827
rect 17684 32784 17736 32793
rect 21916 32988 21968 33040
rect 29920 32988 29972 33040
rect 31760 33031 31812 33040
rect 31760 32997 31769 33031
rect 31769 32997 31803 33031
rect 31803 32997 31812 33031
rect 31760 32988 31812 32997
rect 32956 33031 33008 33040
rect 32956 32997 32965 33031
rect 32965 32997 32999 33031
rect 32999 32997 33008 33031
rect 32956 32988 33008 32997
rect 34612 32988 34664 33040
rect 35900 32988 35952 33040
rect 36820 33056 36872 33108
rect 37648 33056 37700 33108
rect 37740 33099 37792 33108
rect 37740 33065 37749 33099
rect 37749 33065 37783 33099
rect 37783 33065 37792 33099
rect 37740 33056 37792 33065
rect 40960 32988 41012 33040
rect 21272 32920 21324 32972
rect 21640 32963 21692 32972
rect 21640 32929 21649 32963
rect 21649 32929 21683 32963
rect 21683 32929 21692 32963
rect 21640 32920 21692 32929
rect 23756 32920 23808 32972
rect 22100 32852 22152 32904
rect 22468 32895 22520 32904
rect 22468 32861 22477 32895
rect 22477 32861 22511 32895
rect 22511 32861 22520 32895
rect 22468 32852 22520 32861
rect 22560 32895 22612 32904
rect 22560 32861 22569 32895
rect 22569 32861 22603 32895
rect 22603 32861 22612 32895
rect 22560 32852 22612 32861
rect 22652 32895 22704 32904
rect 22652 32861 22661 32895
rect 22661 32861 22695 32895
rect 22695 32861 22704 32895
rect 22652 32852 22704 32861
rect 22836 32895 22888 32904
rect 22836 32861 22845 32895
rect 22845 32861 22879 32895
rect 22879 32861 22888 32895
rect 22836 32852 22888 32861
rect 23848 32852 23900 32904
rect 25136 32920 25188 32972
rect 26148 32920 26200 32972
rect 25688 32852 25740 32904
rect 26332 32852 26384 32904
rect 27804 32920 27856 32972
rect 27988 32920 28040 32972
rect 28540 32920 28592 32972
rect 20904 32784 20956 32836
rect 21732 32784 21784 32836
rect 25320 32784 25372 32836
rect 19984 32716 20036 32768
rect 20352 32759 20404 32768
rect 20352 32725 20361 32759
rect 20361 32725 20395 32759
rect 20395 32725 20404 32759
rect 20352 32716 20404 32725
rect 22376 32716 22428 32768
rect 25044 32716 25096 32768
rect 26792 32827 26844 32836
rect 26792 32793 26801 32827
rect 26801 32793 26835 32827
rect 26835 32793 26844 32827
rect 26792 32784 26844 32793
rect 27436 32716 27488 32768
rect 27712 32895 27764 32904
rect 27712 32861 27721 32895
rect 27721 32861 27755 32895
rect 27755 32861 27764 32895
rect 27712 32852 27764 32861
rect 28816 32784 28868 32836
rect 29460 32852 29512 32904
rect 29920 32852 29972 32904
rect 35348 32920 35400 32972
rect 35624 32963 35676 32972
rect 35624 32929 35633 32963
rect 35633 32929 35667 32963
rect 35667 32929 35676 32963
rect 35624 32920 35676 32929
rect 35992 32920 36044 32972
rect 37648 32920 37700 32972
rect 41052 32920 41104 32972
rect 41328 32963 41380 32972
rect 41328 32929 41337 32963
rect 41337 32929 41371 32963
rect 41371 32929 41380 32963
rect 41328 32920 41380 32929
rect 41604 32963 41656 32972
rect 41604 32929 41613 32963
rect 41613 32929 41647 32963
rect 41647 32929 41656 32963
rect 41604 32920 41656 32929
rect 42800 32920 42852 32972
rect 29276 32784 29328 32836
rect 30288 32852 30340 32904
rect 30564 32895 30616 32904
rect 30564 32861 30573 32895
rect 30573 32861 30607 32895
rect 30607 32861 30616 32895
rect 30564 32852 30616 32861
rect 30748 32895 30800 32904
rect 30748 32861 30757 32895
rect 30757 32861 30791 32895
rect 30791 32861 30800 32895
rect 30748 32852 30800 32861
rect 31944 32895 31996 32904
rect 31944 32861 31953 32895
rect 31953 32861 31987 32895
rect 31987 32861 31996 32895
rect 31944 32852 31996 32861
rect 32036 32895 32088 32904
rect 32036 32861 32045 32895
rect 32045 32861 32079 32895
rect 32079 32861 32088 32895
rect 32036 32852 32088 32861
rect 32220 32852 32272 32904
rect 32312 32895 32364 32904
rect 32312 32861 32321 32895
rect 32321 32861 32355 32895
rect 32355 32861 32364 32895
rect 32312 32852 32364 32861
rect 32680 32852 32732 32904
rect 33968 32895 34020 32904
rect 33968 32861 33977 32895
rect 33977 32861 34011 32895
rect 34011 32861 34020 32895
rect 33968 32852 34020 32861
rect 30196 32784 30248 32836
rect 32404 32784 32456 32836
rect 33784 32827 33836 32836
rect 33784 32793 33793 32827
rect 33793 32793 33827 32827
rect 33827 32793 33836 32827
rect 33784 32784 33836 32793
rect 35808 32852 35860 32904
rect 36084 32895 36136 32904
rect 36084 32861 36093 32895
rect 36093 32861 36127 32895
rect 36127 32861 36136 32895
rect 36084 32852 36136 32861
rect 37372 32895 37424 32904
rect 37372 32861 37381 32895
rect 37381 32861 37415 32895
rect 37415 32861 37424 32895
rect 37372 32852 37424 32861
rect 29000 32716 29052 32768
rect 31208 32759 31260 32768
rect 31208 32725 31217 32759
rect 31217 32725 31251 32759
rect 31251 32725 31260 32759
rect 31208 32716 31260 32725
rect 33968 32716 34020 32768
rect 34060 32716 34112 32768
rect 39396 32895 39448 32904
rect 39396 32861 39405 32895
rect 39405 32861 39439 32895
rect 39439 32861 39448 32895
rect 39396 32852 39448 32861
rect 40040 32895 40092 32904
rect 40040 32861 40049 32895
rect 40049 32861 40083 32895
rect 40083 32861 40092 32895
rect 40040 32852 40092 32861
rect 39948 32784 40000 32836
rect 40776 32852 40828 32904
rect 40868 32895 40920 32904
rect 40868 32861 40877 32895
rect 40877 32861 40911 32895
rect 40911 32861 40920 32895
rect 40868 32852 40920 32861
rect 42708 32852 42760 32904
rect 37648 32716 37700 32768
rect 38200 32759 38252 32768
rect 38200 32725 38209 32759
rect 38209 32725 38243 32759
rect 38243 32725 38252 32759
rect 38200 32716 38252 32725
rect 39304 32759 39356 32768
rect 39304 32725 39313 32759
rect 39313 32725 39347 32759
rect 39347 32725 39356 32759
rect 39304 32716 39356 32725
rect 41144 32784 41196 32836
rect 40500 32716 40552 32768
rect 40684 32716 40736 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15200 32512 15252 32564
rect 16396 32512 16448 32564
rect 13176 32444 13228 32496
rect 14280 32444 14332 32496
rect 18604 32512 18656 32564
rect 20168 32555 20220 32564
rect 20168 32521 20177 32555
rect 20177 32521 20211 32555
rect 20211 32521 20220 32555
rect 20168 32512 20220 32521
rect 20904 32512 20956 32564
rect 22100 32512 22152 32564
rect 22836 32512 22888 32564
rect 13912 32419 13964 32428
rect 13912 32385 13921 32419
rect 13921 32385 13955 32419
rect 13955 32385 13964 32419
rect 13912 32376 13964 32385
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 15016 32376 15068 32428
rect 14464 32240 14516 32292
rect 24860 32512 24912 32564
rect 24952 32512 25004 32564
rect 26240 32512 26292 32564
rect 27160 32555 27212 32564
rect 27160 32521 27169 32555
rect 27169 32521 27203 32555
rect 27203 32521 27212 32555
rect 27160 32512 27212 32521
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 17868 32419 17920 32428
rect 17868 32385 17877 32419
rect 17877 32385 17911 32419
rect 17911 32385 17920 32419
rect 17868 32376 17920 32385
rect 18328 32376 18380 32428
rect 18604 32376 18656 32428
rect 18972 32419 19024 32428
rect 18972 32385 18981 32419
rect 18981 32385 19015 32419
rect 19015 32385 19024 32419
rect 18972 32376 19024 32385
rect 19064 32419 19116 32428
rect 19064 32385 19073 32419
rect 19073 32385 19107 32419
rect 19107 32385 19116 32419
rect 19064 32376 19116 32385
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 19340 32376 19392 32385
rect 15936 32308 15988 32360
rect 16212 32308 16264 32360
rect 24676 32444 24728 32496
rect 16488 32240 16540 32292
rect 19248 32240 19300 32292
rect 20260 32240 20312 32292
rect 20536 32308 20588 32360
rect 22468 32351 22520 32360
rect 22468 32317 22477 32351
rect 22477 32317 22511 32351
rect 22511 32317 22520 32351
rect 22468 32308 22520 32317
rect 23940 32419 23992 32428
rect 23940 32385 23949 32419
rect 23949 32385 23983 32419
rect 23983 32385 23992 32419
rect 23940 32376 23992 32385
rect 24032 32419 24084 32428
rect 24032 32385 24041 32419
rect 24041 32385 24075 32419
rect 24075 32385 24084 32419
rect 24032 32376 24084 32385
rect 24308 32419 24360 32428
rect 24308 32385 24317 32419
rect 24317 32385 24351 32419
rect 24351 32385 24360 32419
rect 24308 32376 24360 32385
rect 24584 32376 24636 32428
rect 24952 32419 25004 32428
rect 24952 32385 24961 32419
rect 24961 32385 24995 32419
rect 24995 32385 25004 32419
rect 24952 32376 25004 32385
rect 25228 32376 25280 32428
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 25872 32376 25924 32428
rect 27252 32444 27304 32496
rect 26976 32376 27028 32428
rect 29000 32512 29052 32564
rect 28264 32444 28316 32496
rect 28540 32444 28592 32496
rect 29276 32512 29328 32564
rect 29552 32512 29604 32564
rect 13084 32172 13136 32224
rect 13452 32172 13504 32224
rect 15200 32172 15252 32224
rect 16948 32172 17000 32224
rect 18696 32172 18748 32224
rect 22560 32215 22612 32224
rect 22560 32181 22569 32215
rect 22569 32181 22603 32215
rect 22603 32181 22612 32215
rect 22560 32172 22612 32181
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 23756 32215 23808 32224
rect 23756 32181 23765 32215
rect 23765 32181 23799 32215
rect 23799 32181 23808 32215
rect 23756 32172 23808 32181
rect 24952 32240 25004 32292
rect 25872 32240 25924 32292
rect 26240 32240 26292 32292
rect 26792 32240 26844 32292
rect 27068 32240 27120 32292
rect 27252 32240 27304 32292
rect 29276 32419 29328 32428
rect 29276 32385 29285 32419
rect 29285 32385 29319 32419
rect 29319 32385 29328 32419
rect 29276 32376 29328 32385
rect 29644 32376 29696 32428
rect 30012 32419 30064 32428
rect 30012 32385 30021 32419
rect 30021 32385 30055 32419
rect 30055 32385 30064 32419
rect 30012 32376 30064 32385
rect 30380 32512 30432 32564
rect 31944 32512 31996 32564
rect 32036 32512 32088 32564
rect 32404 32512 32456 32564
rect 30472 32444 30524 32496
rect 30288 32376 30340 32428
rect 30380 32308 30432 32360
rect 30932 32308 30984 32360
rect 29644 32240 29696 32292
rect 30012 32240 30064 32292
rect 30104 32240 30156 32292
rect 32128 32444 32180 32496
rect 32036 32376 32088 32428
rect 32404 32376 32456 32428
rect 32864 32376 32916 32428
rect 33232 32376 33284 32428
rect 33968 32512 34020 32564
rect 34336 32555 34388 32564
rect 34336 32521 34345 32555
rect 34345 32521 34379 32555
rect 34379 32521 34388 32555
rect 34336 32512 34388 32521
rect 37464 32555 37516 32564
rect 37464 32521 37473 32555
rect 37473 32521 37507 32555
rect 37507 32521 37516 32555
rect 37464 32512 37516 32521
rect 33508 32487 33560 32496
rect 33508 32453 33517 32487
rect 33517 32453 33551 32487
rect 33551 32453 33560 32487
rect 33508 32444 33560 32453
rect 33692 32419 33744 32428
rect 33692 32385 33701 32419
rect 33701 32385 33735 32419
rect 33735 32385 33744 32419
rect 33692 32376 33744 32385
rect 33784 32419 33836 32428
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 37188 32444 37240 32496
rect 35164 32419 35216 32428
rect 35164 32385 35173 32419
rect 35173 32385 35207 32419
rect 35207 32385 35216 32419
rect 35164 32376 35216 32385
rect 35440 32419 35492 32428
rect 35440 32385 35449 32419
rect 35449 32385 35483 32419
rect 35483 32385 35492 32419
rect 35440 32376 35492 32385
rect 34428 32240 34480 32292
rect 36084 32419 36136 32428
rect 36084 32385 36093 32419
rect 36093 32385 36127 32419
rect 36127 32385 36136 32419
rect 36084 32376 36136 32385
rect 36176 32376 36228 32428
rect 39856 32512 39908 32564
rect 40960 32512 41012 32564
rect 42064 32512 42116 32564
rect 43076 32512 43128 32564
rect 43352 32512 43404 32564
rect 37832 32419 37884 32428
rect 37832 32385 37841 32419
rect 37841 32385 37875 32419
rect 37875 32385 37884 32419
rect 37832 32376 37884 32385
rect 38292 32444 38344 32496
rect 39304 32444 39356 32496
rect 39396 32444 39448 32496
rect 25596 32172 25648 32224
rect 28448 32172 28500 32224
rect 28724 32172 28776 32224
rect 30380 32172 30432 32224
rect 32312 32172 32364 32224
rect 32404 32215 32456 32224
rect 32404 32181 32413 32215
rect 32413 32181 32447 32215
rect 32447 32181 32456 32215
rect 32404 32172 32456 32181
rect 32772 32172 32824 32224
rect 33140 32172 33192 32224
rect 33784 32172 33836 32224
rect 34244 32172 34296 32224
rect 36360 32308 36412 32360
rect 36452 32308 36504 32360
rect 37096 32308 37148 32360
rect 39120 32419 39172 32428
rect 39120 32385 39129 32419
rect 39129 32385 39163 32419
rect 39163 32385 39172 32419
rect 39120 32376 39172 32385
rect 41236 32444 41288 32496
rect 40592 32419 40644 32428
rect 40592 32385 40601 32419
rect 40601 32385 40635 32419
rect 40635 32385 40644 32419
rect 40592 32376 40644 32385
rect 40776 32376 40828 32428
rect 41604 32419 41656 32428
rect 41604 32385 41613 32419
rect 41613 32385 41647 32419
rect 41647 32385 41656 32419
rect 41604 32376 41656 32385
rect 43260 32376 43312 32428
rect 40040 32308 40092 32360
rect 35808 32240 35860 32292
rect 39028 32240 39080 32292
rect 39396 32240 39448 32292
rect 39488 32283 39540 32292
rect 39488 32249 39497 32283
rect 39497 32249 39531 32283
rect 39531 32249 39540 32283
rect 39488 32240 39540 32249
rect 35440 32172 35492 32224
rect 40500 32308 40552 32360
rect 42892 32172 42944 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 12624 31968 12676 32020
rect 13268 32011 13320 32020
rect 13268 31977 13277 32011
rect 13277 31977 13311 32011
rect 13311 31977 13320 32011
rect 13268 31968 13320 31977
rect 14280 32011 14332 32020
rect 14280 31977 14289 32011
rect 14289 31977 14323 32011
rect 14323 31977 14332 32011
rect 14280 31968 14332 31977
rect 14556 31968 14608 32020
rect 17040 32011 17092 32020
rect 17040 31977 17049 32011
rect 17049 31977 17083 32011
rect 17083 31977 17092 32011
rect 17040 31968 17092 31977
rect 20720 31968 20772 32020
rect 12716 31900 12768 31952
rect 14096 31900 14148 31952
rect 14188 31832 14240 31884
rect 12624 31807 12676 31816
rect 12624 31773 12633 31807
rect 12633 31773 12667 31807
rect 12667 31773 12676 31807
rect 12624 31764 12676 31773
rect 13360 31764 13412 31816
rect 15384 31943 15436 31952
rect 15384 31909 15393 31943
rect 15393 31909 15427 31943
rect 15427 31909 15436 31943
rect 15384 31900 15436 31909
rect 17224 31900 17276 31952
rect 19064 31900 19116 31952
rect 20628 31900 20680 31952
rect 26976 31968 27028 32020
rect 29828 31968 29880 32020
rect 30288 31968 30340 32020
rect 24768 31900 24820 31952
rect 28816 31900 28868 31952
rect 32312 32011 32364 32020
rect 32312 31977 32321 32011
rect 32321 31977 32355 32011
rect 32355 31977 32364 32011
rect 32312 31968 32364 31977
rect 32772 31968 32824 32020
rect 31944 31900 31996 31952
rect 34244 31968 34296 32020
rect 34612 31968 34664 32020
rect 37096 31968 37148 32020
rect 37648 32011 37700 32020
rect 37648 31977 37657 32011
rect 37657 31977 37691 32011
rect 37691 31977 37700 32011
rect 37648 31968 37700 31977
rect 37832 31968 37884 32020
rect 39212 31968 39264 32020
rect 39856 31968 39908 32020
rect 14464 31807 14516 31816
rect 14464 31773 14473 31807
rect 14473 31773 14507 31807
rect 14507 31773 14516 31807
rect 14464 31764 14516 31773
rect 16304 31832 16356 31884
rect 15200 31807 15252 31816
rect 15200 31773 15209 31807
rect 15209 31773 15243 31807
rect 15243 31773 15252 31807
rect 15200 31764 15252 31773
rect 18052 31807 18104 31816
rect 13452 31739 13504 31748
rect 13452 31705 13461 31739
rect 13461 31705 13495 31739
rect 13495 31705 13504 31739
rect 13452 31696 13504 31705
rect 18052 31773 18061 31807
rect 18061 31773 18095 31807
rect 18095 31773 18104 31807
rect 18052 31764 18104 31773
rect 19984 31875 20036 31884
rect 19984 31841 19993 31875
rect 19993 31841 20027 31875
rect 20027 31841 20036 31875
rect 19984 31832 20036 31841
rect 20352 31832 20404 31884
rect 20904 31832 20956 31884
rect 15936 31628 15988 31680
rect 17868 31696 17920 31748
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 19064 31764 19116 31816
rect 20536 31764 20588 31816
rect 21088 31764 21140 31816
rect 21364 31764 21416 31816
rect 21916 31832 21968 31884
rect 23020 31764 23072 31816
rect 23296 31764 23348 31816
rect 25044 31832 25096 31884
rect 24216 31764 24268 31816
rect 24952 31807 25004 31816
rect 24952 31773 24961 31807
rect 24961 31773 24995 31807
rect 24995 31773 25004 31807
rect 24952 31764 25004 31773
rect 25136 31807 25188 31816
rect 25136 31773 25145 31807
rect 25145 31773 25179 31807
rect 25179 31773 25188 31807
rect 25136 31764 25188 31773
rect 25872 31807 25924 31816
rect 17960 31671 18012 31680
rect 17960 31637 17969 31671
rect 17969 31637 18003 31671
rect 18003 31637 18012 31671
rect 17960 31628 18012 31637
rect 20904 31696 20956 31748
rect 22376 31696 22428 31748
rect 23664 31696 23716 31748
rect 24584 31696 24636 31748
rect 25872 31773 25881 31807
rect 25881 31773 25915 31807
rect 25915 31773 25924 31807
rect 25872 31764 25924 31773
rect 26792 31764 26844 31816
rect 30104 31832 30156 31884
rect 33140 31832 33192 31884
rect 33232 31832 33284 31884
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 18236 31628 18288 31680
rect 19248 31628 19300 31680
rect 19800 31671 19852 31680
rect 19800 31637 19809 31671
rect 19809 31637 19843 31671
rect 19843 31637 19852 31671
rect 19800 31628 19852 31637
rect 20076 31628 20128 31680
rect 22284 31628 22336 31680
rect 22928 31628 22980 31680
rect 24676 31628 24728 31680
rect 24768 31628 24820 31680
rect 25228 31628 25280 31680
rect 25596 31628 25648 31680
rect 26056 31739 26108 31748
rect 26056 31705 26065 31739
rect 26065 31705 26099 31739
rect 26099 31705 26108 31739
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 26056 31696 26108 31705
rect 26240 31628 26292 31680
rect 28540 31696 28592 31748
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 28908 31807 28960 31816
rect 28908 31773 28917 31807
rect 28917 31773 28951 31807
rect 28951 31773 28960 31807
rect 28908 31764 28960 31773
rect 29920 31764 29972 31816
rect 30196 31764 30248 31816
rect 32036 31807 32088 31816
rect 32036 31773 32045 31807
rect 32045 31773 32079 31807
rect 32079 31773 32088 31807
rect 32036 31764 32088 31773
rect 32220 31764 32272 31816
rect 32680 31764 32732 31816
rect 32772 31807 32824 31816
rect 32772 31773 32781 31807
rect 32781 31773 32815 31807
rect 32815 31773 32824 31807
rect 32772 31764 32824 31773
rect 34704 31900 34756 31952
rect 35440 31900 35492 31952
rect 37188 31900 37240 31952
rect 34244 31875 34296 31884
rect 34244 31841 34253 31875
rect 34253 31841 34287 31875
rect 34287 31841 34296 31875
rect 34244 31832 34296 31841
rect 34428 31764 34480 31816
rect 34612 31696 34664 31748
rect 35072 31739 35124 31748
rect 35072 31705 35081 31739
rect 35081 31705 35115 31739
rect 35115 31705 35124 31739
rect 35992 31764 36044 31816
rect 36084 31807 36136 31816
rect 36084 31773 36093 31807
rect 36093 31773 36127 31807
rect 36127 31773 36136 31807
rect 36084 31764 36136 31773
rect 35072 31696 35124 31705
rect 35440 31696 35492 31748
rect 35716 31696 35768 31748
rect 37740 31832 37792 31884
rect 37004 31807 37056 31816
rect 37004 31773 37013 31807
rect 37013 31773 37047 31807
rect 37047 31773 37056 31807
rect 37004 31764 37056 31773
rect 38016 31807 38068 31816
rect 38016 31773 38025 31807
rect 38025 31773 38059 31807
rect 38059 31773 38068 31807
rect 38016 31764 38068 31773
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 40316 31900 40368 31952
rect 40132 31832 40184 31884
rect 40592 31968 40644 32020
rect 41880 31968 41932 32020
rect 40224 31764 40276 31816
rect 41236 31832 41288 31884
rect 42892 31875 42944 31884
rect 42892 31841 42901 31875
rect 42901 31841 42935 31875
rect 42935 31841 42944 31875
rect 42892 31832 42944 31841
rect 43168 31875 43220 31884
rect 43168 31841 43177 31875
rect 43177 31841 43211 31875
rect 43211 31841 43220 31875
rect 43168 31832 43220 31841
rect 39948 31696 40000 31748
rect 40684 31807 40736 31816
rect 40684 31773 40693 31807
rect 40693 31773 40727 31807
rect 40727 31773 40736 31807
rect 40684 31764 40736 31773
rect 42432 31696 42484 31748
rect 29276 31628 29328 31680
rect 32496 31628 32548 31680
rect 33784 31671 33836 31680
rect 33784 31637 33793 31671
rect 33793 31637 33827 31671
rect 33827 31637 33836 31671
rect 33784 31628 33836 31637
rect 39396 31628 39448 31680
rect 40408 31628 40460 31680
rect 41420 31671 41472 31680
rect 41420 31637 41429 31671
rect 41429 31637 41463 31671
rect 41463 31637 41472 31671
rect 41420 31628 41472 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 13268 31356 13320 31408
rect 15384 31424 15436 31476
rect 15660 31467 15712 31476
rect 15660 31433 15669 31467
rect 15669 31433 15703 31467
rect 15703 31433 15712 31467
rect 15660 31424 15712 31433
rect 17960 31424 18012 31476
rect 18512 31424 18564 31476
rect 18880 31424 18932 31476
rect 19156 31424 19208 31476
rect 15016 31356 15068 31408
rect 17224 31399 17276 31408
rect 17224 31365 17233 31399
rect 17233 31365 17267 31399
rect 17267 31365 17276 31399
rect 17224 31356 17276 31365
rect 17776 31356 17828 31408
rect 15936 31288 15988 31340
rect 15844 31263 15896 31272
rect 15844 31229 15853 31263
rect 15853 31229 15887 31263
rect 15887 31229 15896 31263
rect 15844 31220 15896 31229
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 18236 31331 18288 31340
rect 18236 31297 18242 31331
rect 18242 31297 18276 31331
rect 18276 31297 18288 31331
rect 18236 31288 18288 31297
rect 18604 31288 18656 31340
rect 19524 31288 19576 31340
rect 17684 31220 17736 31272
rect 13452 31152 13504 31204
rect 18696 31263 18748 31272
rect 18696 31229 18705 31263
rect 18705 31229 18739 31263
rect 18739 31229 18748 31263
rect 18696 31220 18748 31229
rect 18880 31220 18932 31272
rect 19064 31220 19116 31272
rect 21088 31424 21140 31476
rect 25044 31424 25096 31476
rect 19984 31356 20036 31408
rect 20260 31356 20312 31408
rect 12900 31084 12952 31136
rect 17224 31127 17276 31136
rect 17224 31093 17233 31127
rect 17233 31093 17267 31127
rect 17267 31093 17276 31127
rect 17224 31084 17276 31093
rect 19984 31220 20036 31272
rect 20444 31263 20496 31272
rect 20444 31229 20453 31263
rect 20453 31229 20487 31263
rect 20487 31229 20496 31263
rect 20444 31220 20496 31229
rect 21364 31331 21416 31340
rect 21364 31297 21373 31331
rect 21373 31297 21407 31331
rect 21407 31297 21416 31331
rect 21364 31288 21416 31297
rect 22376 31356 22428 31408
rect 23940 31356 23992 31408
rect 21916 31288 21968 31340
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 24400 31399 24452 31408
rect 24400 31365 24409 31399
rect 24409 31365 24443 31399
rect 24443 31365 24452 31399
rect 24400 31356 24452 31365
rect 24768 31356 24820 31408
rect 26148 31424 26200 31476
rect 25596 31356 25648 31408
rect 26056 31356 26108 31408
rect 28632 31356 28684 31408
rect 20812 31220 20864 31272
rect 21272 31220 21324 31272
rect 21640 31220 21692 31272
rect 22652 31220 22704 31272
rect 23112 31220 23164 31272
rect 23388 31263 23440 31272
rect 23388 31229 23397 31263
rect 23397 31229 23431 31263
rect 23431 31229 23440 31263
rect 23388 31220 23440 31229
rect 23572 31220 23624 31272
rect 20628 31195 20680 31204
rect 20628 31161 20637 31195
rect 20637 31161 20671 31195
rect 20671 31161 20680 31195
rect 20628 31152 20680 31161
rect 22560 31152 22612 31204
rect 24584 31288 24636 31340
rect 24676 31331 24728 31340
rect 24676 31297 24685 31331
rect 24685 31297 24719 31331
rect 24719 31297 24728 31331
rect 24676 31288 24728 31297
rect 25044 31288 25096 31340
rect 26148 31263 26200 31272
rect 26148 31229 26157 31263
rect 26157 31229 26191 31263
rect 26191 31229 26200 31263
rect 26148 31220 26200 31229
rect 28908 31331 28960 31340
rect 28908 31297 28917 31331
rect 28917 31297 28951 31331
rect 28951 31297 28960 31331
rect 28908 31288 28960 31297
rect 29092 31331 29144 31340
rect 29092 31297 29101 31331
rect 29101 31297 29135 31331
rect 29135 31297 29144 31331
rect 29092 31288 29144 31297
rect 37280 31424 37332 31476
rect 29552 31356 29604 31408
rect 30288 31399 30340 31408
rect 30288 31365 30297 31399
rect 30297 31365 30331 31399
rect 30331 31365 30340 31399
rect 30288 31356 30340 31365
rect 29920 31288 29972 31340
rect 30932 31331 30984 31340
rect 30932 31297 30941 31331
rect 30941 31297 30975 31331
rect 30975 31297 30984 31331
rect 30932 31288 30984 31297
rect 32404 31356 32456 31408
rect 33232 31356 33284 31408
rect 33968 31399 34020 31408
rect 33968 31365 33977 31399
rect 33977 31365 34011 31399
rect 34011 31365 34020 31399
rect 33968 31356 34020 31365
rect 35532 31356 35584 31408
rect 35992 31356 36044 31408
rect 31576 31288 31628 31340
rect 31852 31288 31904 31340
rect 32496 31331 32548 31340
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 32864 31331 32916 31340
rect 32864 31297 32873 31331
rect 32873 31297 32907 31331
rect 32907 31297 32916 31331
rect 32864 31288 32916 31297
rect 34704 31288 34756 31340
rect 34980 31288 35032 31340
rect 31760 31220 31812 31272
rect 33692 31220 33744 31272
rect 35716 31263 35768 31272
rect 30380 31152 30432 31204
rect 33600 31152 33652 31204
rect 35716 31229 35725 31263
rect 35725 31229 35759 31263
rect 35759 31229 35768 31263
rect 35716 31220 35768 31229
rect 36452 31220 36504 31272
rect 36636 31331 36688 31340
rect 36636 31297 36645 31331
rect 36645 31297 36679 31331
rect 36679 31297 36688 31331
rect 36636 31288 36688 31297
rect 37004 31356 37056 31408
rect 38752 31399 38804 31408
rect 38752 31365 38761 31399
rect 38761 31365 38795 31399
rect 38795 31365 38804 31399
rect 38752 31356 38804 31365
rect 38292 31288 38344 31340
rect 39120 31288 39172 31340
rect 37372 31220 37424 31272
rect 36084 31152 36136 31204
rect 37280 31152 37332 31204
rect 38384 31220 38436 31272
rect 39396 31331 39448 31340
rect 39396 31297 39405 31331
rect 39405 31297 39439 31331
rect 39439 31297 39448 31331
rect 39396 31288 39448 31297
rect 41880 31467 41932 31476
rect 41880 31433 41889 31467
rect 41889 31433 41923 31467
rect 41923 31433 41932 31467
rect 41880 31424 41932 31433
rect 40040 31356 40092 31408
rect 40316 31356 40368 31408
rect 40500 31288 40552 31340
rect 40960 31288 41012 31340
rect 41328 31331 41380 31340
rect 41328 31297 41337 31331
rect 41337 31297 41371 31331
rect 41371 31297 41380 31331
rect 41328 31288 41380 31297
rect 41420 31288 41472 31340
rect 42892 31288 42944 31340
rect 39580 31220 39632 31272
rect 41696 31220 41748 31272
rect 42708 31220 42760 31272
rect 43996 31220 44048 31272
rect 38108 31152 38160 31204
rect 40040 31152 40092 31204
rect 40132 31152 40184 31204
rect 21640 31084 21692 31136
rect 24032 31084 24084 31136
rect 24952 31084 25004 31136
rect 29736 31084 29788 31136
rect 29920 31127 29972 31136
rect 29920 31093 29929 31127
rect 29929 31093 29963 31127
rect 29963 31093 29972 31127
rect 29920 31084 29972 31093
rect 30012 31084 30064 31136
rect 32312 31127 32364 31136
rect 32312 31093 32321 31127
rect 32321 31093 32355 31127
rect 32355 31093 32364 31127
rect 32312 31084 32364 31093
rect 32772 31127 32824 31136
rect 32772 31093 32781 31127
rect 32781 31093 32815 31127
rect 32815 31093 32824 31127
rect 32772 31084 32824 31093
rect 33324 31127 33376 31136
rect 33324 31093 33333 31127
rect 33333 31093 33367 31127
rect 33367 31093 33376 31127
rect 33324 31084 33376 31093
rect 35716 31084 35768 31136
rect 36268 31084 36320 31136
rect 36728 31127 36780 31136
rect 36728 31093 36737 31127
rect 36737 31093 36771 31127
rect 36771 31093 36780 31127
rect 36728 31084 36780 31093
rect 37648 31084 37700 31136
rect 38384 31127 38436 31136
rect 38384 31093 38393 31127
rect 38393 31093 38427 31127
rect 38427 31093 38436 31127
rect 38384 31084 38436 31093
rect 39212 31084 39264 31136
rect 40224 31127 40276 31136
rect 40224 31093 40233 31127
rect 40233 31093 40267 31127
rect 40267 31093 40276 31127
rect 40224 31084 40276 31093
rect 40868 31084 40920 31136
rect 41972 31084 42024 31136
rect 42800 31084 42852 31136
rect 43260 31084 43312 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 12624 30880 12676 30932
rect 13268 30880 13320 30932
rect 11888 30812 11940 30864
rect 15016 30880 15068 30932
rect 18144 30923 18196 30932
rect 18144 30889 18153 30923
rect 18153 30889 18187 30923
rect 18187 30889 18196 30923
rect 18144 30880 18196 30889
rect 18696 30880 18748 30932
rect 18788 30880 18840 30932
rect 20628 30880 20680 30932
rect 20720 30923 20772 30932
rect 20720 30889 20729 30923
rect 20729 30889 20763 30923
rect 20763 30889 20772 30923
rect 20720 30880 20772 30889
rect 22100 30880 22152 30932
rect 23388 30880 23440 30932
rect 28908 30880 28960 30932
rect 29736 30880 29788 30932
rect 30932 30880 30984 30932
rect 33784 30880 33836 30932
rect 35808 30880 35860 30932
rect 36636 30880 36688 30932
rect 36820 30880 36872 30932
rect 37556 30923 37608 30932
rect 37556 30889 37565 30923
rect 37565 30889 37599 30923
rect 37599 30889 37608 30923
rect 37556 30880 37608 30889
rect 37740 30880 37792 30932
rect 20996 30812 21048 30864
rect 21364 30855 21416 30864
rect 21364 30821 21373 30855
rect 21373 30821 21407 30855
rect 21407 30821 21416 30855
rect 21364 30812 21416 30821
rect 21916 30855 21968 30864
rect 21916 30821 21925 30855
rect 21925 30821 21959 30855
rect 21959 30821 21968 30855
rect 21916 30812 21968 30821
rect 26056 30812 26108 30864
rect 27620 30812 27672 30864
rect 18420 30744 18472 30796
rect 19432 30744 19484 30796
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13452 30676 13504 30728
rect 15844 30676 15896 30728
rect 17776 30608 17828 30660
rect 18880 30719 18932 30728
rect 18880 30685 18889 30719
rect 18889 30685 18923 30719
rect 18923 30685 18932 30719
rect 18880 30676 18932 30685
rect 19340 30676 19392 30728
rect 20444 30744 20496 30796
rect 19708 30719 19760 30728
rect 19708 30685 19717 30719
rect 19717 30685 19751 30719
rect 19751 30685 19760 30719
rect 19708 30676 19760 30685
rect 19892 30719 19944 30728
rect 19892 30685 19901 30719
rect 19901 30685 19935 30719
rect 19935 30685 19944 30719
rect 19892 30676 19944 30685
rect 21088 30676 21140 30728
rect 21180 30676 21232 30728
rect 21640 30676 21692 30728
rect 22376 30719 22428 30728
rect 22376 30685 22385 30719
rect 22385 30685 22419 30719
rect 22419 30685 22428 30719
rect 22376 30676 22428 30685
rect 23112 30676 23164 30728
rect 23756 30676 23808 30728
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 25228 30676 25280 30728
rect 25596 30676 25648 30728
rect 25780 30676 25832 30728
rect 25872 30719 25924 30728
rect 25872 30685 25881 30719
rect 25881 30685 25915 30719
rect 25915 30685 25924 30719
rect 25872 30676 25924 30685
rect 29000 30812 29052 30864
rect 30196 30812 30248 30864
rect 38476 30880 38528 30932
rect 40132 30923 40184 30932
rect 40132 30889 40141 30923
rect 40141 30889 40175 30923
rect 40175 30889 40184 30923
rect 40132 30880 40184 30889
rect 40960 30812 41012 30864
rect 27896 30719 27948 30728
rect 27896 30685 27905 30719
rect 27905 30685 27939 30719
rect 27939 30685 27948 30719
rect 27896 30676 27948 30685
rect 28816 30744 28868 30796
rect 30748 30787 30800 30796
rect 30748 30753 30757 30787
rect 30757 30753 30791 30787
rect 30791 30753 30800 30787
rect 30748 30744 30800 30753
rect 31852 30744 31904 30796
rect 27344 30608 27396 30660
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 29920 30719 29972 30728
rect 29920 30685 29929 30719
rect 29929 30685 29963 30719
rect 29963 30685 29972 30719
rect 29920 30676 29972 30685
rect 30932 30676 30984 30728
rect 32312 30676 32364 30728
rect 32588 30676 32640 30728
rect 34152 30787 34204 30796
rect 34152 30753 34161 30787
rect 34161 30753 34195 30787
rect 34195 30753 34204 30787
rect 34152 30744 34204 30753
rect 36544 30744 36596 30796
rect 32772 30719 32824 30728
rect 32772 30685 32781 30719
rect 32781 30685 32815 30719
rect 32815 30685 32824 30719
rect 32772 30676 32824 30685
rect 33600 30719 33652 30728
rect 33600 30685 33609 30719
rect 33609 30685 33643 30719
rect 33643 30685 33652 30719
rect 33600 30676 33652 30685
rect 34428 30676 34480 30728
rect 34704 30676 34756 30728
rect 35440 30719 35492 30728
rect 35440 30685 35449 30719
rect 35449 30685 35483 30719
rect 35483 30685 35492 30719
rect 35440 30676 35492 30685
rect 35624 30719 35676 30728
rect 35624 30685 35633 30719
rect 35633 30685 35667 30719
rect 35667 30685 35676 30719
rect 35624 30676 35676 30685
rect 36268 30719 36320 30728
rect 36268 30685 36277 30719
rect 36277 30685 36311 30719
rect 36311 30685 36320 30719
rect 36268 30676 36320 30685
rect 30288 30608 30340 30660
rect 32864 30608 32916 30660
rect 37280 30676 37332 30728
rect 38108 30676 38160 30728
rect 36636 30608 36688 30660
rect 39396 30676 39448 30728
rect 41236 30744 41288 30796
rect 42708 30744 42760 30796
rect 42800 30787 42852 30796
rect 42800 30753 42809 30787
rect 42809 30753 42843 30787
rect 42843 30753 42852 30787
rect 42800 30744 42852 30753
rect 39856 30676 39908 30728
rect 40224 30719 40276 30728
rect 40224 30685 40233 30719
rect 40233 30685 40267 30719
rect 40267 30685 40276 30719
rect 40224 30676 40276 30685
rect 40684 30719 40736 30728
rect 40684 30685 40693 30719
rect 40693 30685 40727 30719
rect 40727 30685 40736 30719
rect 40684 30676 40736 30685
rect 40868 30719 40920 30728
rect 40868 30685 40877 30719
rect 40877 30685 40911 30719
rect 40911 30685 40920 30719
rect 40868 30676 40920 30685
rect 41972 30719 42024 30728
rect 41972 30685 41981 30719
rect 41981 30685 42015 30719
rect 42015 30685 42024 30719
rect 41972 30676 42024 30685
rect 11980 30540 12032 30592
rect 13912 30540 13964 30592
rect 15660 30540 15712 30592
rect 15936 30583 15988 30592
rect 15936 30549 15945 30583
rect 15945 30549 15979 30583
rect 15979 30549 15988 30583
rect 15936 30540 15988 30549
rect 16948 30540 17000 30592
rect 19156 30540 19208 30592
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 19708 30540 19760 30592
rect 20076 30540 20128 30592
rect 20536 30540 20588 30592
rect 23112 30540 23164 30592
rect 25136 30540 25188 30592
rect 27252 30583 27304 30592
rect 27252 30549 27261 30583
rect 27261 30549 27295 30583
rect 27295 30549 27304 30583
rect 27252 30540 27304 30549
rect 28908 30540 28960 30592
rect 29184 30540 29236 30592
rect 29920 30540 29972 30592
rect 30656 30540 30708 30592
rect 31944 30583 31996 30592
rect 31944 30549 31953 30583
rect 31953 30549 31987 30583
rect 31987 30549 31996 30583
rect 31944 30540 31996 30549
rect 37372 30540 37424 30592
rect 38568 30540 38620 30592
rect 38844 30540 38896 30592
rect 41328 30540 41380 30592
rect 41696 30583 41748 30592
rect 41696 30549 41705 30583
rect 41705 30549 41739 30583
rect 41739 30549 41748 30583
rect 41696 30540 41748 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17960 30336 18012 30388
rect 12900 30268 12952 30320
rect 12992 30200 13044 30252
rect 16488 30268 16540 30320
rect 18052 30268 18104 30320
rect 18788 30268 18840 30320
rect 19984 30336 20036 30388
rect 20628 30336 20680 30388
rect 27252 30336 27304 30388
rect 27344 30336 27396 30388
rect 31852 30336 31904 30388
rect 32404 30336 32456 30388
rect 35624 30336 35676 30388
rect 16120 30243 16172 30252
rect 16120 30209 16129 30243
rect 16129 30209 16163 30243
rect 16163 30209 16172 30243
rect 16120 30200 16172 30209
rect 16764 30200 16816 30252
rect 19340 30311 19392 30320
rect 19340 30277 19349 30311
rect 19349 30277 19383 30311
rect 19383 30277 19392 30311
rect 19340 30268 19392 30277
rect 21088 30311 21140 30320
rect 21088 30277 21097 30311
rect 21097 30277 21131 30311
rect 21131 30277 21140 30311
rect 21088 30268 21140 30277
rect 13820 30175 13872 30184
rect 13820 30141 13829 30175
rect 13829 30141 13863 30175
rect 13863 30141 13872 30175
rect 13820 30132 13872 30141
rect 14096 30175 14148 30184
rect 14096 30141 14105 30175
rect 14105 30141 14139 30175
rect 14139 30141 14148 30175
rect 14096 30132 14148 30141
rect 18420 30132 18472 30184
rect 19524 30243 19576 30252
rect 19524 30209 19569 30243
rect 19569 30209 19576 30243
rect 19524 30200 19576 30209
rect 13084 30107 13136 30116
rect 13084 30073 13093 30107
rect 13093 30073 13127 30107
rect 13127 30073 13136 30107
rect 13084 30064 13136 30073
rect 16304 30107 16356 30116
rect 16304 30073 16313 30107
rect 16313 30073 16347 30107
rect 16347 30073 16356 30107
rect 16304 30064 16356 30073
rect 17500 30064 17552 30116
rect 19248 30064 19300 30116
rect 19984 30200 20036 30252
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 22008 30243 22060 30252
rect 22008 30209 22017 30243
rect 22017 30209 22051 30243
rect 22051 30209 22060 30243
rect 22008 30200 22060 30209
rect 22468 30268 22520 30320
rect 25780 30268 25832 30320
rect 26700 30268 26752 30320
rect 20260 30132 20312 30184
rect 21180 30132 21232 30184
rect 23388 30132 23440 30184
rect 21272 30064 21324 30116
rect 25044 30064 25096 30116
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25596 30200 25648 30252
rect 25872 30243 25924 30252
rect 25872 30209 25881 30243
rect 25881 30209 25915 30243
rect 25915 30209 25924 30243
rect 25872 30200 25924 30209
rect 27804 30268 27856 30320
rect 29092 30268 29144 30320
rect 29368 30268 29420 30320
rect 29920 30268 29972 30320
rect 30748 30268 30800 30320
rect 31208 30268 31260 30320
rect 32036 30268 32088 30320
rect 27620 30200 27672 30252
rect 28448 30200 28500 30252
rect 27344 30175 27396 30184
rect 27344 30141 27353 30175
rect 27353 30141 27387 30175
rect 27387 30141 27396 30175
rect 27344 30132 27396 30141
rect 28816 30243 28868 30252
rect 28816 30209 28825 30243
rect 28825 30209 28859 30243
rect 28859 30209 28868 30243
rect 28816 30200 28868 30209
rect 30012 30200 30064 30252
rect 30656 30200 30708 30252
rect 37004 30268 37056 30320
rect 29644 30132 29696 30184
rect 31208 30175 31260 30184
rect 31208 30141 31217 30175
rect 31217 30141 31251 30175
rect 31251 30141 31260 30175
rect 31208 30132 31260 30141
rect 32956 30200 33008 30252
rect 33968 30200 34020 30252
rect 34152 30200 34204 30252
rect 34520 30243 34572 30252
rect 34520 30209 34529 30243
rect 34529 30209 34563 30243
rect 34563 30209 34572 30243
rect 34520 30200 34572 30209
rect 35348 30200 35400 30252
rect 31944 30132 31996 30184
rect 13544 29996 13596 30048
rect 17868 30039 17920 30048
rect 17868 30005 17877 30039
rect 17877 30005 17911 30039
rect 17911 30005 17920 30039
rect 17868 29996 17920 30005
rect 18144 29996 18196 30048
rect 20168 29996 20220 30048
rect 20444 29996 20496 30048
rect 21180 29996 21232 30048
rect 22652 30039 22704 30048
rect 22652 30005 22661 30039
rect 22661 30005 22695 30039
rect 22695 30005 22704 30039
rect 22652 29996 22704 30005
rect 24308 29996 24360 30048
rect 24676 29996 24728 30048
rect 26148 29996 26200 30048
rect 26792 29996 26844 30048
rect 27712 30039 27764 30048
rect 27712 30005 27721 30039
rect 27721 30005 27755 30039
rect 27755 30005 27764 30039
rect 27712 29996 27764 30005
rect 29828 29996 29880 30048
rect 33692 30132 33744 30184
rect 35716 30243 35768 30252
rect 35716 30209 35725 30243
rect 35725 30209 35759 30243
rect 35759 30209 35768 30243
rect 35716 30200 35768 30209
rect 35808 30243 35860 30252
rect 35808 30209 35817 30243
rect 35817 30209 35851 30243
rect 35851 30209 35860 30243
rect 35808 30200 35860 30209
rect 36452 30132 36504 30184
rect 33968 30064 34020 30116
rect 37280 30200 37332 30252
rect 38200 30336 38252 30388
rect 40040 30336 40092 30388
rect 40868 30336 40920 30388
rect 41144 30336 41196 30388
rect 41328 30336 41380 30388
rect 41696 30336 41748 30388
rect 37924 30268 37976 30320
rect 38108 30268 38160 30320
rect 40592 30268 40644 30320
rect 41420 30268 41472 30320
rect 37740 30243 37792 30252
rect 37740 30209 37749 30243
rect 37749 30209 37783 30243
rect 37783 30209 37792 30243
rect 37740 30200 37792 30209
rect 37832 30243 37884 30252
rect 37832 30209 37850 30243
rect 37850 30209 37884 30243
rect 37832 30200 37884 30209
rect 38200 30200 38252 30252
rect 38752 30132 38804 30184
rect 39580 30200 39632 30252
rect 40132 30200 40184 30252
rect 43260 30200 43312 30252
rect 39580 30064 39632 30116
rect 40500 30064 40552 30116
rect 42064 30064 42116 30116
rect 32772 29996 32824 30048
rect 38384 29996 38436 30048
rect 39028 30039 39080 30048
rect 39028 30005 39037 30039
rect 39037 30005 39071 30039
rect 39071 30005 39080 30039
rect 39028 29996 39080 30005
rect 39672 29996 39724 30048
rect 42800 30039 42852 30048
rect 42800 30005 42809 30039
rect 42809 30005 42843 30039
rect 42843 30005 42852 30039
rect 42800 29996 42852 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 11980 29835 12032 29844
rect 11980 29801 11989 29835
rect 11989 29801 12023 29835
rect 12023 29801 12032 29835
rect 11980 29792 12032 29801
rect 12992 29792 13044 29844
rect 14096 29792 14148 29844
rect 13636 29724 13688 29776
rect 16120 29656 16172 29708
rect 18604 29792 18656 29844
rect 18696 29792 18748 29844
rect 20352 29792 20404 29844
rect 20996 29792 21048 29844
rect 16856 29724 16908 29776
rect 21916 29835 21968 29844
rect 21916 29801 21925 29835
rect 21925 29801 21959 29835
rect 21959 29801 21968 29835
rect 21916 29792 21968 29801
rect 22376 29835 22428 29844
rect 22376 29801 22385 29835
rect 22385 29801 22419 29835
rect 22419 29801 22428 29835
rect 22376 29792 22428 29801
rect 26056 29792 26108 29844
rect 27620 29792 27672 29844
rect 27712 29792 27764 29844
rect 35992 29792 36044 29844
rect 36912 29792 36964 29844
rect 37004 29835 37056 29844
rect 37004 29801 37013 29835
rect 37013 29801 37047 29835
rect 37047 29801 37056 29835
rect 37004 29792 37056 29801
rect 39212 29835 39264 29844
rect 39212 29801 39221 29835
rect 39221 29801 39255 29835
rect 39255 29801 39264 29835
rect 39212 29792 39264 29801
rect 39580 29792 39632 29844
rect 41328 29792 41380 29844
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 12808 29631 12860 29640
rect 12808 29597 12817 29631
rect 12817 29597 12851 29631
rect 12851 29597 12860 29631
rect 12808 29588 12860 29597
rect 12992 29631 13044 29640
rect 12992 29597 13001 29631
rect 13001 29597 13035 29631
rect 13035 29597 13044 29631
rect 12992 29588 13044 29597
rect 13176 29588 13228 29640
rect 13544 29631 13596 29640
rect 13544 29597 13553 29631
rect 13553 29597 13587 29631
rect 13587 29597 13596 29631
rect 13544 29588 13596 29597
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 15936 29588 15988 29640
rect 16304 29588 16356 29640
rect 16120 29520 16172 29572
rect 17500 29588 17552 29640
rect 17868 29631 17920 29640
rect 17868 29597 17877 29631
rect 17877 29597 17911 29631
rect 17911 29597 17920 29631
rect 17868 29588 17920 29597
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 18880 29631 18932 29640
rect 18880 29597 18889 29631
rect 18889 29597 18923 29631
rect 18923 29597 18932 29631
rect 18880 29588 18932 29597
rect 18972 29588 19024 29640
rect 20076 29631 20128 29640
rect 20076 29597 20085 29631
rect 20085 29597 20119 29631
rect 20119 29597 20128 29631
rect 20076 29588 20128 29597
rect 20168 29631 20220 29640
rect 20168 29597 20177 29631
rect 20177 29597 20211 29631
rect 20211 29597 20220 29631
rect 20168 29588 20220 29597
rect 20352 29631 20404 29640
rect 20352 29597 20361 29631
rect 20361 29597 20395 29631
rect 20395 29597 20404 29631
rect 20352 29588 20404 29597
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 24032 29724 24084 29776
rect 27804 29724 27856 29776
rect 31024 29724 31076 29776
rect 33232 29724 33284 29776
rect 34060 29724 34112 29776
rect 35348 29724 35400 29776
rect 37832 29724 37884 29776
rect 38568 29724 38620 29776
rect 23296 29699 23348 29708
rect 23296 29665 23305 29699
rect 23305 29665 23339 29699
rect 23339 29665 23348 29699
rect 23296 29656 23348 29665
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 22560 29588 22612 29640
rect 22652 29588 22704 29640
rect 12992 29452 13044 29504
rect 15844 29452 15896 29504
rect 16396 29495 16448 29504
rect 16396 29461 16405 29495
rect 16405 29461 16439 29495
rect 16439 29461 16448 29495
rect 16396 29452 16448 29461
rect 17316 29495 17368 29504
rect 17316 29461 17325 29495
rect 17325 29461 17359 29495
rect 17359 29461 17368 29495
rect 17316 29452 17368 29461
rect 17960 29495 18012 29504
rect 19340 29520 19392 29572
rect 20996 29520 21048 29572
rect 23480 29588 23532 29640
rect 24952 29656 25004 29708
rect 24584 29588 24636 29640
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25872 29588 25924 29640
rect 26792 29588 26844 29640
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 29828 29588 29880 29640
rect 33232 29588 33284 29640
rect 33416 29588 33468 29640
rect 33876 29588 33928 29640
rect 37004 29656 37056 29708
rect 38108 29656 38160 29708
rect 40316 29699 40368 29708
rect 40316 29665 40325 29699
rect 40325 29665 40359 29699
rect 40359 29665 40368 29699
rect 40316 29656 40368 29665
rect 40408 29699 40460 29708
rect 40408 29665 40417 29699
rect 40417 29665 40451 29699
rect 40451 29665 40460 29699
rect 40408 29656 40460 29665
rect 40592 29724 40644 29776
rect 42248 29724 42300 29776
rect 42892 29767 42944 29776
rect 42892 29733 42901 29767
rect 42901 29733 42935 29767
rect 42935 29733 42944 29767
rect 42892 29724 42944 29733
rect 41144 29656 41196 29708
rect 41420 29656 41472 29708
rect 34060 29588 34112 29640
rect 34244 29588 34296 29640
rect 34520 29588 34572 29640
rect 36176 29588 36228 29640
rect 37096 29588 37148 29640
rect 37280 29631 37332 29640
rect 37280 29597 37289 29631
rect 37289 29597 37323 29631
rect 37323 29597 37332 29631
rect 37280 29588 37332 29597
rect 37924 29588 37976 29640
rect 38568 29588 38620 29640
rect 24216 29520 24268 29572
rect 25228 29520 25280 29572
rect 28632 29520 28684 29572
rect 31208 29520 31260 29572
rect 17960 29461 17975 29495
rect 17975 29461 18009 29495
rect 18009 29461 18012 29495
rect 17960 29452 18012 29461
rect 19156 29452 19208 29504
rect 22008 29452 22060 29504
rect 23480 29452 23532 29504
rect 24584 29495 24636 29504
rect 24584 29461 24593 29495
rect 24593 29461 24627 29495
rect 24627 29461 24636 29495
rect 24584 29452 24636 29461
rect 28540 29495 28592 29504
rect 28540 29461 28549 29495
rect 28549 29461 28583 29495
rect 28583 29461 28592 29495
rect 28540 29452 28592 29461
rect 31116 29452 31168 29504
rect 34428 29520 34480 29572
rect 36728 29520 36780 29572
rect 37004 29563 37056 29572
rect 37004 29529 37013 29563
rect 37013 29529 37047 29563
rect 37047 29529 37056 29563
rect 37004 29520 37056 29529
rect 39948 29588 40000 29640
rect 31944 29495 31996 29504
rect 31944 29461 31953 29495
rect 31953 29461 31987 29495
rect 31987 29461 31996 29495
rect 31944 29452 31996 29461
rect 34060 29452 34112 29504
rect 34520 29452 34572 29504
rect 35164 29452 35216 29504
rect 39028 29520 39080 29572
rect 41512 29631 41564 29640
rect 41512 29597 41521 29631
rect 41521 29597 41555 29631
rect 41555 29597 41564 29631
rect 41512 29588 41564 29597
rect 41328 29520 41380 29572
rect 42248 29563 42300 29572
rect 42248 29529 42257 29563
rect 42257 29529 42291 29563
rect 42291 29529 42300 29563
rect 42248 29520 42300 29529
rect 42616 29520 42668 29572
rect 42892 29520 42944 29572
rect 43260 29563 43312 29572
rect 43260 29529 43269 29563
rect 43269 29529 43303 29563
rect 43303 29529 43312 29563
rect 43260 29520 43312 29529
rect 37188 29452 37240 29504
rect 39304 29452 39356 29504
rect 39580 29452 39632 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 12808 29248 12860 29300
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 12900 29112 12952 29121
rect 14280 29248 14332 29300
rect 16396 29248 16448 29300
rect 13912 29223 13964 29232
rect 13912 29189 13921 29223
rect 13921 29189 13955 29223
rect 13955 29189 13964 29223
rect 13912 29180 13964 29189
rect 15200 29180 15252 29232
rect 13636 29112 13688 29164
rect 14832 29155 14884 29164
rect 14832 29121 14841 29155
rect 14841 29121 14875 29155
rect 14875 29121 14884 29155
rect 14832 29112 14884 29121
rect 15292 29112 15344 29164
rect 15844 29155 15896 29164
rect 15844 29121 15853 29155
rect 15853 29121 15887 29155
rect 15887 29121 15896 29155
rect 15844 29112 15896 29121
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 16212 29155 16264 29164
rect 16212 29121 16221 29155
rect 16221 29121 16255 29155
rect 16255 29121 16264 29155
rect 16212 29112 16264 29121
rect 16856 29112 16908 29164
rect 18052 29248 18104 29300
rect 18144 29248 18196 29300
rect 17868 29180 17920 29232
rect 18972 29248 19024 29300
rect 20076 29291 20128 29300
rect 20076 29257 20085 29291
rect 20085 29257 20119 29291
rect 20119 29257 20128 29291
rect 20076 29248 20128 29257
rect 20536 29291 20588 29300
rect 18604 29180 18656 29232
rect 19984 29180 20036 29232
rect 12992 28976 13044 29028
rect 13176 28976 13228 29028
rect 16764 29044 16816 29096
rect 16948 29044 17000 29096
rect 18972 29155 19024 29164
rect 18972 29121 18981 29155
rect 18981 29121 19015 29155
rect 19015 29121 19024 29155
rect 18972 29112 19024 29121
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 20536 29257 20545 29291
rect 20545 29257 20579 29291
rect 20579 29257 20588 29291
rect 20536 29248 20588 29257
rect 21456 29291 21508 29300
rect 21456 29257 21465 29291
rect 21465 29257 21499 29291
rect 21499 29257 21508 29291
rect 21456 29248 21508 29257
rect 22192 29248 22244 29300
rect 23480 29248 23532 29300
rect 25136 29291 25188 29300
rect 25136 29257 25145 29291
rect 25145 29257 25179 29291
rect 25179 29257 25188 29291
rect 25136 29248 25188 29257
rect 20352 29180 20404 29232
rect 18144 29044 18196 29096
rect 19340 29044 19392 29096
rect 20260 29044 20312 29096
rect 20536 29112 20588 29164
rect 22744 29180 22796 29232
rect 24860 29180 24912 29232
rect 28356 29248 28408 29300
rect 29644 29248 29696 29300
rect 30012 29291 30064 29300
rect 30012 29257 30021 29291
rect 30021 29257 30055 29291
rect 30055 29257 30064 29291
rect 30012 29248 30064 29257
rect 29460 29180 29512 29232
rect 30656 29180 30708 29232
rect 20628 29087 20680 29096
rect 20628 29053 20637 29087
rect 20637 29053 20671 29087
rect 20671 29053 20680 29087
rect 20628 29044 20680 29053
rect 23020 29155 23072 29164
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 23848 29044 23900 29096
rect 24400 29155 24452 29164
rect 24400 29121 24409 29155
rect 24409 29121 24443 29155
rect 24443 29121 24452 29155
rect 24400 29112 24452 29121
rect 25044 29155 25096 29164
rect 25044 29121 25053 29155
rect 25053 29121 25087 29155
rect 25087 29121 25096 29155
rect 25044 29112 25096 29121
rect 25320 29112 25372 29164
rect 26424 29155 26476 29164
rect 26424 29121 26433 29155
rect 26433 29121 26467 29155
rect 26467 29121 26476 29155
rect 26424 29112 26476 29121
rect 24768 29044 24820 29096
rect 25596 29087 25648 29096
rect 25596 29053 25605 29087
rect 25605 29053 25639 29087
rect 25639 29053 25648 29087
rect 29000 29112 29052 29164
rect 25596 29044 25648 29053
rect 26792 29044 26844 29096
rect 21916 28976 21968 29028
rect 22560 28976 22612 29028
rect 23388 28976 23440 29028
rect 30288 29112 30340 29164
rect 30932 29112 30984 29164
rect 31116 29248 31168 29300
rect 31208 29291 31260 29300
rect 31208 29257 31217 29291
rect 31217 29257 31251 29291
rect 31251 29257 31260 29291
rect 31208 29248 31260 29257
rect 32220 29248 32272 29300
rect 34704 29248 34756 29300
rect 35164 29248 35216 29300
rect 37004 29248 37056 29300
rect 37372 29248 37424 29300
rect 37924 29248 37976 29300
rect 32496 29155 32548 29164
rect 32496 29121 32505 29155
rect 32505 29121 32539 29155
rect 32539 29121 32548 29155
rect 32496 29112 32548 29121
rect 32680 29155 32732 29164
rect 32680 29121 32689 29155
rect 32689 29121 32723 29155
rect 32723 29121 32732 29155
rect 32680 29112 32732 29121
rect 33416 29112 33468 29164
rect 33600 29112 33652 29164
rect 34520 29180 34572 29232
rect 34428 29112 34480 29164
rect 34888 29180 34940 29232
rect 35348 29180 35400 29232
rect 34704 29112 34756 29164
rect 38200 29180 38252 29232
rect 38476 29223 38528 29232
rect 38476 29189 38485 29223
rect 38485 29189 38519 29223
rect 38519 29189 38528 29223
rect 38476 29180 38528 29189
rect 41052 29248 41104 29300
rect 41144 29248 41196 29300
rect 38108 29112 38160 29164
rect 38568 29112 38620 29164
rect 39580 29180 39632 29232
rect 40316 29180 40368 29232
rect 40776 29180 40828 29232
rect 31668 29044 31720 29096
rect 31760 29087 31812 29096
rect 31760 29053 31769 29087
rect 31769 29053 31803 29087
rect 31803 29053 31812 29087
rect 31760 29044 31812 29053
rect 31944 29044 31996 29096
rect 37740 29044 37792 29096
rect 29828 28976 29880 29028
rect 33508 29019 33560 29028
rect 33508 28985 33517 29019
rect 33517 28985 33551 29019
rect 33551 28985 33560 29019
rect 33508 28976 33560 28985
rect 33876 28976 33928 29028
rect 13084 28951 13136 28960
rect 13084 28917 13093 28951
rect 13093 28917 13127 28951
rect 13127 28917 13136 28951
rect 13084 28908 13136 28917
rect 13452 28908 13504 28960
rect 18420 28951 18472 28960
rect 18420 28917 18429 28951
rect 18429 28917 18463 28951
rect 18463 28917 18472 28951
rect 18420 28908 18472 28917
rect 25872 28908 25924 28960
rect 29184 28908 29236 28960
rect 29276 28908 29328 28960
rect 31576 28908 31628 28960
rect 34152 28908 34204 28960
rect 34888 28976 34940 29028
rect 35624 28976 35676 29028
rect 35900 28976 35952 29028
rect 38936 29044 38988 29096
rect 39028 29087 39080 29096
rect 39028 29053 39037 29087
rect 39037 29053 39071 29087
rect 39071 29053 39080 29087
rect 39028 29044 39080 29053
rect 39488 29155 39540 29164
rect 39488 29121 39497 29155
rect 39497 29121 39531 29155
rect 39531 29121 39540 29155
rect 39488 29112 39540 29121
rect 39672 29155 39724 29164
rect 39672 29121 39681 29155
rect 39681 29121 39715 29155
rect 39715 29121 39724 29155
rect 39672 29112 39724 29121
rect 40408 29112 40460 29164
rect 41052 29112 41104 29164
rect 41420 29112 41472 29164
rect 39580 29044 39632 29096
rect 40960 29087 41012 29096
rect 40960 29053 40969 29087
rect 40969 29053 41003 29087
rect 41003 29053 41012 29087
rect 40960 29044 41012 29053
rect 38476 28976 38528 29028
rect 40592 28976 40644 29028
rect 35532 28951 35584 28960
rect 35532 28917 35541 28951
rect 35541 28917 35575 28951
rect 35575 28917 35584 28951
rect 35532 28908 35584 28917
rect 37280 28908 37332 28960
rect 40500 28908 40552 28960
rect 41052 28908 41104 28960
rect 41512 29044 41564 29096
rect 42248 29112 42300 29164
rect 41880 28908 41932 28960
rect 41972 28908 42024 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 14832 28704 14884 28756
rect 16120 28747 16172 28756
rect 16120 28713 16129 28747
rect 16129 28713 16163 28747
rect 16163 28713 16172 28747
rect 16120 28704 16172 28713
rect 16764 28747 16816 28756
rect 16764 28713 16773 28747
rect 16773 28713 16807 28747
rect 16807 28713 16816 28747
rect 16764 28704 16816 28713
rect 13360 28636 13412 28688
rect 16028 28636 16080 28688
rect 18420 28679 18472 28688
rect 16212 28611 16264 28620
rect 16212 28577 16221 28611
rect 16221 28577 16255 28611
rect 16255 28577 16264 28611
rect 16212 28568 16264 28577
rect 17316 28568 17368 28620
rect 18420 28645 18429 28679
rect 18429 28645 18463 28679
rect 18463 28645 18472 28679
rect 18420 28636 18472 28645
rect 19340 28704 19392 28756
rect 20168 28704 20220 28756
rect 20720 28636 20772 28688
rect 17960 28568 18012 28620
rect 20904 28611 20956 28620
rect 13452 28543 13504 28552
rect 13452 28509 13461 28543
rect 13461 28509 13495 28543
rect 13495 28509 13504 28543
rect 13452 28500 13504 28509
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 15844 28500 15896 28552
rect 16948 28500 17000 28552
rect 18052 28500 18104 28552
rect 18512 28500 18564 28552
rect 20904 28577 20913 28611
rect 20913 28577 20947 28611
rect 20947 28577 20956 28611
rect 20904 28568 20956 28577
rect 25872 28636 25924 28688
rect 19984 28500 20036 28552
rect 20536 28543 20588 28552
rect 20536 28509 20545 28543
rect 20545 28509 20579 28543
rect 20579 28509 20588 28543
rect 20536 28500 20588 28509
rect 22192 28500 22244 28552
rect 23388 28568 23440 28620
rect 26332 28568 26384 28620
rect 23572 28500 23624 28552
rect 28356 28704 28408 28756
rect 30288 28704 30340 28756
rect 31392 28704 31444 28756
rect 33784 28704 33836 28756
rect 34060 28704 34112 28756
rect 35348 28747 35400 28756
rect 35348 28713 35357 28747
rect 35357 28713 35391 28747
rect 35391 28713 35400 28747
rect 35348 28704 35400 28713
rect 35900 28747 35952 28756
rect 35900 28713 35909 28747
rect 35909 28713 35943 28747
rect 35943 28713 35952 28747
rect 35900 28704 35952 28713
rect 37004 28704 37056 28756
rect 37556 28704 37608 28756
rect 38752 28704 38804 28756
rect 26516 28636 26568 28688
rect 26700 28611 26752 28620
rect 26700 28577 26709 28611
rect 26709 28577 26743 28611
rect 26743 28577 26752 28611
rect 26700 28568 26752 28577
rect 27712 28636 27764 28688
rect 31484 28636 31536 28688
rect 31576 28636 31628 28688
rect 30748 28611 30800 28620
rect 30748 28577 30757 28611
rect 30757 28577 30791 28611
rect 30791 28577 30800 28611
rect 30748 28568 30800 28577
rect 30840 28568 30892 28620
rect 26976 28543 27028 28552
rect 26976 28509 26985 28543
rect 26985 28509 27019 28543
rect 27019 28509 27028 28543
rect 26976 28500 27028 28509
rect 27068 28543 27120 28552
rect 27068 28509 27102 28543
rect 27102 28509 27120 28543
rect 27068 28500 27120 28509
rect 31024 28500 31076 28552
rect 14740 28432 14792 28484
rect 20352 28432 20404 28484
rect 13912 28364 13964 28416
rect 15108 28364 15160 28416
rect 15200 28364 15252 28416
rect 18236 28364 18288 28416
rect 25964 28432 26016 28484
rect 24032 28407 24084 28416
rect 24032 28373 24041 28407
rect 24041 28373 24075 28407
rect 24075 28373 24084 28407
rect 24032 28364 24084 28373
rect 25044 28407 25096 28416
rect 25044 28373 25053 28407
rect 25053 28373 25087 28407
rect 25087 28373 25096 28407
rect 25044 28364 25096 28373
rect 25688 28364 25740 28416
rect 26976 28364 27028 28416
rect 27068 28364 27120 28416
rect 28080 28432 28132 28484
rect 30104 28432 30156 28484
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 28356 28407 28408 28416
rect 28356 28373 28365 28407
rect 28365 28373 28399 28407
rect 28399 28373 28408 28407
rect 28356 28364 28408 28373
rect 28632 28364 28684 28416
rect 28816 28407 28868 28416
rect 28816 28373 28825 28407
rect 28825 28373 28859 28407
rect 28859 28373 28868 28407
rect 28816 28364 28868 28373
rect 30564 28407 30616 28416
rect 30564 28373 30573 28407
rect 30573 28373 30607 28407
rect 30607 28373 30616 28407
rect 30564 28364 30616 28373
rect 31208 28364 31260 28416
rect 31576 28432 31628 28484
rect 34704 28568 34756 28620
rect 32956 28500 33008 28552
rect 33876 28543 33928 28552
rect 33876 28509 33885 28543
rect 33885 28509 33919 28543
rect 33919 28509 33928 28543
rect 33876 28500 33928 28509
rect 33968 28543 34020 28552
rect 33968 28509 33977 28543
rect 33977 28509 34011 28543
rect 34011 28509 34020 28543
rect 33968 28500 34020 28509
rect 34060 28500 34112 28552
rect 34612 28500 34664 28552
rect 35808 28543 35860 28552
rect 35808 28509 35817 28543
rect 35817 28509 35851 28543
rect 35851 28509 35860 28543
rect 35808 28500 35860 28509
rect 35900 28500 35952 28552
rect 37832 28636 37884 28688
rect 38016 28568 38068 28620
rect 38292 28636 38344 28688
rect 41052 28636 41104 28688
rect 41328 28636 41380 28688
rect 42984 28636 43036 28688
rect 41420 28611 41472 28620
rect 41420 28577 41429 28611
rect 41429 28577 41463 28611
rect 41463 28577 41472 28611
rect 41420 28568 41472 28577
rect 42800 28611 42852 28620
rect 42800 28577 42809 28611
rect 42809 28577 42843 28611
rect 42843 28577 42852 28611
rect 42800 28568 42852 28577
rect 43260 28568 43312 28620
rect 36176 28500 36228 28552
rect 34428 28432 34480 28484
rect 35348 28432 35400 28484
rect 36544 28364 36596 28416
rect 36912 28407 36964 28416
rect 36912 28373 36921 28407
rect 36921 28373 36955 28407
rect 36955 28373 36964 28407
rect 36912 28364 36964 28373
rect 38476 28500 38528 28552
rect 40040 28500 40092 28552
rect 40224 28500 40276 28552
rect 38016 28475 38068 28484
rect 38016 28441 38025 28475
rect 38025 28441 38059 28475
rect 38059 28441 38068 28475
rect 38016 28432 38068 28441
rect 38200 28432 38252 28484
rect 38568 28432 38620 28484
rect 39120 28432 39172 28484
rect 39672 28432 39724 28484
rect 41696 28432 41748 28484
rect 41880 28543 41932 28552
rect 41880 28509 41889 28543
rect 41889 28509 41923 28543
rect 41923 28509 41932 28543
rect 41880 28500 41932 28509
rect 41972 28543 42024 28552
rect 41972 28509 41981 28543
rect 41981 28509 42015 28543
rect 42015 28509 42024 28543
rect 41972 28500 42024 28509
rect 42892 28543 42944 28552
rect 42892 28509 42901 28543
rect 42901 28509 42935 28543
rect 42935 28509 42944 28543
rect 42892 28500 42944 28509
rect 40684 28364 40736 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 14740 28160 14792 28212
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 21456 28160 21508 28212
rect 22100 28160 22152 28212
rect 23020 28160 23072 28212
rect 25688 28160 25740 28212
rect 26424 28160 26476 28212
rect 28356 28160 28408 28212
rect 30840 28160 30892 28212
rect 32772 28160 32824 28212
rect 32956 28203 33008 28212
rect 32956 28169 32965 28203
rect 32965 28169 32999 28203
rect 32999 28169 33008 28203
rect 32956 28160 33008 28169
rect 33232 28160 33284 28212
rect 34428 28160 34480 28212
rect 35440 28160 35492 28212
rect 35900 28203 35952 28212
rect 35900 28169 35909 28203
rect 35909 28169 35943 28203
rect 35943 28169 35952 28203
rect 35900 28160 35952 28169
rect 36360 28203 36412 28212
rect 36360 28169 36369 28203
rect 36369 28169 36403 28203
rect 36403 28169 36412 28203
rect 36360 28160 36412 28169
rect 40868 28160 40920 28212
rect 41788 28160 41840 28212
rect 13176 28024 13228 28076
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 17316 28024 17368 28076
rect 18052 28092 18104 28144
rect 18236 28067 18288 28076
rect 18236 28033 18245 28067
rect 18245 28033 18279 28067
rect 18279 28033 18288 28067
rect 18236 28024 18288 28033
rect 20904 28135 20956 28144
rect 20904 28101 20913 28135
rect 20913 28101 20947 28135
rect 20947 28101 20956 28135
rect 20904 28092 20956 28101
rect 21364 28135 21416 28144
rect 21364 28101 21373 28135
rect 21373 28101 21407 28135
rect 21407 28101 21416 28135
rect 21364 28092 21416 28101
rect 24032 28092 24084 28144
rect 12992 27956 13044 28008
rect 15108 27999 15160 28008
rect 15108 27965 15117 27999
rect 15117 27965 15151 27999
rect 15151 27965 15160 27999
rect 15108 27956 15160 27965
rect 20628 27956 20680 28008
rect 19984 27888 20036 27940
rect 13912 27820 13964 27872
rect 14556 27820 14608 27872
rect 22928 27863 22980 27872
rect 22928 27829 22937 27863
rect 22937 27829 22971 27863
rect 22971 27829 22980 27863
rect 22928 27820 22980 27829
rect 23940 28024 23992 28076
rect 26792 28092 26844 28144
rect 28264 28092 28316 28144
rect 25504 28024 25556 28076
rect 28724 28024 28776 28076
rect 29368 28067 29420 28076
rect 29368 28033 29377 28067
rect 29377 28033 29411 28067
rect 29411 28033 29420 28067
rect 29368 28024 29420 28033
rect 29552 28067 29604 28076
rect 29552 28033 29561 28067
rect 29561 28033 29595 28067
rect 29595 28033 29604 28067
rect 29552 28024 29604 28033
rect 32496 28092 32548 28144
rect 37096 28092 37148 28144
rect 38108 28092 38160 28144
rect 23756 27999 23808 28008
rect 23756 27965 23765 27999
rect 23765 27965 23799 27999
rect 23799 27965 23808 27999
rect 23756 27956 23808 27965
rect 27344 27956 27396 28008
rect 27896 27956 27948 28008
rect 31208 28067 31260 28076
rect 31208 28033 31217 28067
rect 31217 28033 31251 28067
rect 31251 28033 31260 28067
rect 31208 28024 31260 28033
rect 31392 28024 31444 28076
rect 34520 28067 34572 28076
rect 34520 28033 34529 28067
rect 34529 28033 34563 28067
rect 34563 28033 34572 28067
rect 34520 28024 34572 28033
rect 32588 27956 32640 28008
rect 32772 27999 32824 28008
rect 32772 27965 32806 27999
rect 32806 27965 32824 27999
rect 32772 27956 32824 27965
rect 34244 27956 34296 28008
rect 34336 27999 34388 28008
rect 34336 27965 34345 27999
rect 34345 27965 34379 27999
rect 34379 27965 34388 27999
rect 34336 27956 34388 27965
rect 34428 27999 34480 28008
rect 34428 27965 34437 27999
rect 34437 27965 34471 27999
rect 34471 27965 34480 27999
rect 34428 27956 34480 27965
rect 35164 28024 35216 28076
rect 36452 28024 36504 28076
rect 38016 28067 38068 28076
rect 38016 28033 38030 28067
rect 38030 28033 38064 28067
rect 38064 28033 38068 28067
rect 38016 28024 38068 28033
rect 42800 28092 42852 28144
rect 40040 28024 40092 28076
rect 40592 28024 40644 28076
rect 41236 28024 41288 28076
rect 43444 28024 43496 28076
rect 43996 28024 44048 28076
rect 35992 27956 36044 28008
rect 37004 27956 37056 28008
rect 39856 27956 39908 28008
rect 40408 27956 40460 28008
rect 41052 27999 41104 28008
rect 41052 27965 41061 27999
rect 41061 27965 41095 27999
rect 41095 27965 41104 27999
rect 41052 27956 41104 27965
rect 29920 27888 29972 27940
rect 25872 27820 25924 27872
rect 29000 27820 29052 27872
rect 29644 27820 29696 27872
rect 30288 27820 30340 27872
rect 32128 27888 32180 27940
rect 32312 27888 32364 27940
rect 37464 27931 37516 27940
rect 37464 27897 37473 27931
rect 37473 27897 37507 27931
rect 37507 27897 37516 27931
rect 37464 27888 37516 27897
rect 38568 27888 38620 27940
rect 31392 27863 31444 27872
rect 31392 27829 31401 27863
rect 31401 27829 31435 27863
rect 31435 27829 31444 27863
rect 31392 27820 31444 27829
rect 33784 27820 33836 27872
rect 36912 27820 36964 27872
rect 37832 27820 37884 27872
rect 38200 27820 38252 27872
rect 38660 27820 38712 27872
rect 39948 27888 40000 27940
rect 41972 27956 42024 28008
rect 39212 27820 39264 27872
rect 39396 27820 39448 27872
rect 43076 27820 43128 27872
rect 43536 27820 43588 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 20260 27591 20312 27600
rect 20260 27557 20269 27591
rect 20269 27557 20303 27591
rect 20303 27557 20312 27591
rect 20260 27548 20312 27557
rect 20444 27548 20496 27600
rect 23664 27548 23716 27600
rect 26056 27616 26108 27668
rect 27344 27659 27396 27668
rect 27344 27625 27353 27659
rect 27353 27625 27387 27659
rect 27387 27625 27396 27659
rect 27344 27616 27396 27625
rect 23848 27591 23900 27600
rect 23848 27557 23857 27591
rect 23857 27557 23891 27591
rect 23891 27557 23900 27591
rect 23848 27548 23900 27557
rect 25504 27591 25556 27600
rect 25504 27557 25513 27591
rect 25513 27557 25547 27591
rect 25547 27557 25556 27591
rect 25504 27548 25556 27557
rect 13820 27480 13872 27532
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 18972 27412 19024 27464
rect 19432 27344 19484 27396
rect 21456 27412 21508 27464
rect 23756 27455 23808 27464
rect 23756 27421 23765 27455
rect 23765 27421 23799 27455
rect 23799 27421 23808 27455
rect 24400 27480 24452 27532
rect 25044 27480 25096 27532
rect 26700 27548 26752 27600
rect 27988 27616 28040 27668
rect 29368 27616 29420 27668
rect 29552 27616 29604 27668
rect 27804 27548 27856 27600
rect 32772 27616 32824 27668
rect 34428 27616 34480 27668
rect 34980 27616 35032 27668
rect 35348 27616 35400 27668
rect 35532 27616 35584 27668
rect 36360 27616 36412 27668
rect 36636 27616 36688 27668
rect 38108 27616 38160 27668
rect 38844 27616 38896 27668
rect 40408 27616 40460 27668
rect 40500 27616 40552 27668
rect 41420 27659 41472 27668
rect 41420 27625 41429 27659
rect 41429 27625 41463 27659
rect 41463 27625 41472 27659
rect 41420 27616 41472 27625
rect 23756 27412 23808 27421
rect 23940 27455 23992 27464
rect 23940 27421 23949 27455
rect 23949 27421 23983 27455
rect 23983 27421 23992 27455
rect 23940 27412 23992 27421
rect 24768 27412 24820 27464
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 31392 27523 31444 27532
rect 31392 27489 31401 27523
rect 31401 27489 31435 27523
rect 31435 27489 31444 27523
rect 31392 27480 31444 27489
rect 31668 27548 31720 27600
rect 32680 27548 32732 27600
rect 34612 27548 34664 27600
rect 31944 27480 31996 27532
rect 24952 27387 25004 27396
rect 24952 27353 24961 27387
rect 24961 27353 24995 27387
rect 24995 27353 25004 27387
rect 24952 27344 25004 27353
rect 20628 27276 20680 27328
rect 22652 27276 22704 27328
rect 22836 27276 22888 27328
rect 24492 27276 24544 27328
rect 27528 27455 27580 27464
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 27620 27412 27672 27464
rect 27896 27412 27948 27464
rect 28080 27412 28132 27464
rect 29184 27455 29236 27464
rect 29184 27421 29193 27455
rect 29193 27421 29227 27455
rect 29227 27421 29236 27455
rect 29184 27412 29236 27421
rect 30288 27412 30340 27464
rect 33140 27480 33192 27532
rect 34244 27480 34296 27532
rect 32312 27455 32364 27464
rect 32312 27421 32321 27455
rect 32321 27421 32355 27455
rect 32355 27421 32364 27455
rect 32312 27412 32364 27421
rect 32772 27412 32824 27464
rect 33416 27455 33468 27464
rect 33416 27421 33425 27455
rect 33425 27421 33459 27455
rect 33459 27421 33468 27455
rect 33416 27412 33468 27421
rect 34060 27412 34112 27464
rect 34336 27455 34388 27464
rect 34336 27421 34345 27455
rect 34345 27421 34379 27455
rect 34379 27421 34388 27455
rect 34336 27412 34388 27421
rect 35716 27480 35768 27532
rect 35072 27412 35124 27464
rect 35624 27455 35676 27464
rect 35624 27421 35639 27455
rect 35639 27421 35673 27455
rect 35673 27421 35676 27455
rect 35624 27412 35676 27421
rect 36360 27523 36412 27532
rect 36360 27489 36369 27523
rect 36369 27489 36403 27523
rect 36403 27489 36412 27523
rect 36360 27480 36412 27489
rect 36544 27455 36596 27464
rect 26056 27344 26108 27396
rect 28816 27344 28868 27396
rect 30196 27344 30248 27396
rect 32036 27344 32088 27396
rect 32128 27344 32180 27396
rect 33600 27344 33652 27396
rect 27252 27276 27304 27328
rect 27344 27276 27396 27328
rect 28632 27276 28684 27328
rect 30380 27276 30432 27328
rect 32220 27319 32272 27328
rect 32220 27285 32229 27319
rect 32229 27285 32263 27319
rect 32263 27285 32272 27319
rect 32220 27276 32272 27285
rect 35532 27344 35584 27396
rect 36544 27421 36553 27455
rect 36553 27421 36587 27455
rect 36587 27421 36596 27455
rect 36544 27412 36596 27421
rect 37096 27548 37148 27600
rect 37740 27548 37792 27600
rect 39948 27548 40000 27600
rect 41144 27548 41196 27600
rect 42064 27548 42116 27600
rect 38384 27523 38436 27532
rect 38384 27489 38393 27523
rect 38393 27489 38427 27523
rect 38427 27489 38436 27523
rect 38384 27480 38436 27489
rect 37004 27412 37056 27464
rect 38016 27412 38068 27464
rect 38108 27412 38160 27464
rect 38568 27455 38620 27464
rect 38568 27421 38577 27455
rect 38577 27421 38611 27455
rect 38611 27421 38620 27455
rect 38568 27412 38620 27421
rect 39028 27344 39080 27396
rect 39488 27455 39540 27464
rect 39488 27421 39497 27455
rect 39497 27421 39531 27455
rect 39531 27421 39540 27455
rect 39488 27412 39540 27421
rect 41236 27480 41288 27532
rect 40868 27412 40920 27464
rect 41052 27412 41104 27464
rect 41512 27412 41564 27464
rect 42616 27412 42668 27464
rect 34980 27276 35032 27328
rect 35164 27276 35216 27328
rect 36360 27319 36412 27328
rect 36360 27285 36369 27319
rect 36369 27285 36403 27319
rect 36403 27285 36412 27319
rect 36360 27276 36412 27285
rect 36452 27276 36504 27328
rect 38476 27276 38528 27328
rect 40224 27344 40276 27396
rect 41788 27344 41840 27396
rect 40500 27276 40552 27328
rect 41328 27276 41380 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 18144 27072 18196 27124
rect 20720 27072 20772 27124
rect 24952 27072 25004 27124
rect 25688 27115 25740 27124
rect 25688 27081 25697 27115
rect 25697 27081 25731 27115
rect 25731 27081 25740 27115
rect 25688 27072 25740 27081
rect 25780 27072 25832 27124
rect 29184 27115 29236 27124
rect 29184 27081 29193 27115
rect 29193 27081 29227 27115
rect 29227 27081 29236 27115
rect 29184 27072 29236 27081
rect 30380 27115 30432 27124
rect 30380 27081 30389 27115
rect 30389 27081 30423 27115
rect 30423 27081 30432 27115
rect 30380 27072 30432 27081
rect 30840 27072 30892 27124
rect 32220 27072 32272 27124
rect 35808 27072 35860 27124
rect 36176 27115 36228 27124
rect 36176 27081 36185 27115
rect 36185 27081 36219 27115
rect 36219 27081 36228 27115
rect 36176 27072 36228 27081
rect 36544 27072 36596 27124
rect 40684 27072 40736 27124
rect 42616 27115 42668 27124
rect 42616 27081 42625 27115
rect 42625 27081 42659 27115
rect 42659 27081 42668 27115
rect 42616 27072 42668 27081
rect 17224 27004 17276 27056
rect 20444 27047 20496 27056
rect 20444 27013 20453 27047
rect 20453 27013 20487 27047
rect 20487 27013 20496 27047
rect 20444 27004 20496 27013
rect 22836 27004 22888 27056
rect 22928 27004 22980 27056
rect 14280 26868 14332 26920
rect 20628 26936 20680 26988
rect 14832 26868 14884 26920
rect 20260 26868 20312 26920
rect 18512 26732 18564 26784
rect 19800 26775 19852 26784
rect 19800 26741 19809 26775
rect 19809 26741 19843 26775
rect 19843 26741 19852 26775
rect 19800 26732 19852 26741
rect 23388 26936 23440 26988
rect 23664 26979 23716 26988
rect 23664 26945 23673 26979
rect 23673 26945 23707 26979
rect 23707 26945 23716 26979
rect 23664 26936 23716 26945
rect 24768 26936 24820 26988
rect 26332 26936 26384 26988
rect 27252 26936 27304 26988
rect 22376 26911 22428 26920
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 25044 26911 25096 26920
rect 25044 26877 25053 26911
rect 25053 26877 25087 26911
rect 25087 26877 25096 26911
rect 25044 26868 25096 26877
rect 26148 26911 26200 26920
rect 26148 26877 26157 26911
rect 26157 26877 26191 26911
rect 26191 26877 26200 26911
rect 26148 26868 26200 26877
rect 26240 26911 26292 26920
rect 26240 26877 26249 26911
rect 26249 26877 26283 26911
rect 26283 26877 26292 26911
rect 26240 26868 26292 26877
rect 28172 26979 28224 26988
rect 28172 26945 28181 26979
rect 28181 26945 28215 26979
rect 28215 26945 28224 26979
rect 28172 26936 28224 26945
rect 28540 27004 28592 27056
rect 29828 27004 29880 27056
rect 31392 27047 31444 27056
rect 31392 27013 31401 27047
rect 31401 27013 31435 27047
rect 31435 27013 31444 27047
rect 31392 27004 31444 27013
rect 31944 27004 31996 27056
rect 28448 26979 28500 26988
rect 28448 26945 28457 26979
rect 28457 26945 28491 26979
rect 28491 26945 28500 26979
rect 28448 26936 28500 26945
rect 29368 26979 29420 26988
rect 29368 26945 29377 26979
rect 29377 26945 29411 26979
rect 29411 26945 29420 26979
rect 29368 26936 29420 26945
rect 29460 26979 29512 26988
rect 29460 26945 29469 26979
rect 29469 26945 29503 26979
rect 29503 26945 29512 26979
rect 29460 26936 29512 26945
rect 29552 26979 29604 26988
rect 29552 26945 29561 26979
rect 29561 26945 29595 26979
rect 29595 26945 29604 26979
rect 29552 26936 29604 26945
rect 31668 26936 31720 26988
rect 32680 27004 32732 27056
rect 33968 27004 34020 27056
rect 34704 27004 34756 27056
rect 37096 27004 37148 27056
rect 29828 26911 29880 26920
rect 29828 26877 29837 26911
rect 29837 26877 29871 26911
rect 29871 26877 29880 26911
rect 29828 26868 29880 26877
rect 33508 26936 33560 26988
rect 34244 26979 34296 26988
rect 34244 26945 34253 26979
rect 34253 26945 34287 26979
rect 34287 26945 34296 26979
rect 34244 26936 34296 26945
rect 34796 26936 34848 26988
rect 35164 26979 35216 26988
rect 35164 26945 35173 26979
rect 35173 26945 35207 26979
rect 35207 26945 35216 26979
rect 35164 26936 35216 26945
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 32404 26800 32456 26852
rect 33048 26800 33100 26852
rect 22744 26732 22796 26784
rect 23480 26775 23532 26784
rect 23480 26741 23489 26775
rect 23489 26741 23523 26775
rect 23523 26741 23532 26775
rect 23480 26732 23532 26741
rect 24492 26732 24544 26784
rect 27068 26732 27120 26784
rect 27804 26732 27856 26784
rect 33140 26775 33192 26784
rect 33140 26741 33149 26775
rect 33149 26741 33183 26775
rect 33183 26741 33192 26775
rect 33140 26732 33192 26741
rect 33876 26843 33928 26852
rect 33876 26809 33885 26843
rect 33885 26809 33919 26843
rect 33919 26809 33928 26843
rect 33876 26800 33928 26809
rect 34336 26868 34388 26920
rect 36176 26868 36228 26920
rect 37740 26979 37792 26988
rect 37740 26945 37749 26979
rect 37749 26945 37783 26979
rect 37783 26945 37792 26979
rect 37740 26936 37792 26945
rect 37924 26979 37976 26988
rect 37924 26945 37933 26979
rect 37933 26945 37967 26979
rect 37967 26945 37976 26979
rect 37924 26936 37976 26945
rect 38384 27004 38436 27056
rect 39396 27047 39448 27056
rect 39396 27013 39405 27047
rect 39405 27013 39439 27047
rect 39439 27013 39448 27047
rect 39396 27004 39448 27013
rect 39856 27004 39908 27056
rect 38292 26936 38344 26988
rect 40040 26936 40092 26988
rect 40224 26936 40276 26988
rect 40960 26936 41012 26988
rect 36636 26868 36688 26920
rect 34428 26800 34480 26852
rect 35808 26800 35860 26852
rect 37004 26800 37056 26852
rect 37740 26800 37792 26852
rect 38476 26868 38528 26920
rect 38752 26868 38804 26920
rect 39212 26868 39264 26920
rect 40316 26868 40368 26920
rect 40868 26868 40920 26920
rect 39120 26800 39172 26852
rect 39580 26800 39632 26852
rect 43352 27004 43404 27056
rect 41512 26936 41564 26988
rect 41420 26868 41472 26920
rect 43076 26979 43128 26988
rect 43076 26945 43085 26979
rect 43085 26945 43119 26979
rect 43119 26945 43128 26979
rect 43076 26936 43128 26945
rect 34060 26775 34112 26784
rect 34060 26741 34069 26775
rect 34069 26741 34103 26775
rect 34103 26741 34112 26775
rect 34060 26732 34112 26741
rect 34704 26732 34756 26784
rect 36452 26732 36504 26784
rect 37280 26732 37332 26784
rect 38108 26732 38160 26784
rect 38844 26775 38896 26784
rect 38844 26741 38853 26775
rect 38853 26741 38887 26775
rect 38887 26741 38896 26775
rect 38844 26732 38896 26741
rect 40224 26732 40276 26784
rect 41236 26732 41288 26784
rect 42432 26732 42484 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 22836 26528 22888 26580
rect 23572 26528 23624 26580
rect 25872 26528 25924 26580
rect 26148 26528 26200 26580
rect 29552 26528 29604 26580
rect 30564 26571 30616 26580
rect 30564 26537 30573 26571
rect 30573 26537 30607 26571
rect 30607 26537 30616 26571
rect 30564 26528 30616 26537
rect 31484 26528 31536 26580
rect 34520 26528 34572 26580
rect 37096 26528 37148 26580
rect 20352 26460 20404 26512
rect 20628 26460 20680 26512
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 15292 26324 15344 26376
rect 19800 26435 19852 26444
rect 19800 26401 19809 26435
rect 19809 26401 19843 26435
rect 19843 26401 19852 26435
rect 19800 26392 19852 26401
rect 23388 26392 23440 26444
rect 13268 26188 13320 26240
rect 14372 26256 14424 26308
rect 17776 26256 17828 26308
rect 19340 26324 19392 26376
rect 22468 26367 22520 26376
rect 22468 26333 22477 26367
rect 22477 26333 22511 26367
rect 22511 26333 22520 26367
rect 22468 26324 22520 26333
rect 22744 26324 22796 26376
rect 26056 26460 26108 26512
rect 26332 26460 26384 26512
rect 24860 26392 24912 26444
rect 25964 26435 26016 26444
rect 25964 26401 25973 26435
rect 25973 26401 26007 26435
rect 26007 26401 26016 26435
rect 25964 26392 26016 26401
rect 27344 26435 27396 26444
rect 27344 26401 27353 26435
rect 27353 26401 27387 26435
rect 27387 26401 27396 26435
rect 27344 26392 27396 26401
rect 27988 26392 28040 26444
rect 28448 26435 28500 26444
rect 28448 26401 28457 26435
rect 28457 26401 28491 26435
rect 28491 26401 28500 26435
rect 28448 26392 28500 26401
rect 29092 26392 29144 26444
rect 21272 26256 21324 26308
rect 22376 26256 22428 26308
rect 25228 26324 25280 26376
rect 25596 26324 25648 26376
rect 26148 26324 26200 26376
rect 27068 26367 27120 26376
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 29276 26324 29328 26376
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 30932 26392 30984 26444
rect 33140 26392 33192 26444
rect 33876 26460 33928 26512
rect 25780 26299 25832 26308
rect 25780 26265 25789 26299
rect 25789 26265 25823 26299
rect 25823 26265 25832 26299
rect 25780 26256 25832 26265
rect 25872 26256 25924 26308
rect 29092 26256 29144 26308
rect 29184 26299 29236 26308
rect 29184 26265 29193 26299
rect 29193 26265 29227 26299
rect 29227 26265 29236 26299
rect 29184 26256 29236 26265
rect 30656 26256 30708 26308
rect 32680 26256 32732 26308
rect 33784 26367 33836 26376
rect 33784 26333 33793 26367
rect 33793 26333 33827 26367
rect 33827 26333 33836 26367
rect 33784 26324 33836 26333
rect 18604 26188 18656 26240
rect 21456 26231 21508 26240
rect 21456 26197 21465 26231
rect 21465 26197 21499 26231
rect 21499 26197 21508 26231
rect 21456 26188 21508 26197
rect 24584 26188 24636 26240
rect 25688 26188 25740 26240
rect 26056 26188 26108 26240
rect 29000 26188 29052 26240
rect 31024 26231 31076 26240
rect 31024 26197 31033 26231
rect 31033 26197 31067 26231
rect 31067 26197 31076 26231
rect 31024 26188 31076 26197
rect 32312 26188 32364 26240
rect 33232 26256 33284 26308
rect 33508 26256 33560 26308
rect 34060 26324 34112 26376
rect 34612 26324 34664 26376
rect 35716 26392 35768 26444
rect 37004 26392 37056 26444
rect 36176 26324 36228 26376
rect 36636 26367 36688 26376
rect 36636 26333 36645 26367
rect 36645 26333 36679 26367
rect 36679 26333 36688 26367
rect 36636 26324 36688 26333
rect 34520 26188 34572 26240
rect 35256 26299 35308 26308
rect 35256 26265 35265 26299
rect 35265 26265 35299 26299
rect 35299 26265 35308 26299
rect 35256 26256 35308 26265
rect 37464 26256 37516 26308
rect 38384 26460 38436 26512
rect 39120 26392 39172 26444
rect 38384 26324 38436 26376
rect 38568 26324 38620 26376
rect 39396 26435 39448 26444
rect 39396 26401 39405 26435
rect 39405 26401 39439 26435
rect 39439 26401 39448 26435
rect 39396 26392 39448 26401
rect 40040 26435 40092 26444
rect 40040 26401 40049 26435
rect 40049 26401 40083 26435
rect 40083 26401 40092 26435
rect 40040 26392 40092 26401
rect 39672 26324 39724 26376
rect 39948 26324 40000 26376
rect 40408 26367 40460 26376
rect 40408 26333 40417 26367
rect 40417 26333 40451 26367
rect 40451 26333 40460 26367
rect 40408 26324 40460 26333
rect 40500 26367 40552 26376
rect 40500 26333 40509 26367
rect 40509 26333 40543 26367
rect 40543 26333 40552 26367
rect 41052 26392 41104 26444
rect 41880 26392 41932 26444
rect 40500 26324 40552 26333
rect 40684 26367 40736 26376
rect 40684 26333 40693 26367
rect 40693 26333 40727 26367
rect 40727 26333 40736 26367
rect 40684 26324 40736 26333
rect 40960 26324 41012 26376
rect 41788 26367 41840 26376
rect 41788 26333 41797 26367
rect 41797 26333 41831 26367
rect 41831 26333 41840 26367
rect 41788 26324 41840 26333
rect 43076 26392 43128 26444
rect 41972 26256 42024 26308
rect 35808 26188 35860 26240
rect 35900 26188 35952 26240
rect 37924 26188 37976 26240
rect 38752 26231 38804 26240
rect 38752 26197 38761 26231
rect 38761 26197 38795 26231
rect 38795 26197 38804 26231
rect 38752 26188 38804 26197
rect 41236 26188 41288 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 20536 26027 20588 26036
rect 20536 25993 20545 26027
rect 20545 25993 20579 26027
rect 20579 25993 20588 26027
rect 20536 25984 20588 25993
rect 20444 25959 20496 25968
rect 20444 25925 20453 25959
rect 20453 25925 20487 25959
rect 20487 25925 20496 25959
rect 20444 25916 20496 25925
rect 14280 25848 14332 25900
rect 15844 25891 15896 25900
rect 15844 25857 15853 25891
rect 15853 25857 15887 25891
rect 15887 25857 15896 25891
rect 15844 25848 15896 25857
rect 18512 25891 18564 25900
rect 18512 25857 18521 25891
rect 18521 25857 18555 25891
rect 18555 25857 18564 25891
rect 18512 25848 18564 25857
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 22468 25984 22520 26036
rect 25136 25984 25188 26036
rect 25872 25984 25924 26036
rect 26056 25984 26108 26036
rect 26240 25984 26292 26036
rect 28540 25984 28592 26036
rect 25228 25916 25280 25968
rect 27160 25916 27212 25968
rect 30012 25916 30064 25968
rect 31024 26027 31076 26036
rect 31024 25993 31033 26027
rect 31033 25993 31067 26027
rect 31067 25993 31076 26027
rect 31024 25984 31076 25993
rect 31300 25984 31352 26036
rect 31944 25984 31996 26036
rect 32312 25984 32364 26036
rect 32496 25984 32548 26036
rect 33232 25984 33284 26036
rect 33692 25984 33744 26036
rect 34060 26027 34112 26036
rect 34060 25993 34069 26027
rect 34069 25993 34103 26027
rect 34103 25993 34112 26027
rect 34060 25984 34112 25993
rect 22836 25848 22888 25900
rect 23480 25848 23532 25900
rect 23664 25848 23716 25900
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 27252 25848 27304 25900
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 13268 25780 13320 25832
rect 18604 25823 18656 25832
rect 18604 25789 18613 25823
rect 18613 25789 18647 25823
rect 18647 25789 18656 25823
rect 18604 25780 18656 25789
rect 19340 25780 19392 25832
rect 20996 25780 21048 25832
rect 23388 25823 23440 25832
rect 23388 25789 23397 25823
rect 23397 25789 23431 25823
rect 23431 25789 23440 25823
rect 23388 25780 23440 25789
rect 26056 25823 26108 25832
rect 26056 25789 26065 25823
rect 26065 25789 26099 25823
rect 26099 25789 26108 25823
rect 26056 25780 26108 25789
rect 27988 25848 28040 25900
rect 28172 25780 28224 25832
rect 28448 25780 28500 25832
rect 33048 25916 33100 25968
rect 34704 25916 34756 25968
rect 31760 25848 31812 25900
rect 32404 25891 32456 25900
rect 32404 25857 32413 25891
rect 32413 25857 32447 25891
rect 32447 25857 32456 25891
rect 32404 25848 32456 25857
rect 31484 25823 31536 25832
rect 31484 25789 31493 25823
rect 31493 25789 31527 25823
rect 31527 25789 31536 25823
rect 31484 25780 31536 25789
rect 33140 25891 33192 25900
rect 33140 25857 33149 25891
rect 33149 25857 33183 25891
rect 33183 25857 33192 25891
rect 33140 25848 33192 25857
rect 38108 25984 38160 26036
rect 39212 25984 39264 26036
rect 39396 25984 39448 26036
rect 40040 25984 40092 26036
rect 40316 26027 40368 26036
rect 40316 25993 40325 26027
rect 40325 25993 40359 26027
rect 40359 25993 40368 26027
rect 40316 25984 40368 25993
rect 41236 25984 41288 26036
rect 35992 25916 36044 25968
rect 36452 25916 36504 25968
rect 39488 25916 39540 25968
rect 41052 25959 41104 25968
rect 41052 25925 41061 25959
rect 41061 25925 41095 25959
rect 41095 25925 41104 25959
rect 41052 25916 41104 25925
rect 41696 25959 41748 25968
rect 41696 25925 41705 25959
rect 41705 25925 41739 25959
rect 41739 25925 41748 25959
rect 41696 25916 41748 25925
rect 37372 25848 37424 25900
rect 37832 25848 37884 25900
rect 38292 25848 38344 25900
rect 39120 25891 39172 25900
rect 39120 25857 39129 25891
rect 39129 25857 39163 25891
rect 39163 25857 39172 25891
rect 39120 25848 39172 25857
rect 39212 25891 39264 25900
rect 39212 25857 39221 25891
rect 39221 25857 39255 25891
rect 39255 25857 39264 25891
rect 39212 25848 39264 25857
rect 40500 25891 40552 25900
rect 40500 25857 40509 25891
rect 40509 25857 40543 25891
rect 40543 25857 40552 25891
rect 40500 25848 40552 25857
rect 27252 25712 27304 25764
rect 14832 25687 14884 25696
rect 14832 25653 14841 25687
rect 14841 25653 14875 25687
rect 14875 25653 14884 25687
rect 14832 25644 14884 25653
rect 15568 25644 15620 25696
rect 16028 25644 16080 25696
rect 21364 25644 21416 25696
rect 22376 25687 22428 25696
rect 22376 25653 22385 25687
rect 22385 25653 22419 25687
rect 22419 25653 22428 25687
rect 22376 25644 22428 25653
rect 23020 25644 23072 25696
rect 23756 25687 23808 25696
rect 23756 25653 23765 25687
rect 23765 25653 23799 25687
rect 23799 25653 23808 25687
rect 23756 25644 23808 25653
rect 26976 25644 27028 25696
rect 27712 25644 27764 25696
rect 31392 25712 31444 25764
rect 34152 25712 34204 25764
rect 34612 25755 34664 25764
rect 34612 25721 34621 25755
rect 34621 25721 34655 25755
rect 34655 25721 34664 25755
rect 34612 25712 34664 25721
rect 35808 25823 35860 25832
rect 35808 25789 35817 25823
rect 35817 25789 35851 25823
rect 35851 25789 35860 25823
rect 35808 25780 35860 25789
rect 37556 25780 37608 25832
rect 41512 25780 41564 25832
rect 37832 25712 37884 25764
rect 33416 25644 33468 25696
rect 35348 25644 35400 25696
rect 36360 25644 36412 25696
rect 37740 25687 37792 25696
rect 37740 25653 37749 25687
rect 37749 25653 37783 25687
rect 37783 25653 37792 25687
rect 37740 25644 37792 25653
rect 39488 25644 39540 25696
rect 41696 25644 41748 25696
rect 42524 25848 42576 25900
rect 42800 25712 42852 25764
rect 42984 25644 43036 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 14280 25483 14332 25492
rect 14280 25449 14289 25483
rect 14289 25449 14323 25483
rect 14323 25449 14332 25483
rect 14280 25440 14332 25449
rect 19432 25440 19484 25492
rect 23020 25440 23072 25492
rect 23480 25440 23532 25492
rect 23848 25440 23900 25492
rect 24952 25440 25004 25492
rect 25228 25483 25280 25492
rect 25228 25449 25237 25483
rect 25237 25449 25271 25483
rect 25271 25449 25280 25483
rect 25228 25440 25280 25449
rect 27344 25440 27396 25492
rect 27988 25440 28040 25492
rect 29092 25440 29144 25492
rect 18144 25372 18196 25424
rect 20904 25372 20956 25424
rect 15292 25347 15344 25356
rect 15292 25313 15301 25347
rect 15301 25313 15335 25347
rect 15335 25313 15344 25347
rect 15292 25304 15344 25313
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 15568 25279 15620 25288
rect 15568 25245 15602 25279
rect 15602 25245 15620 25279
rect 15568 25236 15620 25245
rect 17684 25279 17736 25288
rect 17684 25245 17693 25279
rect 17693 25245 17727 25279
rect 17727 25245 17736 25279
rect 17684 25236 17736 25245
rect 20812 25236 20864 25288
rect 21456 25236 21508 25288
rect 26056 25372 26108 25424
rect 29184 25372 29236 25424
rect 30288 25440 30340 25492
rect 30748 25440 30800 25492
rect 31484 25440 31536 25492
rect 32404 25440 32456 25492
rect 32772 25440 32824 25492
rect 34060 25440 34112 25492
rect 37372 25440 37424 25492
rect 39120 25440 39172 25492
rect 42616 25440 42668 25492
rect 23756 25304 23808 25356
rect 24768 25304 24820 25356
rect 24952 25347 25004 25356
rect 24952 25313 24961 25347
rect 24961 25313 24995 25347
rect 24995 25313 25004 25347
rect 24952 25304 25004 25313
rect 25964 25304 26016 25356
rect 29460 25304 29512 25356
rect 32680 25372 32732 25424
rect 35532 25372 35584 25424
rect 35900 25372 35952 25424
rect 19432 25168 19484 25220
rect 23480 25236 23532 25288
rect 23848 25279 23900 25288
rect 23848 25245 23857 25279
rect 23857 25245 23891 25279
rect 23891 25245 23900 25279
rect 23848 25236 23900 25245
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 22744 25211 22796 25220
rect 22744 25177 22753 25211
rect 22753 25177 22787 25211
rect 22787 25177 22796 25211
rect 22744 25168 22796 25177
rect 17040 25100 17092 25152
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 17500 25100 17552 25109
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 22836 25100 22888 25152
rect 23112 25168 23164 25220
rect 23940 25168 23992 25220
rect 25136 25236 25188 25288
rect 27620 25236 27672 25288
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 28172 25279 28224 25288
rect 28172 25245 28181 25279
rect 28181 25245 28215 25279
rect 28215 25245 28224 25279
rect 28172 25236 28224 25245
rect 28632 25279 28684 25288
rect 28632 25245 28641 25279
rect 28641 25245 28675 25279
rect 28675 25245 28684 25279
rect 28632 25236 28684 25245
rect 29552 25236 29604 25288
rect 30380 25304 30432 25356
rect 31300 25304 31352 25356
rect 34520 25304 34572 25356
rect 35072 25304 35124 25356
rect 36820 25304 36872 25356
rect 30840 25236 30892 25288
rect 31392 25279 31444 25288
rect 31392 25245 31401 25279
rect 31401 25245 31435 25279
rect 31435 25245 31444 25279
rect 31392 25236 31444 25245
rect 32312 25236 32364 25288
rect 32404 25279 32456 25288
rect 32404 25245 32413 25279
rect 32413 25245 32447 25279
rect 32447 25245 32456 25279
rect 32404 25236 32456 25245
rect 32680 25236 32732 25288
rect 33508 25236 33560 25288
rect 33784 25236 33836 25288
rect 34980 25279 35032 25288
rect 34980 25245 34989 25279
rect 34989 25245 35023 25279
rect 35023 25245 35032 25279
rect 34980 25236 35032 25245
rect 35256 25236 35308 25288
rect 27436 25168 27488 25220
rect 29000 25168 29052 25220
rect 29368 25168 29420 25220
rect 25688 25143 25740 25152
rect 25688 25109 25697 25143
rect 25697 25109 25731 25143
rect 25731 25109 25740 25143
rect 25688 25100 25740 25109
rect 26148 25100 26200 25152
rect 26884 25143 26936 25152
rect 26884 25109 26893 25143
rect 26893 25109 26927 25143
rect 26927 25109 26936 25143
rect 26884 25100 26936 25109
rect 28816 25143 28868 25152
rect 28816 25109 28825 25143
rect 28825 25109 28859 25143
rect 28859 25109 28868 25143
rect 28816 25100 28868 25109
rect 29644 25100 29696 25152
rect 33692 25168 33744 25220
rect 34612 25168 34664 25220
rect 35348 25168 35400 25220
rect 36268 25236 36320 25288
rect 36636 25236 36688 25288
rect 37832 25236 37884 25288
rect 38384 25279 38436 25288
rect 38384 25245 38393 25279
rect 38393 25245 38427 25279
rect 38427 25245 38436 25279
rect 38384 25236 38436 25245
rect 36728 25168 36780 25220
rect 37372 25168 37424 25220
rect 38292 25211 38344 25220
rect 38292 25177 38301 25211
rect 38301 25177 38335 25211
rect 38335 25177 38344 25211
rect 38292 25168 38344 25177
rect 39212 25372 39264 25424
rect 40040 25372 40092 25424
rect 39212 25279 39264 25288
rect 39212 25245 39221 25279
rect 39221 25245 39255 25279
rect 39255 25245 39264 25279
rect 39212 25236 39264 25245
rect 39304 25236 39356 25288
rect 35440 25100 35492 25152
rect 37464 25143 37516 25152
rect 37464 25109 37473 25143
rect 37473 25109 37507 25143
rect 37507 25109 37516 25143
rect 37464 25100 37516 25109
rect 39120 25100 39172 25152
rect 39580 25168 39632 25220
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40500 25372 40552 25424
rect 40040 25236 40092 25245
rect 41880 25372 41932 25424
rect 41236 25347 41288 25356
rect 41236 25313 41245 25347
rect 41245 25313 41279 25347
rect 41279 25313 41288 25347
rect 41236 25304 41288 25313
rect 41512 25236 41564 25288
rect 42064 25236 42116 25288
rect 42432 25168 42484 25220
rect 41972 25100 42024 25152
rect 42524 25100 42576 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 15844 24896 15896 24948
rect 19432 24939 19484 24948
rect 19432 24905 19441 24939
rect 19441 24905 19475 24939
rect 19475 24905 19484 24939
rect 19432 24896 19484 24905
rect 20904 24896 20956 24948
rect 21916 24896 21968 24948
rect 17040 24828 17092 24880
rect 17500 24871 17552 24880
rect 17500 24837 17534 24871
rect 17534 24837 17552 24871
rect 17500 24828 17552 24837
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 16028 24803 16080 24812
rect 16028 24769 16037 24803
rect 16037 24769 16071 24803
rect 16071 24769 16080 24803
rect 16028 24760 16080 24769
rect 13268 24692 13320 24744
rect 18328 24760 18380 24812
rect 20812 24760 20864 24812
rect 20904 24803 20956 24812
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 20904 24760 20956 24769
rect 24032 24896 24084 24948
rect 24584 24896 24636 24948
rect 14648 24556 14700 24608
rect 21364 24692 21416 24744
rect 23112 24760 23164 24812
rect 23480 24828 23532 24880
rect 24952 24896 25004 24948
rect 27620 24896 27672 24948
rect 31576 24896 31628 24948
rect 31760 24896 31812 24948
rect 32312 24939 32364 24948
rect 32312 24905 32321 24939
rect 32321 24905 32355 24939
rect 32355 24905 32364 24939
rect 32312 24896 32364 24905
rect 34704 24896 34756 24948
rect 28816 24828 28868 24880
rect 29092 24828 29144 24880
rect 23572 24692 23624 24744
rect 23848 24735 23900 24744
rect 23848 24701 23857 24735
rect 23857 24701 23891 24735
rect 23891 24701 23900 24735
rect 23848 24692 23900 24701
rect 24216 24735 24268 24744
rect 24216 24701 24225 24735
rect 24225 24701 24259 24735
rect 24259 24701 24268 24735
rect 24216 24692 24268 24701
rect 24032 24624 24084 24676
rect 24584 24692 24636 24744
rect 26700 24760 26752 24812
rect 27160 24760 27212 24812
rect 27252 24803 27304 24812
rect 27252 24769 27261 24803
rect 27261 24769 27295 24803
rect 27295 24769 27304 24803
rect 27252 24760 27304 24769
rect 28172 24760 28224 24812
rect 25228 24735 25280 24744
rect 25228 24701 25237 24735
rect 25237 24701 25271 24735
rect 25271 24701 25280 24735
rect 25228 24692 25280 24701
rect 29368 24760 29420 24812
rect 29736 24760 29788 24812
rect 29920 24803 29972 24812
rect 29920 24769 29929 24803
rect 29929 24769 29963 24803
rect 29963 24769 29972 24803
rect 29920 24760 29972 24769
rect 30380 24828 30432 24880
rect 30104 24760 30156 24812
rect 30840 24760 30892 24812
rect 31392 24760 31444 24812
rect 32128 24760 32180 24812
rect 32404 24760 32456 24812
rect 32680 24735 32732 24744
rect 32680 24701 32689 24735
rect 32689 24701 32723 24735
rect 32723 24701 32732 24735
rect 32680 24692 32732 24701
rect 18420 24556 18472 24608
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 20812 24556 20864 24608
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 21456 24556 21508 24608
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23664 24599 23716 24608
rect 23664 24565 23673 24599
rect 23673 24565 23707 24599
rect 23707 24565 23716 24599
rect 23664 24556 23716 24565
rect 24216 24556 24268 24608
rect 24860 24556 24912 24608
rect 25136 24624 25188 24676
rect 28080 24624 28132 24676
rect 29460 24624 29512 24676
rect 32588 24667 32640 24676
rect 32588 24633 32597 24667
rect 32597 24633 32631 24667
rect 32631 24633 32640 24667
rect 32588 24624 32640 24633
rect 33784 24760 33836 24812
rect 33600 24692 33652 24744
rect 34520 24803 34572 24812
rect 34520 24769 34529 24803
rect 34529 24769 34563 24803
rect 34563 24769 34572 24803
rect 34520 24760 34572 24769
rect 35900 24828 35952 24880
rect 37832 24896 37884 24948
rect 34980 24760 35032 24812
rect 35348 24760 35400 24812
rect 35624 24760 35676 24812
rect 36544 24760 36596 24812
rect 36636 24803 36688 24812
rect 36636 24769 36645 24803
rect 36645 24769 36679 24803
rect 36679 24769 36688 24803
rect 36636 24760 36688 24769
rect 37740 24760 37792 24812
rect 35992 24735 36044 24744
rect 35992 24701 36001 24735
rect 36001 24701 36035 24735
rect 36035 24701 36044 24735
rect 35992 24692 36044 24701
rect 37096 24692 37148 24744
rect 40040 24760 40092 24812
rect 40132 24803 40184 24812
rect 40132 24769 40141 24803
rect 40141 24769 40175 24803
rect 40175 24769 40184 24803
rect 40132 24760 40184 24769
rect 34428 24624 34480 24676
rect 35072 24624 35124 24676
rect 35256 24624 35308 24676
rect 35624 24624 35676 24676
rect 37740 24667 37792 24676
rect 37740 24633 37749 24667
rect 37749 24633 37783 24667
rect 37783 24633 37792 24667
rect 37740 24624 37792 24633
rect 37832 24624 37884 24676
rect 38016 24624 38068 24676
rect 39488 24735 39540 24744
rect 39488 24701 39497 24735
rect 39497 24701 39531 24735
rect 39531 24701 39540 24735
rect 39488 24692 39540 24701
rect 39672 24692 39724 24744
rect 41788 24828 41840 24880
rect 42984 24871 43036 24880
rect 42984 24837 42993 24871
rect 42993 24837 43027 24871
rect 43027 24837 43036 24871
rect 42984 24828 43036 24837
rect 40316 24803 40368 24812
rect 40316 24769 40325 24803
rect 40325 24769 40359 24803
rect 40359 24769 40368 24803
rect 40316 24760 40368 24769
rect 40500 24760 40552 24812
rect 41144 24760 41196 24812
rect 28264 24556 28316 24608
rect 29736 24599 29788 24608
rect 29736 24565 29745 24599
rect 29745 24565 29779 24599
rect 29779 24565 29788 24599
rect 29736 24556 29788 24565
rect 30748 24556 30800 24608
rect 31668 24556 31720 24608
rect 34520 24556 34572 24608
rect 34704 24599 34756 24608
rect 34704 24565 34713 24599
rect 34713 24565 34747 24599
rect 34747 24565 34756 24599
rect 34704 24556 34756 24565
rect 35716 24556 35768 24608
rect 36452 24599 36504 24608
rect 36452 24565 36461 24599
rect 36461 24565 36495 24599
rect 36495 24565 36504 24599
rect 36452 24556 36504 24565
rect 36912 24599 36964 24608
rect 36912 24565 36921 24599
rect 36921 24565 36955 24599
rect 36955 24565 36964 24599
rect 36912 24556 36964 24565
rect 39028 24556 39080 24608
rect 39488 24556 39540 24608
rect 41236 24692 41288 24744
rect 41972 24803 42024 24812
rect 41972 24769 41981 24803
rect 41981 24769 42015 24803
rect 42015 24769 42024 24803
rect 41972 24760 42024 24769
rect 42616 24803 42668 24812
rect 42616 24769 42625 24803
rect 42625 24769 42659 24803
rect 42659 24769 42668 24803
rect 42616 24760 42668 24769
rect 42892 24803 42944 24812
rect 42892 24769 42901 24803
rect 42901 24769 42935 24803
rect 42935 24769 42944 24803
rect 42892 24760 42944 24769
rect 43076 24803 43128 24812
rect 43076 24769 43085 24803
rect 43085 24769 43119 24803
rect 43119 24769 43128 24803
rect 43076 24760 43128 24769
rect 42432 24692 42484 24744
rect 40500 24624 40552 24676
rect 41880 24599 41932 24608
rect 41880 24565 41889 24599
rect 41889 24565 41923 24599
rect 41923 24565 41932 24599
rect 41880 24556 41932 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12900 24352 12952 24404
rect 17684 24395 17736 24404
rect 17684 24361 17693 24395
rect 17693 24361 17727 24395
rect 17727 24361 17736 24395
rect 17684 24352 17736 24361
rect 20352 24352 20404 24404
rect 20628 24284 20680 24336
rect 15108 24216 15160 24268
rect 18328 24259 18380 24268
rect 18328 24225 18337 24259
rect 18337 24225 18371 24259
rect 18371 24225 18380 24259
rect 18328 24216 18380 24225
rect 21732 24352 21784 24404
rect 23664 24352 23716 24404
rect 23848 24352 23900 24404
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 24860 24352 24912 24404
rect 28632 24352 28684 24404
rect 29920 24352 29972 24404
rect 33048 24352 33100 24404
rect 35348 24352 35400 24404
rect 35808 24352 35860 24404
rect 35900 24352 35952 24404
rect 36544 24352 36596 24404
rect 21824 24284 21876 24336
rect 22560 24284 22612 24336
rect 23112 24327 23164 24336
rect 23112 24293 23121 24327
rect 23121 24293 23155 24327
rect 23155 24293 23164 24327
rect 23112 24284 23164 24293
rect 16028 24148 16080 24200
rect 20076 24148 20128 24200
rect 18604 24080 18656 24132
rect 20720 24191 20772 24200
rect 20720 24157 20729 24191
rect 20729 24157 20763 24191
rect 20763 24157 20772 24191
rect 20720 24148 20772 24157
rect 21088 24080 21140 24132
rect 21824 24191 21876 24200
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 22560 24191 22612 24200
rect 22560 24157 22569 24191
rect 22569 24157 22603 24191
rect 22603 24157 22612 24191
rect 22560 24148 22612 24157
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 24032 24191 24084 24200
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 24492 24148 24544 24200
rect 25228 24148 25280 24200
rect 22928 24080 22980 24132
rect 24216 24080 24268 24132
rect 26608 24191 26660 24200
rect 26608 24157 26617 24191
rect 26617 24157 26651 24191
rect 26651 24157 26660 24191
rect 26608 24148 26660 24157
rect 32496 24284 32548 24336
rect 33508 24284 33560 24336
rect 28172 24216 28224 24268
rect 29736 24216 29788 24268
rect 27160 24148 27212 24200
rect 27712 24191 27764 24200
rect 27712 24157 27721 24191
rect 27721 24157 27755 24191
rect 27755 24157 27764 24191
rect 27712 24148 27764 24157
rect 27896 24191 27948 24200
rect 27896 24157 27905 24191
rect 27905 24157 27939 24191
rect 27939 24157 27948 24191
rect 27896 24148 27948 24157
rect 28080 24148 28132 24200
rect 29460 24148 29512 24200
rect 30932 24216 30984 24268
rect 31484 24216 31536 24268
rect 31576 24259 31628 24268
rect 31576 24225 31585 24259
rect 31585 24225 31619 24259
rect 31619 24225 31628 24259
rect 31576 24216 31628 24225
rect 33232 24216 33284 24268
rect 30196 24148 30248 24200
rect 31300 24148 31352 24200
rect 32772 24148 32824 24200
rect 33600 24191 33652 24200
rect 33600 24157 33609 24191
rect 33609 24157 33643 24191
rect 33643 24157 33652 24191
rect 33600 24148 33652 24157
rect 33876 24259 33928 24268
rect 33876 24225 33885 24259
rect 33885 24225 33919 24259
rect 33919 24225 33928 24259
rect 33876 24216 33928 24225
rect 35716 24284 35768 24336
rect 37096 24284 37148 24336
rect 37372 24395 37424 24404
rect 37372 24361 37381 24395
rect 37381 24361 37415 24395
rect 37415 24361 37424 24395
rect 37372 24352 37424 24361
rect 37464 24352 37516 24404
rect 40040 24395 40092 24404
rect 40040 24361 40049 24395
rect 40049 24361 40083 24395
rect 40083 24361 40092 24395
rect 40040 24352 40092 24361
rect 40408 24395 40460 24404
rect 40408 24361 40417 24395
rect 40417 24361 40451 24395
rect 40451 24361 40460 24395
rect 40408 24352 40460 24361
rect 41236 24395 41288 24404
rect 41236 24361 41245 24395
rect 41245 24361 41279 24395
rect 41279 24361 41288 24395
rect 41236 24352 41288 24361
rect 42064 24395 42116 24404
rect 42064 24361 42073 24395
rect 42073 24361 42107 24395
rect 42107 24361 42116 24395
rect 42064 24352 42116 24361
rect 34336 24216 34388 24268
rect 34244 24191 34296 24200
rect 34244 24157 34253 24191
rect 34253 24157 34287 24191
rect 34287 24157 34296 24191
rect 34244 24148 34296 24157
rect 34428 24148 34480 24200
rect 29184 24080 29236 24132
rect 14648 24055 14700 24064
rect 14648 24021 14657 24055
rect 14657 24021 14691 24055
rect 14691 24021 14700 24055
rect 14648 24012 14700 24021
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 20720 24012 20772 24064
rect 20904 24055 20956 24064
rect 20904 24021 20913 24055
rect 20913 24021 20947 24055
rect 20947 24021 20956 24055
rect 20904 24012 20956 24021
rect 21364 24055 21416 24064
rect 21364 24021 21373 24055
rect 21373 24021 21407 24055
rect 21407 24021 21416 24055
rect 21364 24012 21416 24021
rect 22560 24012 22612 24064
rect 25136 24055 25188 24064
rect 25136 24021 25145 24055
rect 25145 24021 25179 24055
rect 25179 24021 25188 24055
rect 25136 24012 25188 24021
rect 27344 24012 27396 24064
rect 30288 24012 30340 24064
rect 31392 24080 31444 24132
rect 34152 24012 34204 24064
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 36268 24148 36320 24200
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 37004 24148 37056 24200
rect 37648 24191 37700 24200
rect 37648 24157 37657 24191
rect 37657 24157 37691 24191
rect 37691 24157 37700 24191
rect 37648 24148 37700 24157
rect 38016 24148 38068 24200
rect 38384 24148 38436 24200
rect 41328 24216 41380 24268
rect 41696 24216 41748 24268
rect 42892 24216 42944 24268
rect 39396 24148 39448 24200
rect 39672 24148 39724 24200
rect 40132 24191 40184 24200
rect 40132 24157 40141 24191
rect 40141 24157 40175 24191
rect 40175 24157 40184 24191
rect 40132 24148 40184 24157
rect 41788 24148 41840 24200
rect 42432 24148 42484 24200
rect 43352 24148 43404 24200
rect 43996 24148 44048 24200
rect 36452 24012 36504 24064
rect 37832 24080 37884 24132
rect 41696 24080 41748 24132
rect 38016 24012 38068 24064
rect 38476 24055 38528 24064
rect 38476 24021 38485 24055
rect 38485 24021 38519 24055
rect 38519 24021 38528 24055
rect 38476 24012 38528 24021
rect 38568 24012 38620 24064
rect 40960 24012 41012 24064
rect 42340 24012 42392 24064
rect 42524 24012 42576 24064
rect 42984 24012 43036 24064
rect 43168 24055 43220 24064
rect 43168 24021 43177 24055
rect 43177 24021 43211 24055
rect 43211 24021 43220 24055
rect 43168 24012 43220 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 14464 23808 14516 23860
rect 14740 23808 14792 23860
rect 18144 23808 18196 23860
rect 21732 23808 21784 23860
rect 14648 23740 14700 23792
rect 14832 23672 14884 23724
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 17868 23740 17920 23792
rect 15108 23604 15160 23656
rect 15384 23604 15436 23656
rect 17684 23715 17736 23724
rect 17684 23681 17693 23715
rect 17693 23681 17727 23715
rect 17727 23681 17736 23715
rect 17684 23672 17736 23681
rect 20996 23783 21048 23792
rect 20996 23749 21005 23783
rect 21005 23749 21039 23783
rect 21039 23749 21048 23783
rect 20996 23740 21048 23749
rect 21824 23740 21876 23792
rect 25872 23808 25924 23860
rect 26424 23808 26476 23860
rect 17224 23604 17276 23656
rect 18972 23715 19024 23724
rect 18972 23681 18981 23715
rect 18981 23681 19015 23715
rect 19015 23681 19024 23715
rect 18972 23672 19024 23681
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 21364 23672 21416 23724
rect 22376 23783 22428 23792
rect 22376 23749 22385 23783
rect 22385 23749 22419 23783
rect 22419 23749 22428 23783
rect 22376 23740 22428 23749
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 18604 23647 18656 23656
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 21272 23604 21324 23656
rect 24308 23740 24360 23792
rect 24952 23740 25004 23792
rect 27620 23740 27672 23792
rect 24492 23672 24544 23724
rect 25964 23672 26016 23724
rect 27804 23672 27856 23724
rect 27896 23715 27948 23724
rect 27896 23681 27905 23715
rect 27905 23681 27939 23715
rect 27939 23681 27948 23715
rect 27896 23672 27948 23681
rect 23756 23604 23808 23656
rect 27712 23604 27764 23656
rect 29184 23740 29236 23792
rect 29460 23740 29512 23792
rect 30288 23851 30340 23860
rect 30288 23817 30297 23851
rect 30297 23817 30331 23851
rect 30331 23817 30340 23851
rect 30288 23808 30340 23817
rect 30748 23851 30800 23860
rect 30748 23817 30757 23851
rect 30757 23817 30791 23851
rect 30791 23817 30800 23851
rect 30748 23808 30800 23817
rect 34336 23851 34388 23860
rect 34336 23817 34345 23851
rect 34345 23817 34379 23851
rect 34379 23817 34388 23851
rect 34336 23808 34388 23817
rect 34796 23808 34848 23860
rect 35348 23808 35400 23860
rect 28908 23672 28960 23724
rect 28632 23604 28684 23656
rect 30104 23740 30156 23792
rect 30196 23740 30248 23792
rect 31852 23740 31904 23792
rect 32496 23740 32548 23792
rect 33692 23740 33744 23792
rect 30380 23672 30432 23724
rect 30840 23672 30892 23724
rect 31208 23715 31260 23724
rect 31208 23681 31217 23715
rect 31217 23681 31251 23715
rect 31251 23681 31260 23715
rect 31208 23672 31260 23681
rect 32680 23672 32732 23724
rect 33508 23715 33560 23724
rect 33508 23681 33517 23715
rect 33517 23681 33551 23715
rect 33551 23681 33560 23715
rect 33508 23672 33560 23681
rect 34152 23672 34204 23724
rect 34244 23715 34296 23724
rect 34244 23681 34253 23715
rect 34253 23681 34287 23715
rect 34287 23681 34296 23715
rect 34244 23672 34296 23681
rect 34704 23740 34756 23792
rect 16304 23468 16356 23520
rect 20076 23468 20128 23520
rect 22560 23468 22612 23520
rect 23480 23468 23532 23520
rect 24952 23536 25004 23588
rect 26608 23536 26660 23588
rect 27436 23536 27488 23588
rect 26700 23468 26752 23520
rect 27160 23511 27212 23520
rect 27160 23477 27169 23511
rect 27169 23477 27203 23511
rect 27203 23477 27212 23511
rect 27160 23468 27212 23477
rect 27252 23468 27304 23520
rect 27620 23468 27672 23520
rect 29000 23536 29052 23588
rect 30288 23604 30340 23656
rect 31116 23647 31168 23656
rect 31116 23613 31125 23647
rect 31125 23613 31159 23647
rect 31159 23613 31168 23647
rect 31116 23604 31168 23613
rect 32036 23604 32088 23656
rect 35440 23672 35492 23724
rect 35716 23672 35768 23724
rect 36268 23672 36320 23724
rect 36544 23672 36596 23724
rect 37832 23740 37884 23792
rect 39028 23783 39080 23792
rect 39028 23749 39037 23783
rect 39037 23749 39071 23783
rect 39071 23749 39080 23783
rect 39028 23740 39080 23749
rect 39212 23740 39264 23792
rect 38292 23672 38344 23724
rect 39488 23715 39540 23724
rect 39488 23681 39497 23715
rect 39497 23681 39531 23715
rect 39531 23681 39540 23715
rect 39488 23672 39540 23681
rect 39672 23851 39724 23860
rect 39672 23817 39681 23851
rect 39681 23817 39715 23851
rect 39715 23817 39724 23851
rect 39672 23808 39724 23817
rect 40684 23851 40736 23860
rect 40684 23817 40693 23851
rect 40693 23817 40727 23851
rect 40727 23817 40736 23851
rect 40684 23808 40736 23817
rect 42984 23851 43036 23860
rect 42984 23817 42993 23851
rect 42993 23817 43027 23851
rect 43027 23817 43036 23851
rect 42984 23808 43036 23817
rect 42340 23740 42392 23792
rect 41512 23715 41564 23724
rect 41512 23681 41521 23715
rect 41521 23681 41555 23715
rect 41555 23681 41564 23715
rect 41512 23672 41564 23681
rect 42800 23715 42852 23724
rect 42800 23681 42809 23715
rect 42809 23681 42843 23715
rect 42843 23681 42852 23715
rect 42800 23672 42852 23681
rect 35348 23604 35400 23656
rect 35624 23604 35676 23656
rect 37096 23604 37148 23656
rect 37464 23604 37516 23656
rect 37832 23604 37884 23656
rect 40684 23604 40736 23656
rect 32864 23536 32916 23588
rect 35440 23536 35492 23588
rect 35808 23536 35860 23588
rect 36452 23536 36504 23588
rect 41144 23536 41196 23588
rect 29552 23468 29604 23520
rect 32312 23468 32364 23520
rect 32404 23511 32456 23520
rect 32404 23477 32413 23511
rect 32413 23477 32447 23511
rect 32447 23477 32456 23511
rect 32404 23468 32456 23477
rect 35900 23468 35952 23520
rect 37464 23511 37516 23520
rect 37464 23477 37473 23511
rect 37473 23477 37507 23511
rect 37507 23477 37516 23511
rect 37464 23468 37516 23477
rect 37648 23511 37700 23520
rect 37648 23477 37657 23511
rect 37657 23477 37691 23511
rect 37691 23477 37700 23511
rect 37648 23468 37700 23477
rect 38384 23468 38436 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17684 23264 17736 23316
rect 15476 23196 15528 23248
rect 18236 23196 18288 23248
rect 14280 23060 14332 23112
rect 15752 23128 15804 23180
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 20812 23264 20864 23316
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 22836 23264 22888 23316
rect 25964 23307 26016 23316
rect 25964 23273 25973 23307
rect 25973 23273 26007 23307
rect 26007 23273 26016 23307
rect 25964 23264 26016 23273
rect 28908 23264 28960 23316
rect 31392 23264 31444 23316
rect 33232 23264 33284 23316
rect 33508 23264 33560 23316
rect 33968 23307 34020 23316
rect 33968 23273 33977 23307
rect 33977 23273 34011 23307
rect 34011 23273 34020 23307
rect 33968 23264 34020 23273
rect 36728 23264 36780 23316
rect 38476 23264 38528 23316
rect 38660 23264 38712 23316
rect 39212 23264 39264 23316
rect 40224 23307 40276 23316
rect 40224 23273 40233 23307
rect 40233 23273 40267 23307
rect 40267 23273 40276 23307
rect 40224 23264 40276 23273
rect 41512 23264 41564 23316
rect 41788 23264 41840 23316
rect 42892 23264 42944 23316
rect 31300 23196 31352 23248
rect 37096 23196 37148 23248
rect 23756 23171 23808 23180
rect 23756 23137 23765 23171
rect 23765 23137 23799 23171
rect 23799 23137 23808 23171
rect 23756 23128 23808 23137
rect 24768 23171 24820 23180
rect 24768 23137 24777 23171
rect 24777 23137 24811 23171
rect 24811 23137 24820 23171
rect 24768 23128 24820 23137
rect 25136 23128 25188 23180
rect 27160 23128 27212 23180
rect 27804 23128 27856 23180
rect 31944 23128 31996 23180
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 15568 22992 15620 23044
rect 13544 22924 13596 22976
rect 14832 22924 14884 22976
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 17224 23103 17276 23112
rect 17224 23069 17233 23103
rect 17233 23069 17267 23103
rect 17267 23069 17276 23103
rect 17224 23060 17276 23069
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 18604 23060 18656 23112
rect 19340 23060 19392 23112
rect 19984 23060 20036 23112
rect 20904 23060 20956 23112
rect 23480 23103 23532 23112
rect 23480 23069 23498 23103
rect 23498 23069 23532 23103
rect 23480 23060 23532 23069
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 26424 23060 26476 23112
rect 27344 23103 27396 23112
rect 27344 23069 27353 23103
rect 27353 23069 27387 23103
rect 27387 23069 27396 23103
rect 27344 23060 27396 23069
rect 28356 23060 28408 23112
rect 17684 22992 17736 23044
rect 19064 22992 19116 23044
rect 28908 23060 28960 23112
rect 18512 22924 18564 22976
rect 20996 22967 21048 22976
rect 20996 22933 21005 22967
rect 21005 22933 21039 22967
rect 21039 22933 21048 22967
rect 20996 22924 21048 22933
rect 24032 22924 24084 22976
rect 28172 22967 28224 22976
rect 28172 22933 28181 22967
rect 28181 22933 28215 22967
rect 28215 22933 28224 22967
rect 28172 22924 28224 22933
rect 28908 22924 28960 22976
rect 33140 23060 33192 23112
rect 33876 23060 33928 23112
rect 34704 23128 34756 23180
rect 34796 23060 34848 23112
rect 30288 22992 30340 23044
rect 30196 22924 30248 22976
rect 31668 22967 31720 22976
rect 31668 22933 31677 22967
rect 31677 22933 31711 22967
rect 31711 22933 31720 22967
rect 31668 22924 31720 22933
rect 31944 23035 31996 23044
rect 31944 23001 31953 23035
rect 31953 23001 31987 23035
rect 31987 23001 31996 23035
rect 31944 22992 31996 23001
rect 33600 23035 33652 23044
rect 33600 23001 33609 23035
rect 33609 23001 33643 23035
rect 33643 23001 33652 23035
rect 33600 22992 33652 23001
rect 33784 23035 33836 23044
rect 33784 23001 33793 23035
rect 33793 23001 33827 23035
rect 33827 23001 33836 23035
rect 33784 22992 33836 23001
rect 34980 23103 35032 23112
rect 34980 23069 34989 23103
rect 34989 23069 35023 23103
rect 35023 23069 35032 23103
rect 34980 23060 35032 23069
rect 37832 23128 37884 23180
rect 35992 23060 36044 23112
rect 35624 22992 35676 23044
rect 36820 23035 36872 23044
rect 36820 23001 36829 23035
rect 36829 23001 36863 23035
rect 36863 23001 36872 23035
rect 36820 22992 36872 23001
rect 37188 23060 37240 23112
rect 37556 23060 37608 23112
rect 38752 23128 38804 23180
rect 38844 23128 38896 23180
rect 39304 23128 39356 23180
rect 43076 23196 43128 23248
rect 41972 23128 42024 23180
rect 42892 23128 42944 23180
rect 38568 23060 38620 23112
rect 39212 23103 39264 23112
rect 39212 23069 39221 23103
rect 39221 23069 39255 23103
rect 39255 23069 39264 23103
rect 39212 23060 39264 23069
rect 36268 22924 36320 22976
rect 37556 22924 37608 22976
rect 37648 22924 37700 22976
rect 38292 22992 38344 23044
rect 39304 22924 39356 22976
rect 39488 23060 39540 23112
rect 41880 23103 41932 23112
rect 41880 23069 41889 23103
rect 41889 23069 41923 23103
rect 41923 23069 41932 23103
rect 41880 23060 41932 23069
rect 42708 23060 42760 23112
rect 39764 22992 39816 23044
rect 42432 22992 42484 23044
rect 43076 22992 43128 23044
rect 39672 22924 39724 22976
rect 39948 22924 40000 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 15476 22720 15528 22772
rect 16028 22763 16080 22772
rect 16028 22729 16037 22763
rect 16037 22729 16071 22763
rect 16071 22729 16080 22763
rect 16028 22720 16080 22729
rect 18972 22720 19024 22772
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 24492 22720 24544 22772
rect 17592 22652 17644 22704
rect 18420 22652 18472 22704
rect 13544 22627 13596 22636
rect 13544 22593 13578 22627
rect 13578 22593 13596 22627
rect 13544 22584 13596 22593
rect 13268 22559 13320 22568
rect 13268 22525 13277 22559
rect 13277 22525 13311 22559
rect 13311 22525 13320 22559
rect 13268 22516 13320 22525
rect 18052 22584 18104 22636
rect 18512 22627 18564 22636
rect 19984 22652 20036 22704
rect 18512 22593 18530 22627
rect 18530 22593 18564 22627
rect 18512 22584 18564 22593
rect 20812 22584 20864 22636
rect 14372 22448 14424 22500
rect 14924 22448 14976 22500
rect 20904 22448 20956 22500
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 27620 22652 27672 22704
rect 28356 22763 28408 22772
rect 28356 22729 28365 22763
rect 28365 22729 28399 22763
rect 28399 22729 28408 22763
rect 28356 22720 28408 22729
rect 29368 22763 29420 22772
rect 29368 22729 29377 22763
rect 29377 22729 29411 22763
rect 29411 22729 29420 22763
rect 29368 22720 29420 22729
rect 30288 22720 30340 22772
rect 30380 22763 30432 22772
rect 30380 22729 30389 22763
rect 30389 22729 30423 22763
rect 30423 22729 30432 22763
rect 30380 22720 30432 22729
rect 30472 22720 30524 22772
rect 32220 22720 32272 22772
rect 32496 22763 32548 22772
rect 32496 22729 32505 22763
rect 32505 22729 32539 22763
rect 32539 22729 32548 22763
rect 32496 22720 32548 22729
rect 33416 22720 33468 22772
rect 30104 22652 30156 22704
rect 25412 22627 25464 22636
rect 25412 22593 25421 22627
rect 25421 22593 25455 22627
rect 25455 22593 25464 22627
rect 25412 22584 25464 22593
rect 27252 22627 27304 22636
rect 27252 22593 27261 22627
rect 27261 22593 27295 22627
rect 27295 22593 27304 22627
rect 27252 22584 27304 22593
rect 28172 22584 28224 22636
rect 31300 22652 31352 22704
rect 32956 22652 33008 22704
rect 30748 22627 30800 22636
rect 30748 22593 30757 22627
rect 30757 22593 30791 22627
rect 30791 22593 30800 22627
rect 30748 22584 30800 22593
rect 33140 22584 33192 22636
rect 34060 22720 34112 22772
rect 34336 22720 34388 22772
rect 34796 22720 34848 22772
rect 34888 22720 34940 22772
rect 33784 22652 33836 22704
rect 33968 22652 34020 22704
rect 36820 22763 36872 22772
rect 36820 22729 36829 22763
rect 36829 22729 36863 22763
rect 36863 22729 36872 22763
rect 36820 22720 36872 22729
rect 37924 22720 37976 22772
rect 38384 22720 38436 22772
rect 38936 22720 38988 22772
rect 39488 22720 39540 22772
rect 42340 22720 42392 22772
rect 39672 22652 39724 22704
rect 41788 22652 41840 22704
rect 42064 22652 42116 22704
rect 22928 22559 22980 22568
rect 22928 22525 22937 22559
rect 22937 22525 22971 22559
rect 22971 22525 22980 22559
rect 22928 22516 22980 22525
rect 24860 22516 24912 22568
rect 25688 22448 25740 22500
rect 26332 22448 26384 22500
rect 27804 22491 27856 22500
rect 27804 22457 27813 22491
rect 27813 22457 27847 22491
rect 27847 22457 27856 22491
rect 27804 22448 27856 22457
rect 28816 22448 28868 22500
rect 31024 22559 31076 22568
rect 31024 22525 31033 22559
rect 31033 22525 31067 22559
rect 31067 22525 31076 22559
rect 31024 22516 31076 22525
rect 14464 22380 14516 22432
rect 15200 22380 15252 22432
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 22376 22380 22428 22432
rect 22652 22380 22704 22432
rect 26884 22380 26936 22432
rect 30472 22380 30524 22432
rect 31576 22423 31628 22432
rect 31576 22389 31585 22423
rect 31585 22389 31619 22423
rect 31619 22389 31628 22423
rect 31576 22380 31628 22389
rect 32312 22491 32364 22500
rect 32312 22457 32321 22491
rect 32321 22457 32355 22491
rect 32355 22457 32364 22491
rect 32312 22448 32364 22457
rect 32864 22423 32916 22432
rect 32864 22389 32873 22423
rect 32873 22389 32907 22423
rect 32907 22389 32916 22423
rect 32864 22380 32916 22389
rect 33600 22448 33652 22500
rect 35624 22627 35676 22636
rect 35624 22593 35633 22627
rect 35633 22593 35667 22627
rect 35667 22593 35676 22627
rect 35624 22584 35676 22593
rect 35900 22627 35952 22636
rect 35900 22593 35909 22627
rect 35909 22593 35943 22627
rect 35943 22593 35952 22627
rect 35900 22584 35952 22593
rect 36084 22627 36136 22636
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 36636 22627 36688 22636
rect 36636 22593 36645 22627
rect 36645 22593 36679 22627
rect 36679 22593 36688 22627
rect 36636 22584 36688 22593
rect 36820 22627 36872 22636
rect 36820 22593 36829 22627
rect 36829 22593 36863 22627
rect 36863 22593 36872 22627
rect 36820 22584 36872 22593
rect 37004 22584 37056 22636
rect 37556 22584 37608 22636
rect 37924 22584 37976 22636
rect 38200 22584 38252 22636
rect 39212 22627 39264 22636
rect 39212 22593 39221 22627
rect 39221 22593 39255 22627
rect 39255 22593 39264 22627
rect 39212 22584 39264 22593
rect 39396 22584 39448 22636
rect 40868 22627 40920 22636
rect 40868 22593 40877 22627
rect 40877 22593 40911 22627
rect 40911 22593 40920 22627
rect 40868 22584 40920 22593
rect 42248 22584 42300 22636
rect 43076 22627 43128 22636
rect 43076 22593 43085 22627
rect 43085 22593 43119 22627
rect 43119 22593 43128 22627
rect 43076 22584 43128 22593
rect 43260 22584 43312 22636
rect 35808 22516 35860 22568
rect 42984 22559 43036 22568
rect 42984 22525 42993 22559
rect 42993 22525 43027 22559
rect 43027 22525 43036 22559
rect 42984 22516 43036 22525
rect 38844 22448 38896 22500
rect 39304 22448 39356 22500
rect 39488 22448 39540 22500
rect 34888 22380 34940 22432
rect 34980 22380 35032 22432
rect 35900 22380 35952 22432
rect 35992 22423 36044 22432
rect 35992 22389 36001 22423
rect 36001 22389 36035 22423
rect 36035 22389 36044 22423
rect 35992 22380 36044 22389
rect 36544 22380 36596 22432
rect 39028 22380 39080 22432
rect 40408 22448 40460 22500
rect 40040 22380 40092 22432
rect 41788 22380 41840 22432
rect 42156 22380 42208 22432
rect 42708 22423 42760 22432
rect 42708 22389 42717 22423
rect 42717 22389 42751 22423
rect 42751 22389 42760 22423
rect 42708 22380 42760 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 15476 22176 15528 22228
rect 14372 22108 14424 22160
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 14924 22083 14976 22092
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 15844 22176 15896 22228
rect 17592 22108 17644 22160
rect 18604 22151 18656 22160
rect 18604 22117 18613 22151
rect 18613 22117 18647 22151
rect 18647 22117 18656 22151
rect 18604 22108 18656 22117
rect 19340 22176 19392 22228
rect 22008 22176 22060 22228
rect 24860 22176 24912 22228
rect 18052 22083 18104 22092
rect 18052 22049 18061 22083
rect 18061 22049 18095 22083
rect 18095 22049 18104 22083
rect 18052 22040 18104 22049
rect 18144 22083 18196 22092
rect 18144 22049 18153 22083
rect 18153 22049 18187 22083
rect 18187 22049 18196 22083
rect 18144 22040 18196 22049
rect 20812 22040 20864 22092
rect 21916 22040 21968 22092
rect 14464 21972 14516 22024
rect 18972 21972 19024 22024
rect 20720 21972 20772 22024
rect 15384 21904 15436 21956
rect 20260 21904 20312 21956
rect 22100 22015 22152 22024
rect 22100 21981 22109 22015
rect 22109 21981 22143 22015
rect 22143 21981 22152 22015
rect 22100 21972 22152 21981
rect 23756 22108 23808 22160
rect 28908 22176 28960 22228
rect 29000 22108 29052 22160
rect 29736 22151 29788 22160
rect 29736 22117 29745 22151
rect 29745 22117 29779 22151
rect 29779 22117 29788 22151
rect 29736 22108 29788 22117
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 26792 21972 26844 22024
rect 28540 21972 28592 22024
rect 30748 22176 30800 22228
rect 34796 22176 34848 22228
rect 35164 22176 35216 22228
rect 35440 22176 35492 22228
rect 39028 22176 39080 22228
rect 39304 22219 39356 22228
rect 39304 22185 39313 22219
rect 39313 22185 39347 22219
rect 39347 22185 39356 22219
rect 39304 22176 39356 22185
rect 42524 22176 42576 22228
rect 42984 22176 43036 22228
rect 31576 22108 31628 22160
rect 32036 22151 32088 22160
rect 32036 22117 32045 22151
rect 32045 22117 32079 22151
rect 32079 22117 32088 22151
rect 32036 22108 32088 22117
rect 35808 22108 35860 22160
rect 30104 22040 30156 22092
rect 33876 22083 33928 22092
rect 33876 22049 33885 22083
rect 33885 22049 33919 22083
rect 33919 22049 33928 22083
rect 33876 22040 33928 22049
rect 35624 22040 35676 22092
rect 36452 22108 36504 22160
rect 36084 22040 36136 22092
rect 36544 22083 36596 22092
rect 36544 22049 36553 22083
rect 36553 22049 36587 22083
rect 36587 22049 36596 22083
rect 36544 22040 36596 22049
rect 23848 21904 23900 21956
rect 25412 21904 25464 21956
rect 28080 21904 28132 21956
rect 28908 21904 28960 21956
rect 30196 21904 30248 21956
rect 14740 21836 14792 21888
rect 19432 21836 19484 21888
rect 19984 21836 20036 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23020 21836 23072 21888
rect 25688 21836 25740 21888
rect 28724 21879 28776 21888
rect 28724 21845 28733 21879
rect 28733 21845 28767 21879
rect 28767 21845 28776 21879
rect 28724 21836 28776 21845
rect 30932 22015 30984 22024
rect 30932 21981 30941 22015
rect 30941 21981 30975 22015
rect 30975 21981 30984 22015
rect 30932 21972 30984 21981
rect 31116 21972 31168 22024
rect 32036 21972 32088 22024
rect 32496 22015 32548 22024
rect 32496 21981 32505 22015
rect 32505 21981 32539 22015
rect 32539 21981 32548 22015
rect 32496 21972 32548 21981
rect 32956 22015 33008 22024
rect 32956 21981 32965 22015
rect 32965 21981 32999 22015
rect 32999 21981 33008 22015
rect 32956 21972 33008 21981
rect 33416 22015 33468 22024
rect 33416 21981 33425 22015
rect 33425 21981 33459 22015
rect 33459 21981 33468 22015
rect 33416 21972 33468 21981
rect 36360 22015 36412 22024
rect 36360 21981 36369 22015
rect 36369 21981 36403 22015
rect 36403 21981 36412 22015
rect 36360 21972 36412 21981
rect 36636 22015 36688 22024
rect 36636 21981 36645 22015
rect 36645 21981 36679 22015
rect 36679 21981 36688 22015
rect 36636 21972 36688 21981
rect 39948 22108 40000 22160
rect 38200 22040 38252 22092
rect 37188 21972 37240 22024
rect 37464 21972 37516 22024
rect 31392 21836 31444 21888
rect 31668 21836 31720 21888
rect 34336 21836 34388 21888
rect 36084 21904 36136 21956
rect 37740 21904 37792 21956
rect 38016 21972 38068 22024
rect 38568 22015 38620 22024
rect 38568 21981 38577 22015
rect 38577 21981 38611 22015
rect 38611 21981 38620 22015
rect 38568 21972 38620 21981
rect 39120 22040 39172 22092
rect 38844 21972 38896 22024
rect 40316 22040 40368 22092
rect 41788 22083 41840 22092
rect 41788 22049 41797 22083
rect 41797 22049 41831 22083
rect 41831 22049 41840 22083
rect 41788 22040 41840 22049
rect 38108 21879 38160 21888
rect 38108 21845 38117 21879
rect 38117 21845 38151 21879
rect 38151 21845 38160 21879
rect 38108 21836 38160 21845
rect 39120 21904 39172 21956
rect 40224 22015 40276 22024
rect 40224 21981 40233 22015
rect 40233 21981 40267 22015
rect 40267 21981 40276 22015
rect 40224 21972 40276 21981
rect 42156 21904 42208 21956
rect 39304 21836 39356 21888
rect 39672 21836 39724 21888
rect 40684 21879 40736 21888
rect 40684 21845 40693 21879
rect 40693 21845 40727 21879
rect 40727 21845 40736 21879
rect 40684 21836 40736 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 14740 21675 14792 21684
rect 14740 21641 14749 21675
rect 14749 21641 14783 21675
rect 14783 21641 14792 21675
rect 14740 21632 14792 21641
rect 15292 21632 15344 21684
rect 20996 21632 21048 21684
rect 13268 21564 13320 21616
rect 15844 21564 15896 21616
rect 19432 21564 19484 21616
rect 20904 21607 20956 21616
rect 20904 21573 20913 21607
rect 20913 21573 20947 21607
rect 20947 21573 20956 21607
rect 20904 21564 20956 21573
rect 22284 21607 22336 21616
rect 22284 21573 22318 21607
rect 22318 21573 22336 21607
rect 22284 21564 22336 21573
rect 23848 21675 23900 21684
rect 23848 21641 23857 21675
rect 23857 21641 23891 21675
rect 23891 21641 23900 21675
rect 23848 21632 23900 21641
rect 25504 21632 25556 21684
rect 28080 21632 28132 21684
rect 28908 21632 28960 21684
rect 29828 21632 29880 21684
rect 30104 21632 30156 21684
rect 12532 21428 12584 21480
rect 14740 21496 14792 21548
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 15752 21496 15804 21548
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 17132 21539 17184 21548
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 19984 21496 20036 21548
rect 29736 21564 29788 21616
rect 34612 21632 34664 21684
rect 36084 21632 36136 21684
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 22008 21471 22060 21480
rect 22008 21437 22017 21471
rect 22017 21437 22051 21471
rect 22051 21437 22060 21471
rect 22008 21428 22060 21437
rect 18236 21360 18288 21412
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 17500 21292 17552 21344
rect 18052 21292 18104 21344
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 20352 21292 20404 21344
rect 23388 21335 23440 21344
rect 23388 21301 23397 21335
rect 23397 21301 23431 21335
rect 23431 21301 23440 21335
rect 23388 21292 23440 21301
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 26884 21496 26936 21548
rect 27068 21496 27120 21548
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 29368 21496 29420 21548
rect 30564 21539 30616 21548
rect 30564 21505 30573 21539
rect 30573 21505 30607 21539
rect 30607 21505 30616 21539
rect 30564 21496 30616 21505
rect 32404 21564 32456 21616
rect 31024 21496 31076 21548
rect 32864 21539 32916 21548
rect 32864 21505 32873 21539
rect 32873 21505 32907 21539
rect 32907 21505 32916 21539
rect 32864 21496 32916 21505
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 33140 21471 33192 21480
rect 33140 21437 33149 21471
rect 33149 21437 33183 21471
rect 33183 21437 33192 21471
rect 33140 21428 33192 21437
rect 35716 21607 35768 21616
rect 35716 21573 35725 21607
rect 35725 21573 35759 21607
rect 35759 21573 35768 21607
rect 35716 21564 35768 21573
rect 36912 21564 36964 21616
rect 33600 21496 33652 21548
rect 33968 21496 34020 21548
rect 34796 21496 34848 21548
rect 35164 21496 35216 21548
rect 35440 21539 35492 21548
rect 35440 21505 35449 21539
rect 35449 21505 35483 21539
rect 35483 21505 35492 21539
rect 35440 21496 35492 21505
rect 28172 21360 28224 21412
rect 30840 21360 30892 21412
rect 31576 21360 31628 21412
rect 32680 21360 32732 21412
rect 33508 21360 33560 21412
rect 35808 21539 35860 21548
rect 35808 21505 35817 21539
rect 35817 21505 35851 21539
rect 35851 21505 35860 21539
rect 35808 21496 35860 21505
rect 35992 21496 36044 21548
rect 35716 21428 35768 21480
rect 37372 21428 37424 21480
rect 34060 21360 34112 21412
rect 38844 21632 38896 21684
rect 40868 21632 40920 21684
rect 42064 21675 42116 21684
rect 42064 21641 42073 21675
rect 42073 21641 42107 21675
rect 42107 21641 42116 21675
rect 42064 21632 42116 21641
rect 43352 21675 43404 21684
rect 43352 21641 43361 21675
rect 43361 21641 43395 21675
rect 43395 21641 43404 21675
rect 43352 21632 43404 21641
rect 40040 21564 40092 21616
rect 40500 21564 40552 21616
rect 40684 21564 40736 21616
rect 38108 21496 38160 21548
rect 38752 21496 38804 21548
rect 39580 21496 39632 21548
rect 40316 21539 40368 21548
rect 40316 21505 40325 21539
rect 40325 21505 40359 21539
rect 40359 21505 40368 21539
rect 40316 21496 40368 21505
rect 42248 21496 42300 21548
rect 38476 21471 38528 21480
rect 38476 21437 38485 21471
rect 38485 21437 38519 21471
rect 38519 21437 38528 21471
rect 38476 21428 38528 21437
rect 33048 21292 33100 21344
rect 35532 21292 35584 21344
rect 35624 21292 35676 21344
rect 35900 21292 35952 21344
rect 37004 21292 37056 21344
rect 37464 21335 37516 21344
rect 37464 21301 37473 21335
rect 37473 21301 37507 21335
rect 37507 21301 37516 21335
rect 37464 21292 37516 21301
rect 39212 21292 39264 21344
rect 39672 21335 39724 21344
rect 39672 21301 39681 21335
rect 39681 21301 39715 21335
rect 39715 21301 39724 21335
rect 39672 21292 39724 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 15384 21131 15436 21140
rect 15384 21097 15393 21131
rect 15393 21097 15427 21131
rect 15427 21097 15436 21131
rect 15384 21088 15436 21097
rect 17132 21088 17184 21140
rect 22100 21131 22152 21140
rect 22100 21097 22109 21131
rect 22109 21097 22143 21131
rect 22143 21097 22152 21131
rect 22100 21088 22152 21097
rect 22284 21088 22336 21140
rect 24860 21088 24912 21140
rect 25504 21088 25556 21140
rect 25964 21131 26016 21140
rect 25964 21097 25973 21131
rect 25973 21097 26007 21131
rect 26007 21097 26016 21131
rect 25964 21088 26016 21097
rect 26332 21088 26384 21140
rect 27620 21088 27672 21140
rect 28172 21131 28224 21140
rect 28172 21097 28181 21131
rect 28181 21097 28215 21131
rect 28215 21097 28224 21131
rect 28172 21088 28224 21097
rect 28540 21088 28592 21140
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18236 20952 18288 20961
rect 18328 20952 18380 21004
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 16120 20927 16172 20936
rect 16120 20893 16154 20927
rect 16154 20893 16172 20927
rect 16120 20884 16172 20893
rect 19064 20884 19116 20936
rect 15108 20816 15160 20868
rect 20444 20816 20496 20868
rect 13820 20748 13872 20800
rect 14372 20748 14424 20800
rect 16580 20748 16632 20800
rect 17776 20748 17828 20800
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 22284 20884 22336 20936
rect 22744 20884 22796 20936
rect 23388 20884 23440 20936
rect 23480 20927 23532 20936
rect 23480 20893 23489 20927
rect 23489 20893 23523 20927
rect 23523 20893 23532 20927
rect 23480 20884 23532 20893
rect 23572 20927 23624 20936
rect 23572 20893 23581 20927
rect 23581 20893 23615 20927
rect 23615 20893 23624 20927
rect 23572 20884 23624 20893
rect 22560 20859 22612 20868
rect 22560 20825 22569 20859
rect 22569 20825 22603 20859
rect 22603 20825 22612 20859
rect 22560 20816 22612 20825
rect 24584 20995 24636 21004
rect 24584 20961 24593 20995
rect 24593 20961 24627 20995
rect 24627 20961 24636 20995
rect 24584 20952 24636 20961
rect 24308 20884 24360 20936
rect 24676 20884 24728 20936
rect 29092 20952 29144 21004
rect 27620 20884 27672 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 28816 20884 28868 20936
rect 27160 20816 27212 20868
rect 33140 21088 33192 21140
rect 34336 21131 34388 21140
rect 34336 21097 34345 21131
rect 34345 21097 34379 21131
rect 34379 21097 34388 21131
rect 34336 21088 34388 21097
rect 31484 21020 31536 21072
rect 35808 21088 35860 21140
rect 35900 21088 35952 21140
rect 36360 21020 36412 21072
rect 36728 21131 36780 21140
rect 36728 21097 36737 21131
rect 36737 21097 36771 21131
rect 36771 21097 36780 21131
rect 36728 21088 36780 21097
rect 37464 21088 37516 21140
rect 39856 21088 39908 21140
rect 40040 21088 40092 21140
rect 40224 21088 40276 21140
rect 31760 20884 31812 20936
rect 32220 20884 32272 20936
rect 33140 20952 33192 21004
rect 32864 20884 32916 20936
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 33048 20927 33100 20936
rect 33048 20893 33057 20927
rect 33057 20893 33091 20927
rect 33091 20893 33100 20927
rect 33048 20884 33100 20893
rect 35624 20952 35676 21004
rect 35992 20952 36044 21004
rect 37832 21020 37884 21072
rect 40500 21020 40552 21072
rect 38476 20952 38528 21004
rect 39028 20995 39080 21004
rect 39028 20961 39037 20995
rect 39037 20961 39071 20995
rect 39071 20961 39080 20995
rect 39028 20952 39080 20961
rect 35532 20884 35584 20936
rect 36728 20927 36780 20936
rect 36728 20893 36737 20927
rect 36737 20893 36771 20927
rect 36771 20893 36780 20927
rect 36728 20884 36780 20893
rect 37924 20884 37976 20936
rect 38752 20884 38804 20936
rect 24768 20748 24820 20800
rect 30380 20816 30432 20868
rect 35900 20816 35952 20868
rect 37556 20859 37608 20868
rect 37556 20825 37565 20859
rect 37565 20825 37599 20859
rect 37599 20825 37608 20859
rect 37556 20816 37608 20825
rect 37740 20816 37792 20868
rect 39212 20884 39264 20936
rect 40132 20884 40184 20936
rect 40500 20927 40552 20936
rect 40500 20893 40509 20927
rect 40509 20893 40543 20927
rect 40543 20893 40552 20927
rect 40500 20884 40552 20893
rect 29092 20748 29144 20800
rect 31024 20748 31076 20800
rect 32772 20748 32824 20800
rect 35440 20748 35492 20800
rect 35808 20748 35860 20800
rect 38016 20748 38068 20800
rect 39028 20748 39080 20800
rect 40408 20816 40460 20868
rect 41328 20816 41380 20868
rect 43352 20816 43404 20868
rect 43996 20816 44048 20868
rect 42248 20791 42300 20800
rect 42248 20757 42257 20791
rect 42257 20757 42291 20791
rect 42291 20757 42300 20791
rect 42248 20748 42300 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 17224 20544 17276 20596
rect 19984 20544 20036 20596
rect 20444 20587 20496 20596
rect 20444 20553 20453 20587
rect 20453 20553 20487 20587
rect 20487 20553 20496 20587
rect 20444 20544 20496 20553
rect 22744 20544 22796 20596
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 13452 20340 13504 20392
rect 18236 20476 18288 20528
rect 20720 20476 20772 20528
rect 20904 20476 20956 20528
rect 15108 20340 15160 20392
rect 15568 20408 15620 20460
rect 15936 20408 15988 20460
rect 17684 20451 17736 20460
rect 17684 20417 17693 20451
rect 17693 20417 17727 20451
rect 17727 20417 17736 20451
rect 17684 20408 17736 20417
rect 17776 20408 17828 20460
rect 19064 20408 19116 20460
rect 19432 20408 19484 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 23664 20476 23716 20528
rect 15752 20340 15804 20392
rect 15476 20272 15528 20324
rect 15660 20272 15712 20324
rect 17960 20340 18012 20392
rect 21640 20340 21692 20392
rect 23756 20408 23808 20460
rect 27436 20544 27488 20596
rect 27528 20544 27580 20596
rect 28356 20544 28408 20596
rect 25688 20519 25740 20528
rect 25688 20485 25697 20519
rect 25697 20485 25731 20519
rect 25731 20485 25740 20519
rect 25688 20476 25740 20485
rect 27160 20476 27212 20528
rect 29092 20519 29144 20528
rect 29092 20485 29101 20519
rect 29101 20485 29135 20519
rect 29135 20485 29144 20519
rect 29092 20476 29144 20485
rect 30564 20587 30616 20596
rect 30564 20553 30573 20587
rect 30573 20553 30607 20587
rect 30607 20553 30616 20587
rect 30564 20544 30616 20553
rect 32220 20544 32272 20596
rect 34796 20544 34848 20596
rect 37464 20544 37516 20596
rect 40132 20544 40184 20596
rect 40316 20544 40368 20596
rect 42708 20544 42760 20596
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 27620 20408 27672 20460
rect 13176 20247 13228 20256
rect 13176 20213 13185 20247
rect 13185 20213 13219 20247
rect 13219 20213 13228 20247
rect 13176 20204 13228 20213
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 15292 20204 15344 20256
rect 18144 20272 18196 20324
rect 18788 20272 18840 20324
rect 18328 20204 18380 20256
rect 19340 20272 19392 20324
rect 23572 20272 23624 20324
rect 27896 20340 27948 20392
rect 27988 20340 28040 20392
rect 28908 20408 28960 20460
rect 30748 20340 30800 20392
rect 31668 20476 31720 20528
rect 31116 20451 31168 20460
rect 31116 20417 31125 20451
rect 31125 20417 31159 20451
rect 31159 20417 31168 20451
rect 31116 20408 31168 20417
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 32404 20408 32456 20460
rect 32588 20451 32640 20460
rect 32588 20417 32597 20451
rect 32597 20417 32631 20451
rect 32631 20417 32640 20451
rect 32588 20408 32640 20417
rect 32772 20408 32824 20460
rect 33048 20408 33100 20460
rect 33876 20451 33928 20460
rect 33876 20417 33910 20451
rect 33910 20417 33928 20451
rect 33876 20408 33928 20417
rect 35348 20408 35400 20460
rect 36912 20451 36964 20460
rect 36912 20417 36921 20451
rect 36921 20417 36955 20451
rect 36955 20417 36964 20451
rect 36912 20408 36964 20417
rect 37648 20451 37700 20460
rect 37648 20417 37657 20451
rect 37657 20417 37691 20451
rect 37691 20417 37700 20451
rect 37648 20408 37700 20417
rect 38016 20408 38068 20460
rect 33508 20340 33560 20392
rect 34612 20340 34664 20392
rect 36176 20340 36228 20392
rect 38936 20383 38988 20392
rect 38936 20349 38945 20383
rect 38945 20349 38979 20383
rect 38979 20349 38988 20383
rect 38936 20340 38988 20349
rect 39212 20408 39264 20460
rect 41880 20476 41932 20528
rect 42248 20408 42300 20460
rect 40500 20383 40552 20392
rect 40500 20349 40509 20383
rect 40509 20349 40543 20383
rect 40543 20349 40552 20383
rect 40500 20340 40552 20349
rect 28816 20272 28868 20324
rect 32404 20272 32456 20324
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 22468 20204 22520 20256
rect 27344 20247 27396 20256
rect 27344 20213 27353 20247
rect 27353 20213 27387 20247
rect 27387 20213 27396 20247
rect 27344 20204 27396 20213
rect 28356 20247 28408 20256
rect 28356 20213 28365 20247
rect 28365 20213 28399 20247
rect 28399 20213 28408 20247
rect 28356 20204 28408 20213
rect 28908 20204 28960 20256
rect 30104 20247 30156 20256
rect 30104 20213 30113 20247
rect 30113 20213 30147 20247
rect 30147 20213 30156 20247
rect 30104 20204 30156 20213
rect 31024 20247 31076 20256
rect 31024 20213 31033 20247
rect 31033 20213 31067 20247
rect 31067 20213 31076 20247
rect 31024 20204 31076 20213
rect 31392 20204 31444 20256
rect 32772 20204 32824 20256
rect 37372 20272 37424 20324
rect 34612 20204 34664 20256
rect 34704 20204 34756 20256
rect 35624 20204 35676 20256
rect 37464 20204 37516 20256
rect 37648 20247 37700 20256
rect 37648 20213 37657 20247
rect 37657 20213 37691 20247
rect 37691 20213 37700 20247
rect 37648 20204 37700 20213
rect 38016 20247 38068 20256
rect 38016 20213 38025 20247
rect 38025 20213 38059 20247
rect 38059 20213 38068 20247
rect 38016 20204 38068 20213
rect 39120 20272 39172 20324
rect 42892 20247 42944 20256
rect 42892 20213 42901 20247
rect 42901 20213 42935 20247
rect 42935 20213 42944 20247
rect 42892 20204 42944 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 12992 20043 13044 20052
rect 12992 20009 13001 20043
rect 13001 20009 13035 20043
rect 13035 20009 13044 20043
rect 12992 20000 13044 20009
rect 14648 20000 14700 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 16304 20000 16356 20052
rect 18788 20043 18840 20052
rect 18788 20009 18797 20043
rect 18797 20009 18831 20043
rect 18831 20009 18840 20043
rect 18788 20000 18840 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 21640 20043 21692 20052
rect 21640 20009 21649 20043
rect 21649 20009 21683 20043
rect 21683 20009 21692 20043
rect 21640 20000 21692 20009
rect 22192 20000 22244 20052
rect 23664 20000 23716 20052
rect 23940 20000 23992 20052
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 16948 19864 17000 19916
rect 13360 19796 13412 19848
rect 13820 19728 13872 19780
rect 15844 19796 15896 19848
rect 17500 19796 17552 19848
rect 19984 19864 20036 19916
rect 24308 19932 24360 19984
rect 26148 19932 26200 19984
rect 28264 20043 28316 20052
rect 28264 20009 28273 20043
rect 28273 20009 28307 20043
rect 28307 20009 28316 20043
rect 28264 20000 28316 20009
rect 28724 20043 28776 20052
rect 28724 20009 28733 20043
rect 28733 20009 28767 20043
rect 28767 20009 28776 20043
rect 28724 20000 28776 20009
rect 30104 20000 30156 20052
rect 30380 20043 30432 20052
rect 30380 20009 30389 20043
rect 30389 20009 30423 20043
rect 30423 20009 30432 20043
rect 30380 20000 30432 20009
rect 32128 20000 32180 20052
rect 33876 20043 33928 20052
rect 33876 20009 33885 20043
rect 33885 20009 33919 20043
rect 33919 20009 33928 20043
rect 33876 20000 33928 20009
rect 34888 20000 34940 20052
rect 31576 19932 31628 19984
rect 34612 19932 34664 19984
rect 36728 20000 36780 20052
rect 38568 20000 38620 20052
rect 40500 20000 40552 20052
rect 43260 20043 43312 20052
rect 43260 20009 43269 20043
rect 43269 20009 43303 20043
rect 43303 20009 43312 20043
rect 43260 20000 43312 20009
rect 23572 19907 23624 19916
rect 23572 19873 23581 19907
rect 23581 19873 23615 19907
rect 23615 19873 23624 19907
rect 23572 19864 23624 19873
rect 16856 19728 16908 19780
rect 17868 19728 17920 19780
rect 22008 19796 22060 19848
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22468 19796 22520 19805
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 23756 19796 23808 19848
rect 24492 19796 24544 19848
rect 24860 19864 24912 19916
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 27436 19796 27488 19848
rect 28816 19864 28868 19916
rect 28908 19864 28960 19916
rect 31116 19864 31168 19916
rect 34796 19864 34848 19916
rect 37648 19932 37700 19984
rect 37832 19932 37884 19984
rect 40408 19932 40460 19984
rect 20904 19728 20956 19780
rect 15568 19660 15620 19712
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 18236 19660 18288 19712
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 23664 19660 23716 19712
rect 27252 19660 27304 19712
rect 27988 19771 28040 19780
rect 27988 19737 27997 19771
rect 27997 19737 28031 19771
rect 28031 19737 28040 19771
rect 27988 19728 28040 19737
rect 29184 19796 29236 19848
rect 30840 19796 30892 19848
rect 31024 19796 31076 19848
rect 31760 19839 31812 19848
rect 31760 19805 31769 19839
rect 31769 19805 31803 19839
rect 31803 19805 31812 19839
rect 31760 19796 31812 19805
rect 33048 19796 33100 19848
rect 38016 19864 38068 19916
rect 28172 19728 28224 19780
rect 29368 19728 29420 19780
rect 31852 19728 31904 19780
rect 34704 19728 34756 19780
rect 36452 19839 36504 19848
rect 36452 19805 36461 19839
rect 36461 19805 36495 19839
rect 36495 19805 36504 19839
rect 36452 19796 36504 19805
rect 36544 19796 36596 19848
rect 37188 19796 37240 19848
rect 37280 19796 37332 19848
rect 37740 19796 37792 19848
rect 36912 19728 36964 19780
rect 37372 19728 37424 19780
rect 38660 19796 38712 19848
rect 38568 19728 38620 19780
rect 39028 19839 39080 19848
rect 39028 19805 39037 19839
rect 39037 19805 39071 19839
rect 39071 19805 39080 19839
rect 39028 19796 39080 19805
rect 40316 19864 40368 19916
rect 42892 19796 42944 19848
rect 35440 19660 35492 19712
rect 39304 19660 39356 19712
rect 39948 19660 40000 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 15568 19456 15620 19508
rect 15936 19499 15988 19508
rect 15936 19465 15945 19499
rect 15945 19465 15979 19499
rect 15979 19465 15988 19499
rect 15936 19456 15988 19465
rect 17960 19456 18012 19508
rect 18604 19456 18656 19508
rect 19984 19456 20036 19508
rect 20076 19456 20128 19508
rect 22744 19499 22796 19508
rect 22744 19465 22753 19499
rect 22753 19465 22787 19499
rect 22787 19465 22796 19499
rect 22744 19456 22796 19465
rect 23664 19499 23716 19508
rect 23664 19465 23673 19499
rect 23673 19465 23707 19499
rect 23707 19465 23716 19499
rect 23664 19456 23716 19465
rect 24124 19499 24176 19508
rect 24124 19465 24133 19499
rect 24133 19465 24167 19499
rect 24167 19465 24176 19499
rect 24124 19456 24176 19465
rect 26516 19456 26568 19508
rect 27988 19456 28040 19508
rect 28356 19456 28408 19508
rect 28908 19456 28960 19508
rect 13176 19388 13228 19440
rect 15384 19388 15436 19440
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 15292 19320 15344 19329
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 15752 19388 15804 19440
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16948 19320 17000 19372
rect 20720 19388 20772 19440
rect 21180 19388 21232 19440
rect 28264 19431 28316 19440
rect 28264 19397 28282 19431
rect 28282 19397 28316 19431
rect 28264 19388 28316 19397
rect 29368 19431 29420 19440
rect 29368 19397 29377 19431
rect 29377 19397 29411 19431
rect 29411 19397 29420 19431
rect 29368 19388 29420 19397
rect 30104 19388 30156 19440
rect 31668 19456 31720 19508
rect 31852 19456 31904 19508
rect 33968 19456 34020 19508
rect 35808 19456 35860 19508
rect 18328 19363 18380 19372
rect 18328 19329 18337 19363
rect 18337 19329 18371 19363
rect 18371 19329 18380 19363
rect 18328 19320 18380 19329
rect 19984 19320 20036 19372
rect 22008 19320 22060 19372
rect 22284 19320 22336 19372
rect 18972 19252 19024 19304
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 23940 19252 23992 19304
rect 24584 19252 24636 19304
rect 27804 19320 27856 19372
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 30380 19320 30432 19372
rect 31576 19363 31628 19372
rect 31576 19329 31585 19363
rect 31585 19329 31619 19363
rect 31619 19329 31628 19363
rect 31576 19320 31628 19329
rect 33508 19388 33560 19440
rect 36912 19456 36964 19508
rect 38292 19456 38344 19508
rect 37096 19388 37148 19440
rect 39120 19456 39172 19508
rect 40132 19456 40184 19508
rect 41880 19499 41932 19508
rect 41880 19465 41889 19499
rect 41889 19465 41923 19499
rect 41923 19465 41932 19499
rect 41880 19456 41932 19465
rect 32128 19320 32180 19372
rect 28540 19295 28592 19304
rect 28540 19261 28549 19295
rect 28549 19261 28583 19295
rect 28583 19261 28592 19295
rect 28540 19252 28592 19261
rect 29000 19252 29052 19304
rect 30012 19252 30064 19304
rect 33048 19320 33100 19372
rect 34060 19363 34112 19372
rect 34060 19329 34094 19363
rect 34094 19329 34112 19363
rect 34060 19320 34112 19329
rect 35992 19320 36044 19372
rect 37740 19320 37792 19372
rect 38568 19388 38620 19440
rect 39672 19388 39724 19440
rect 39948 19388 40000 19440
rect 39028 19320 39080 19372
rect 35900 19252 35952 19304
rect 37188 19252 37240 19304
rect 38936 19252 38988 19304
rect 39212 19363 39264 19372
rect 39212 19329 39221 19363
rect 39221 19329 39255 19363
rect 39255 19329 39264 19363
rect 39212 19320 39264 19329
rect 39304 19320 39356 19372
rect 39672 19252 39724 19304
rect 40132 19320 40184 19372
rect 40684 19363 40736 19372
rect 40684 19329 40693 19363
rect 40693 19329 40727 19363
rect 40727 19329 40736 19363
rect 40684 19320 40736 19329
rect 40776 19363 40828 19372
rect 40776 19329 40785 19363
rect 40785 19329 40819 19363
rect 40819 19329 40828 19363
rect 40776 19320 40828 19329
rect 41052 19320 41104 19372
rect 42248 19320 42300 19372
rect 40316 19252 40368 19304
rect 21272 19184 21324 19236
rect 31760 19184 31812 19236
rect 32312 19184 32364 19236
rect 39764 19184 39816 19236
rect 40040 19227 40092 19236
rect 40040 19193 40049 19227
rect 40049 19193 40083 19227
rect 40083 19193 40092 19227
rect 40040 19184 40092 19193
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 29092 19116 29144 19168
rect 37648 19159 37700 19168
rect 37648 19125 37657 19159
rect 37657 19125 37691 19159
rect 37691 19125 37700 19159
rect 37648 19116 37700 19125
rect 40960 19159 41012 19168
rect 40960 19125 40969 19159
rect 40969 19125 41003 19159
rect 41003 19125 41012 19159
rect 40960 19116 41012 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 15200 18955 15252 18964
rect 15200 18921 15209 18955
rect 15209 18921 15243 18955
rect 15243 18921 15252 18955
rect 15200 18912 15252 18921
rect 21088 18912 21140 18964
rect 17960 18776 18012 18828
rect 21272 18776 21324 18828
rect 17040 18708 17092 18760
rect 15384 18640 15436 18692
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 19156 18708 19208 18760
rect 20720 18708 20772 18760
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 22652 18708 22704 18760
rect 23848 18912 23900 18964
rect 29000 18912 29052 18964
rect 28356 18844 28408 18896
rect 31208 18912 31260 18964
rect 34060 18912 34112 18964
rect 35532 18912 35584 18964
rect 35624 18955 35676 18964
rect 35624 18921 35633 18955
rect 35633 18921 35667 18955
rect 35667 18921 35676 18955
rect 35624 18912 35676 18921
rect 36452 18912 36504 18964
rect 36912 18955 36964 18964
rect 36912 18921 36921 18955
rect 36921 18921 36955 18955
rect 36955 18921 36964 18955
rect 36912 18912 36964 18921
rect 37556 18955 37608 18964
rect 37556 18921 37565 18955
rect 37565 18921 37599 18955
rect 37599 18921 37608 18955
rect 37556 18912 37608 18921
rect 37924 18912 37976 18964
rect 39304 18955 39356 18964
rect 39304 18921 39313 18955
rect 39313 18921 39347 18955
rect 39347 18921 39356 18955
rect 39304 18912 39356 18921
rect 40684 18912 40736 18964
rect 40776 18912 40828 18964
rect 41788 18912 41840 18964
rect 19248 18640 19300 18692
rect 22008 18640 22060 18692
rect 24584 18708 24636 18760
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 28816 18776 28868 18828
rect 37372 18844 37424 18896
rect 38844 18844 38896 18896
rect 39672 18844 39724 18896
rect 17132 18572 17184 18624
rect 19432 18572 19484 18624
rect 19984 18572 20036 18624
rect 29184 18708 29236 18760
rect 29460 18708 29512 18760
rect 29552 18708 29604 18760
rect 32772 18751 32824 18760
rect 32772 18717 32790 18751
rect 32790 18717 32824 18751
rect 32772 18708 32824 18717
rect 32956 18708 33008 18760
rect 33600 18708 33652 18760
rect 28356 18640 28408 18692
rect 29092 18572 29144 18624
rect 31024 18640 31076 18692
rect 33968 18751 34020 18760
rect 33968 18717 33977 18751
rect 33977 18717 34011 18751
rect 34011 18717 34020 18751
rect 33968 18708 34020 18717
rect 40224 18776 40276 18828
rect 32588 18572 32640 18624
rect 34796 18640 34848 18692
rect 35624 18751 35676 18760
rect 35624 18717 35633 18751
rect 35633 18717 35667 18751
rect 35667 18717 35676 18751
rect 35624 18708 35676 18717
rect 35992 18640 36044 18692
rect 37096 18708 37148 18760
rect 37372 18751 37424 18760
rect 37372 18717 37381 18751
rect 37381 18717 37415 18751
rect 37415 18717 37424 18751
rect 37372 18708 37424 18717
rect 37556 18751 37608 18760
rect 37556 18717 37565 18751
rect 37565 18717 37599 18751
rect 37599 18717 37608 18751
rect 37556 18708 37608 18717
rect 37924 18708 37976 18760
rect 40132 18751 40184 18760
rect 40132 18717 40141 18751
rect 40141 18717 40175 18751
rect 40175 18717 40184 18751
rect 40132 18708 40184 18717
rect 41696 18708 41748 18760
rect 42616 18751 42668 18760
rect 42616 18717 42625 18751
rect 42625 18717 42659 18751
rect 42659 18717 42668 18751
rect 42616 18708 42668 18717
rect 37740 18640 37792 18692
rect 38660 18640 38712 18692
rect 39948 18640 40000 18692
rect 40776 18683 40828 18692
rect 40776 18649 40785 18683
rect 40785 18649 40819 18683
rect 40819 18649 40828 18683
rect 40776 18640 40828 18649
rect 41052 18640 41104 18692
rect 34704 18572 34756 18624
rect 36360 18572 36412 18624
rect 38936 18615 38988 18624
rect 38936 18581 38945 18615
rect 38945 18581 38979 18615
rect 38979 18581 38988 18615
rect 38936 18572 38988 18581
rect 39028 18615 39080 18624
rect 39028 18581 39037 18615
rect 39037 18581 39071 18615
rect 39071 18581 39080 18615
rect 39028 18572 39080 18581
rect 39120 18615 39172 18624
rect 39120 18581 39129 18615
rect 39129 18581 39163 18615
rect 39163 18581 39172 18615
rect 39120 18572 39172 18581
rect 41144 18615 41196 18624
rect 41144 18581 41153 18615
rect 41153 18581 41187 18615
rect 41187 18581 41196 18615
rect 41144 18572 41196 18581
rect 42248 18572 42300 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 15292 18368 15344 18420
rect 15752 18368 15804 18420
rect 19984 18368 20036 18420
rect 22560 18368 22612 18420
rect 25044 18411 25096 18420
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 27620 18368 27672 18420
rect 32312 18368 32364 18420
rect 34612 18368 34664 18420
rect 36452 18368 36504 18420
rect 37464 18368 37516 18420
rect 38016 18368 38068 18420
rect 39028 18368 39080 18420
rect 39212 18368 39264 18420
rect 42616 18411 42668 18420
rect 42616 18377 42625 18411
rect 42625 18377 42659 18411
rect 42659 18377 42668 18411
rect 42616 18368 42668 18377
rect 15384 18300 15436 18352
rect 20260 18300 20312 18352
rect 23480 18300 23532 18352
rect 29000 18343 29052 18352
rect 29000 18309 29009 18343
rect 29009 18309 29043 18343
rect 29043 18309 29052 18343
rect 29000 18300 29052 18309
rect 30748 18300 30800 18352
rect 31484 18343 31536 18352
rect 31484 18309 31493 18343
rect 31493 18309 31527 18343
rect 31527 18309 31536 18343
rect 33048 18343 33100 18352
rect 31484 18300 31536 18309
rect 33048 18309 33057 18343
rect 33057 18309 33091 18343
rect 33091 18309 33100 18343
rect 33048 18300 33100 18309
rect 35624 18300 35676 18352
rect 37924 18343 37976 18352
rect 37924 18309 37927 18343
rect 37927 18309 37961 18343
rect 37961 18309 37976 18343
rect 37924 18300 37976 18309
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 15568 18232 15620 18284
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 14924 18164 14976 18216
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 17960 18232 18012 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 19248 18232 19300 18284
rect 19892 18232 19944 18284
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 20812 18232 20864 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 21088 18232 21140 18284
rect 22744 18275 22796 18284
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 22836 18207 22888 18216
rect 22836 18173 22845 18207
rect 22845 18173 22879 18207
rect 22879 18173 22888 18207
rect 22836 18164 22888 18173
rect 22928 18207 22980 18216
rect 22928 18173 22937 18207
rect 22937 18173 22971 18207
rect 22971 18173 22980 18207
rect 23756 18232 23808 18284
rect 27436 18232 27488 18284
rect 29920 18275 29972 18284
rect 29920 18241 29954 18275
rect 29954 18241 29972 18275
rect 29920 18232 29972 18241
rect 22928 18164 22980 18173
rect 26700 18164 26752 18216
rect 27160 18164 27212 18216
rect 28540 18164 28592 18216
rect 29552 18164 29604 18216
rect 31944 18164 31996 18216
rect 32588 18232 32640 18284
rect 34428 18275 34480 18284
rect 34428 18241 34437 18275
rect 34437 18241 34471 18275
rect 34471 18241 34480 18275
rect 34428 18232 34480 18241
rect 34704 18232 34756 18284
rect 37740 18232 37792 18284
rect 40960 18300 41012 18352
rect 38844 18232 38896 18284
rect 32956 18164 33008 18216
rect 33600 18164 33652 18216
rect 15476 18028 15528 18080
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 20996 18096 21048 18148
rect 32496 18096 32548 18148
rect 34428 18096 34480 18148
rect 35716 18096 35768 18148
rect 36360 18139 36412 18148
rect 36360 18105 36369 18139
rect 36369 18105 36403 18139
rect 36403 18105 36412 18139
rect 36360 18096 36412 18105
rect 37556 18164 37608 18216
rect 39212 18232 39264 18284
rect 43536 18232 43588 18284
rect 39304 18164 39356 18216
rect 43076 18207 43128 18216
rect 43076 18173 43085 18207
rect 43085 18173 43119 18207
rect 43119 18173 43128 18207
rect 43076 18164 43128 18173
rect 21180 18028 21232 18080
rect 28172 18028 28224 18080
rect 28908 18028 28960 18080
rect 30656 18028 30708 18080
rect 30932 18028 30984 18080
rect 34520 18071 34572 18080
rect 34520 18037 34529 18071
rect 34529 18037 34563 18071
rect 34563 18037 34572 18071
rect 34520 18028 34572 18037
rect 36176 18071 36228 18080
rect 36176 18037 36185 18071
rect 36185 18037 36219 18071
rect 36219 18037 36228 18071
rect 36176 18028 36228 18037
rect 37188 18028 37240 18080
rect 37556 18071 37608 18080
rect 37556 18037 37565 18071
rect 37565 18037 37599 18071
rect 37599 18037 37608 18071
rect 37556 18028 37608 18037
rect 38752 18028 38804 18080
rect 42984 18096 43036 18148
rect 41328 18028 41380 18080
rect 41696 18028 41748 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19892 17867 19944 17876
rect 19892 17833 19901 17867
rect 19901 17833 19935 17867
rect 19935 17833 19944 17867
rect 19892 17824 19944 17833
rect 20076 17824 20128 17876
rect 20904 17824 20956 17876
rect 22284 17867 22336 17876
rect 22284 17833 22293 17867
rect 22293 17833 22327 17867
rect 22327 17833 22336 17867
rect 22284 17824 22336 17833
rect 23572 17867 23624 17876
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 23940 17756 23992 17808
rect 24492 17756 24544 17808
rect 13636 17688 13688 17740
rect 15016 17688 15068 17740
rect 17316 17731 17368 17740
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 17316 17688 17368 17697
rect 20536 17688 20588 17740
rect 24768 17824 24820 17876
rect 25320 17824 25372 17876
rect 25780 17824 25832 17876
rect 27436 17867 27488 17876
rect 27436 17833 27445 17867
rect 27445 17833 27479 17867
rect 27479 17833 27488 17867
rect 27436 17824 27488 17833
rect 27896 17824 27948 17876
rect 28816 17824 28868 17876
rect 29920 17824 29972 17876
rect 31484 17867 31536 17876
rect 31484 17833 31493 17867
rect 31493 17833 31527 17867
rect 31527 17833 31536 17867
rect 31484 17824 31536 17833
rect 33048 17824 33100 17876
rect 34612 17824 34664 17876
rect 35808 17867 35860 17876
rect 35808 17833 35817 17867
rect 35817 17833 35851 17867
rect 35851 17833 35860 17867
rect 35808 17824 35860 17833
rect 36268 17824 36320 17876
rect 37648 17824 37700 17876
rect 37924 17824 37976 17876
rect 39028 17824 39080 17876
rect 40132 17867 40184 17876
rect 40132 17833 40141 17867
rect 40141 17833 40175 17867
rect 40175 17833 40184 17867
rect 40132 17824 40184 17833
rect 42984 17824 43036 17876
rect 43076 17824 43128 17876
rect 27620 17756 27672 17808
rect 29460 17756 29512 17808
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17224 17620 17276 17672
rect 17960 17620 18012 17672
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 18604 17620 18656 17672
rect 19984 17552 20036 17604
rect 20536 17552 20588 17604
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 14648 17527 14700 17536
rect 14648 17493 14657 17527
rect 14657 17493 14691 17527
rect 14691 17493 14700 17527
rect 14648 17484 14700 17493
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 20904 17527 20956 17536
rect 20904 17493 20913 17527
rect 20913 17493 20947 17527
rect 20947 17493 20956 17527
rect 20904 17484 20956 17493
rect 21088 17527 21140 17536
rect 21088 17493 21115 17527
rect 21115 17493 21140 17527
rect 22928 17620 22980 17672
rect 21088 17484 21140 17493
rect 21456 17484 21508 17536
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 23940 17663 23992 17672
rect 23940 17629 23949 17663
rect 23949 17629 23983 17663
rect 23983 17629 23992 17663
rect 23940 17620 23992 17629
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 23388 17552 23440 17604
rect 25044 17552 25096 17604
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28356 17620 28408 17672
rect 30656 17688 30708 17740
rect 27804 17595 27856 17604
rect 27804 17561 27813 17595
rect 27813 17561 27847 17595
rect 27847 17561 27856 17595
rect 27804 17552 27856 17561
rect 30380 17663 30432 17672
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 30380 17620 30432 17629
rect 31944 17756 31996 17808
rect 34520 17688 34572 17740
rect 36268 17731 36320 17740
rect 36268 17697 36277 17731
rect 36277 17697 36311 17731
rect 36311 17697 36320 17731
rect 36268 17688 36320 17697
rect 37832 17731 37884 17740
rect 37832 17697 37841 17731
rect 37841 17697 37875 17731
rect 37875 17697 37884 17731
rect 37832 17688 37884 17697
rect 32864 17620 32916 17672
rect 33048 17663 33100 17672
rect 33048 17629 33057 17663
rect 33057 17629 33091 17663
rect 33091 17629 33100 17663
rect 33048 17620 33100 17629
rect 34152 17663 34204 17672
rect 34152 17629 34161 17663
rect 34161 17629 34195 17663
rect 34195 17629 34204 17663
rect 34152 17620 34204 17629
rect 34336 17663 34388 17672
rect 34336 17629 34345 17663
rect 34345 17629 34379 17663
rect 34379 17629 34388 17663
rect 34336 17620 34388 17629
rect 34428 17620 34480 17672
rect 36636 17663 36688 17672
rect 36636 17629 36645 17663
rect 36645 17629 36679 17663
rect 36679 17629 36688 17663
rect 36636 17620 36688 17629
rect 27988 17484 28040 17536
rect 28172 17484 28224 17536
rect 28632 17527 28684 17536
rect 28632 17493 28659 17527
rect 28659 17493 28684 17527
rect 28632 17484 28684 17493
rect 35900 17552 35952 17604
rect 37648 17663 37700 17672
rect 37648 17629 37657 17663
rect 37657 17629 37691 17663
rect 37691 17629 37700 17663
rect 37648 17620 37700 17629
rect 37740 17663 37792 17672
rect 37740 17629 37749 17663
rect 37749 17629 37783 17663
rect 37783 17629 37792 17663
rect 37740 17620 37792 17629
rect 37924 17620 37976 17672
rect 39120 17756 39172 17808
rect 41420 17688 41472 17740
rect 41972 17731 42024 17740
rect 41972 17697 41981 17731
rect 41981 17697 42015 17731
rect 42015 17697 42024 17731
rect 41972 17688 42024 17697
rect 38476 17552 38528 17604
rect 38844 17663 38896 17672
rect 38844 17629 38853 17663
rect 38853 17629 38887 17663
rect 38887 17629 38896 17663
rect 38844 17620 38896 17629
rect 40224 17620 40276 17672
rect 40316 17663 40368 17672
rect 40316 17629 40325 17663
rect 40325 17629 40359 17663
rect 40359 17629 40368 17663
rect 40316 17620 40368 17629
rect 41144 17663 41196 17672
rect 41144 17629 41153 17663
rect 41153 17629 41187 17663
rect 41187 17629 41196 17663
rect 41144 17620 41196 17629
rect 42248 17663 42300 17672
rect 42248 17629 42282 17663
rect 42282 17629 42300 17663
rect 42248 17620 42300 17629
rect 28908 17484 28960 17536
rect 32128 17484 32180 17536
rect 34796 17484 34848 17536
rect 36544 17527 36596 17536
rect 36544 17493 36553 17527
rect 36553 17493 36587 17527
rect 36587 17493 36596 17527
rect 36544 17484 36596 17493
rect 37740 17484 37792 17536
rect 37924 17484 37976 17536
rect 43536 17552 43588 17604
rect 38752 17484 38804 17536
rect 39488 17484 39540 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 14924 17280 14976 17332
rect 15568 17280 15620 17332
rect 18236 17323 18288 17332
rect 18236 17289 18245 17323
rect 18245 17289 18279 17323
rect 18279 17289 18288 17323
rect 18236 17280 18288 17289
rect 18696 17280 18748 17332
rect 20536 17323 20588 17332
rect 20536 17289 20545 17323
rect 20545 17289 20579 17323
rect 20579 17289 20588 17323
rect 20536 17280 20588 17289
rect 14280 17212 14332 17264
rect 14648 17212 14700 17264
rect 13544 17144 13596 17196
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 19248 17212 19300 17264
rect 24032 17280 24084 17332
rect 28356 17280 28408 17332
rect 28540 17323 28592 17332
rect 28540 17289 28549 17323
rect 28549 17289 28583 17323
rect 28583 17289 28592 17323
rect 28540 17280 28592 17289
rect 17132 17187 17184 17196
rect 16856 17144 16908 17153
rect 17132 17153 17166 17187
rect 17166 17153 17184 17187
rect 17132 17144 17184 17153
rect 19156 17187 19208 17196
rect 19156 17153 19165 17187
rect 19165 17153 19199 17187
rect 19199 17153 19208 17187
rect 19156 17144 19208 17153
rect 20904 17144 20956 17196
rect 24584 17212 24636 17264
rect 25136 17212 25188 17264
rect 29092 17212 29144 17264
rect 30748 17255 30800 17264
rect 30748 17221 30757 17255
rect 30757 17221 30791 17255
rect 30791 17221 30800 17255
rect 30748 17212 30800 17221
rect 13360 17076 13412 17128
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 25688 17144 25740 17196
rect 25780 17187 25832 17196
rect 25780 17153 25789 17187
rect 25789 17153 25823 17187
rect 25823 17153 25832 17187
rect 25780 17144 25832 17153
rect 27436 17187 27488 17196
rect 27436 17153 27470 17187
rect 27470 17153 27488 17187
rect 27436 17144 27488 17153
rect 29000 17187 29052 17196
rect 29000 17153 29009 17187
rect 29009 17153 29043 17187
rect 29043 17153 29052 17187
rect 29000 17144 29052 17153
rect 29736 17144 29788 17196
rect 31852 17280 31904 17332
rect 32864 17280 32916 17332
rect 36176 17280 36228 17332
rect 37648 17280 37700 17332
rect 39396 17280 39448 17332
rect 41052 17280 41104 17332
rect 41880 17280 41932 17332
rect 43076 17280 43128 17332
rect 34520 17212 34572 17264
rect 31392 17187 31444 17196
rect 31392 17153 31401 17187
rect 31401 17153 31435 17187
rect 31435 17153 31444 17187
rect 31392 17144 31444 17153
rect 32128 17144 32180 17196
rect 34428 17187 34480 17196
rect 34428 17153 34437 17187
rect 34437 17153 34471 17187
rect 34471 17153 34480 17187
rect 34428 17144 34480 17153
rect 34612 17187 34664 17196
rect 34612 17153 34621 17187
rect 34621 17153 34655 17187
rect 34655 17153 34664 17187
rect 34612 17144 34664 17153
rect 35992 17212 36044 17264
rect 37096 17212 37148 17264
rect 36728 17144 36780 17196
rect 37372 17144 37424 17196
rect 38752 17212 38804 17264
rect 41512 17212 41564 17264
rect 41696 17212 41748 17264
rect 38384 17144 38436 17196
rect 38936 17187 38988 17196
rect 38936 17153 38945 17187
rect 38945 17153 38979 17187
rect 38979 17153 38988 17187
rect 38936 17144 38988 17153
rect 40040 17144 40092 17196
rect 40132 17187 40184 17196
rect 40132 17153 40153 17187
rect 40153 17153 40184 17187
rect 40132 17144 40184 17153
rect 27160 17119 27212 17128
rect 27160 17085 27169 17119
rect 27169 17085 27203 17119
rect 27203 17085 27212 17119
rect 27160 17076 27212 17085
rect 28724 17076 28776 17128
rect 25044 17008 25096 17060
rect 29552 17076 29604 17128
rect 34336 17076 34388 17128
rect 36912 17076 36964 17128
rect 22192 16940 22244 16992
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 23388 16940 23440 16949
rect 26516 16940 26568 16992
rect 28632 16940 28684 16992
rect 31944 17008 31996 17060
rect 37464 17051 37516 17060
rect 37464 17017 37473 17051
rect 37473 17017 37507 17051
rect 37507 17017 37516 17051
rect 37464 17008 37516 17017
rect 29184 16940 29236 16992
rect 31024 16940 31076 16992
rect 34612 16940 34664 16992
rect 37556 16940 37608 16992
rect 38844 17119 38896 17128
rect 38844 17085 38853 17119
rect 38853 17085 38887 17119
rect 38887 17085 38896 17119
rect 38844 17076 38896 17085
rect 39120 17076 39172 17128
rect 42248 17144 42300 17196
rect 43996 17144 44048 17196
rect 39948 17051 40000 17060
rect 39948 17017 39957 17051
rect 39957 17017 39991 17051
rect 39991 17017 40000 17051
rect 39948 17008 40000 17017
rect 43536 17076 43588 17128
rect 38292 16940 38344 16992
rect 38476 16940 38528 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 14740 16668 14792 16720
rect 15200 16600 15252 16652
rect 15476 16600 15528 16652
rect 17960 16668 18012 16720
rect 19248 16668 19300 16720
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 19064 16600 19116 16652
rect 20168 16668 20220 16720
rect 14924 16532 14976 16584
rect 15568 16532 15620 16584
rect 18236 16532 18288 16584
rect 18604 16532 18656 16584
rect 20536 16600 20588 16652
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 22192 16779 22244 16788
rect 22192 16745 22201 16779
rect 22201 16745 22235 16779
rect 22235 16745 22244 16779
rect 22192 16736 22244 16745
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 21640 16711 21692 16720
rect 21640 16677 21649 16711
rect 21649 16677 21683 16711
rect 21683 16677 21692 16711
rect 21640 16668 21692 16677
rect 27436 16736 27488 16788
rect 27804 16736 27856 16788
rect 29000 16736 29052 16788
rect 30196 16779 30248 16788
rect 30196 16745 30205 16779
rect 30205 16745 30239 16779
rect 30239 16745 30248 16779
rect 30196 16736 30248 16745
rect 30380 16736 30432 16788
rect 23388 16532 23440 16584
rect 25136 16532 25188 16584
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 27620 16532 27672 16584
rect 28540 16600 28592 16652
rect 30656 16668 30708 16720
rect 32404 16779 32456 16788
rect 32404 16745 32413 16779
rect 32413 16745 32447 16779
rect 32447 16745 32456 16779
rect 32404 16736 32456 16745
rect 33416 16736 33468 16788
rect 29092 16600 29144 16652
rect 28632 16532 28684 16584
rect 16948 16464 17000 16516
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 17040 16396 17092 16448
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 22376 16464 22428 16516
rect 28908 16575 28960 16584
rect 28908 16541 28917 16575
rect 28917 16541 28951 16575
rect 28951 16541 28960 16575
rect 32496 16600 32548 16652
rect 35072 16736 35124 16788
rect 35532 16736 35584 16788
rect 36268 16779 36320 16788
rect 36268 16745 36277 16779
rect 36277 16745 36311 16779
rect 36311 16745 36320 16779
rect 36268 16736 36320 16745
rect 37740 16736 37792 16788
rect 37832 16736 37884 16788
rect 38384 16736 38436 16788
rect 39856 16736 39908 16788
rect 37188 16668 37240 16720
rect 34980 16643 35032 16652
rect 34980 16609 34989 16643
rect 34989 16609 35023 16643
rect 35023 16609 35032 16643
rect 34980 16600 35032 16609
rect 28908 16532 28960 16541
rect 32312 16532 32364 16584
rect 26976 16396 27028 16448
rect 29184 16464 29236 16516
rect 30656 16464 30708 16516
rect 31300 16464 31352 16516
rect 28816 16396 28868 16448
rect 30012 16396 30064 16448
rect 31484 16396 31536 16448
rect 31944 16507 31996 16516
rect 31944 16473 31953 16507
rect 31953 16473 31987 16507
rect 31987 16473 31996 16507
rect 31944 16464 31996 16473
rect 32864 16464 32916 16516
rect 33784 16464 33836 16516
rect 34336 16532 34388 16584
rect 37372 16600 37424 16652
rect 38476 16600 38528 16652
rect 35164 16575 35216 16584
rect 35164 16541 35173 16575
rect 35173 16541 35207 16575
rect 35207 16541 35216 16575
rect 35164 16532 35216 16541
rect 35256 16532 35308 16584
rect 34888 16507 34940 16516
rect 34888 16473 34897 16507
rect 34897 16473 34931 16507
rect 34931 16473 34940 16507
rect 34888 16464 34940 16473
rect 37188 16575 37240 16584
rect 37188 16541 37197 16575
rect 37197 16541 37231 16575
rect 37231 16541 37240 16575
rect 37188 16532 37240 16541
rect 37280 16575 37332 16584
rect 37280 16541 37289 16575
rect 37289 16541 37323 16575
rect 37323 16541 37332 16575
rect 37280 16532 37332 16541
rect 38108 16575 38160 16584
rect 38108 16541 38117 16575
rect 38117 16541 38151 16575
rect 38151 16541 38160 16575
rect 38108 16532 38160 16541
rect 38752 16532 38804 16584
rect 39212 16575 39264 16584
rect 39212 16541 39221 16575
rect 39221 16541 39255 16575
rect 39255 16541 39264 16575
rect 39212 16532 39264 16541
rect 41696 16643 41748 16652
rect 41696 16609 41705 16643
rect 41705 16609 41739 16643
rect 41739 16609 41748 16643
rect 41696 16600 41748 16609
rect 40224 16532 40276 16584
rect 40316 16532 40368 16584
rect 42892 16600 42944 16652
rect 42984 16532 43036 16584
rect 34428 16396 34480 16448
rect 35348 16439 35400 16448
rect 35348 16405 35357 16439
rect 35357 16405 35391 16439
rect 35391 16405 35400 16439
rect 35348 16396 35400 16405
rect 35624 16396 35676 16448
rect 35992 16396 36044 16448
rect 36452 16464 36504 16516
rect 37648 16464 37700 16516
rect 38016 16464 38068 16516
rect 36820 16396 36872 16448
rect 37924 16396 37976 16448
rect 41512 16464 41564 16516
rect 41052 16439 41104 16448
rect 41052 16405 41061 16439
rect 41061 16405 41095 16439
rect 41095 16405 41104 16439
rect 41052 16396 41104 16405
rect 42800 16396 42852 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 14648 16235 14700 16244
rect 14648 16201 14657 16235
rect 14657 16201 14691 16235
rect 14691 16201 14700 16235
rect 14648 16192 14700 16201
rect 15568 16235 15620 16244
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 17316 16192 17368 16244
rect 18144 16192 18196 16244
rect 19432 16192 19484 16244
rect 21456 16192 21508 16244
rect 22192 16192 22244 16244
rect 22744 16192 22796 16244
rect 26608 16235 26660 16244
rect 26608 16201 26617 16235
rect 26617 16201 26651 16235
rect 26651 16201 26660 16235
rect 26608 16192 26660 16201
rect 27620 16235 27672 16244
rect 27620 16201 27629 16235
rect 27629 16201 27663 16235
rect 27663 16201 27672 16235
rect 27620 16192 27672 16201
rect 12992 16124 13044 16176
rect 15752 16124 15804 16176
rect 16948 16167 17000 16176
rect 16948 16133 16957 16167
rect 16957 16133 16991 16167
rect 16991 16133 17000 16167
rect 16948 16124 17000 16133
rect 18512 16167 18564 16176
rect 18512 16133 18530 16167
rect 18530 16133 18564 16167
rect 18512 16124 18564 16133
rect 22652 16124 22704 16176
rect 34980 16192 35032 16244
rect 36728 16192 36780 16244
rect 37188 16192 37240 16244
rect 38660 16235 38712 16244
rect 38660 16201 38669 16235
rect 38669 16201 38703 16235
rect 38703 16201 38712 16235
rect 38660 16192 38712 16201
rect 40960 16192 41012 16244
rect 13360 16056 13412 16108
rect 15108 16056 15160 16108
rect 17684 16056 17736 16108
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 19156 16056 19208 16108
rect 19340 16056 19392 16108
rect 22376 16056 22428 16108
rect 23388 16056 23440 16108
rect 27804 16099 27856 16108
rect 27804 16065 27813 16099
rect 27813 16065 27847 16099
rect 27847 16065 27856 16099
rect 27804 16056 27856 16065
rect 34612 16167 34664 16176
rect 34612 16133 34621 16167
rect 34621 16133 34655 16167
rect 34655 16133 34664 16167
rect 34612 16124 34664 16133
rect 36176 16167 36228 16176
rect 36176 16133 36185 16167
rect 36185 16133 36219 16167
rect 36219 16133 36228 16167
rect 36176 16124 36228 16133
rect 39212 16124 39264 16176
rect 43168 16124 43220 16176
rect 29184 16056 29236 16108
rect 30104 16056 30156 16108
rect 21272 16031 21324 16040
rect 21272 15997 21281 16031
rect 21281 15997 21315 16031
rect 21315 15997 21324 16031
rect 21272 15988 21324 15997
rect 19340 15920 19392 15972
rect 21640 15920 21692 15972
rect 25136 15988 25188 16040
rect 27252 15988 27304 16040
rect 20260 15852 20312 15904
rect 22008 15895 22060 15904
rect 22008 15861 22017 15895
rect 22017 15861 22051 15895
rect 22051 15861 22060 15895
rect 22008 15852 22060 15861
rect 23664 15852 23716 15904
rect 28080 15895 28132 15904
rect 28080 15861 28089 15895
rect 28089 15861 28123 15895
rect 28123 15861 28132 15895
rect 28080 15852 28132 15861
rect 29552 16031 29604 16040
rect 29552 15997 29561 16031
rect 29561 15997 29595 16031
rect 29595 15997 29604 16031
rect 29552 15988 29604 15997
rect 31668 16056 31720 16108
rect 31576 15920 31628 15972
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 33232 16056 33284 16108
rect 33416 16099 33468 16108
rect 33416 16065 33425 16099
rect 33425 16065 33459 16099
rect 33459 16065 33468 16099
rect 33416 16056 33468 16065
rect 33876 16056 33928 16108
rect 35992 16099 36044 16108
rect 35992 16065 36001 16099
rect 36001 16065 36035 16099
rect 36035 16065 36044 16099
rect 35992 16056 36044 16065
rect 38200 16099 38252 16108
rect 38200 16065 38209 16099
rect 38209 16065 38243 16099
rect 38243 16065 38252 16099
rect 38200 16056 38252 16065
rect 38384 16099 38436 16108
rect 38384 16065 38393 16099
rect 38393 16065 38427 16099
rect 38427 16065 38436 16099
rect 38384 16056 38436 16065
rect 38476 16099 38528 16108
rect 38476 16065 38485 16099
rect 38485 16065 38519 16099
rect 38519 16065 38528 16099
rect 38476 16056 38528 16065
rect 39304 16099 39356 16108
rect 39304 16065 39313 16099
rect 39313 16065 39347 16099
rect 39347 16065 39356 16099
rect 39304 16056 39356 16065
rect 41236 16056 41288 16108
rect 31944 15988 31996 16040
rect 34336 15988 34388 16040
rect 35900 15988 35952 16040
rect 39856 15988 39908 16040
rect 33232 15920 33284 15972
rect 31392 15895 31444 15904
rect 31392 15861 31401 15895
rect 31401 15861 31435 15895
rect 31435 15861 31444 15895
rect 31392 15852 31444 15861
rect 32772 15852 32824 15904
rect 33140 15895 33192 15904
rect 33140 15861 33149 15895
rect 33149 15861 33183 15895
rect 33183 15861 33192 15895
rect 33140 15852 33192 15861
rect 34796 15920 34848 15972
rect 34980 15920 35032 15972
rect 36728 15920 36780 15972
rect 37280 15920 37332 15972
rect 37924 15920 37976 15972
rect 34612 15895 34664 15904
rect 34612 15861 34621 15895
rect 34621 15861 34655 15895
rect 34655 15861 34664 15895
rect 34612 15852 34664 15861
rect 35164 15852 35216 15904
rect 37188 15852 37240 15904
rect 39028 15852 39080 15904
rect 40224 15852 40276 15904
rect 42984 15920 43036 15972
rect 41328 15852 41380 15904
rect 41604 15852 41656 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17316 15648 17368 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 22192 15691 22244 15700
rect 22192 15657 22201 15691
rect 22201 15657 22235 15691
rect 22235 15657 22244 15691
rect 22192 15648 22244 15657
rect 23388 15691 23440 15700
rect 23388 15657 23397 15691
rect 23397 15657 23431 15691
rect 23431 15657 23440 15691
rect 23388 15648 23440 15657
rect 27252 15648 27304 15700
rect 27896 15648 27948 15700
rect 30104 15691 30156 15700
rect 30104 15657 30113 15691
rect 30113 15657 30147 15691
rect 30147 15657 30156 15691
rect 30104 15648 30156 15657
rect 31484 15648 31536 15700
rect 31760 15691 31812 15700
rect 31760 15657 31769 15691
rect 31769 15657 31803 15691
rect 31803 15657 31812 15691
rect 31760 15648 31812 15657
rect 16212 15512 16264 15564
rect 19064 15512 19116 15564
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 15660 15444 15712 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 18144 15444 18196 15496
rect 20260 15512 20312 15564
rect 20720 15512 20772 15564
rect 22376 15512 22428 15564
rect 25688 15512 25740 15564
rect 26240 15580 26292 15632
rect 30012 15580 30064 15632
rect 32864 15648 32916 15700
rect 28080 15512 28132 15564
rect 29920 15512 29972 15564
rect 31392 15512 31444 15564
rect 33140 15580 33192 15632
rect 32772 15555 32824 15564
rect 32772 15521 32781 15555
rect 32781 15521 32815 15555
rect 32815 15521 32824 15555
rect 32772 15512 32824 15521
rect 32864 15555 32916 15564
rect 32864 15521 32873 15555
rect 32873 15521 32907 15555
rect 32907 15521 32916 15555
rect 32864 15512 32916 15521
rect 22008 15444 22060 15496
rect 22836 15444 22888 15496
rect 28540 15444 28592 15496
rect 28908 15444 28960 15496
rect 30288 15487 30340 15496
rect 30288 15453 30297 15487
rect 30297 15453 30331 15487
rect 30331 15453 30340 15487
rect 30288 15444 30340 15453
rect 15292 15376 15344 15428
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17960 15308 18012 15360
rect 20076 15308 20128 15360
rect 22652 15376 22704 15428
rect 31116 15444 31168 15496
rect 31760 15444 31812 15496
rect 33508 15487 33560 15496
rect 33508 15453 33517 15487
rect 33517 15453 33551 15487
rect 33551 15453 33560 15487
rect 33508 15444 33560 15453
rect 35900 15648 35952 15700
rect 36636 15648 36688 15700
rect 38200 15691 38252 15700
rect 38200 15657 38209 15691
rect 38209 15657 38243 15691
rect 38243 15657 38252 15691
rect 38200 15648 38252 15657
rect 42892 15648 42944 15700
rect 38936 15623 38988 15632
rect 34244 15444 34296 15496
rect 34520 15444 34572 15496
rect 34704 15444 34756 15496
rect 35348 15512 35400 15564
rect 34796 15376 34848 15428
rect 35532 15444 35584 15496
rect 36268 15512 36320 15564
rect 37188 15512 37240 15564
rect 36636 15487 36688 15496
rect 36636 15453 36645 15487
rect 36645 15453 36679 15487
rect 36679 15453 36688 15487
rect 36636 15444 36688 15453
rect 36820 15487 36872 15496
rect 36820 15453 36829 15487
rect 36829 15453 36863 15487
rect 36863 15453 36872 15487
rect 36820 15444 36872 15453
rect 38936 15589 38945 15623
rect 38945 15589 38979 15623
rect 38979 15589 38988 15623
rect 38936 15580 38988 15589
rect 38384 15512 38436 15564
rect 40960 15555 41012 15564
rect 40960 15521 40969 15555
rect 40969 15521 41003 15555
rect 41003 15521 41012 15555
rect 40960 15512 41012 15521
rect 41144 15555 41196 15564
rect 41144 15521 41153 15555
rect 41153 15521 41187 15555
rect 41187 15521 41196 15555
rect 41144 15512 41196 15521
rect 41696 15512 41748 15564
rect 41972 15555 42024 15564
rect 41972 15521 41981 15555
rect 41981 15521 42015 15555
rect 42015 15521 42024 15555
rect 41972 15512 42024 15521
rect 37924 15487 37976 15496
rect 37924 15453 37933 15487
rect 37933 15453 37967 15487
rect 37967 15453 37976 15487
rect 37924 15444 37976 15453
rect 35624 15376 35676 15428
rect 36084 15376 36136 15428
rect 39212 15487 39264 15496
rect 39212 15453 39221 15487
rect 39221 15453 39255 15487
rect 39255 15453 39264 15487
rect 39212 15444 39264 15453
rect 41328 15444 41380 15496
rect 25228 15308 25280 15360
rect 26056 15308 26108 15360
rect 27620 15308 27672 15360
rect 27988 15308 28040 15360
rect 32404 15308 32456 15360
rect 34152 15351 34204 15360
rect 34152 15317 34161 15351
rect 34161 15317 34195 15351
rect 34195 15317 34204 15351
rect 34152 15308 34204 15317
rect 40500 15351 40552 15360
rect 40500 15317 40509 15351
rect 40509 15317 40543 15351
rect 40543 15317 40552 15351
rect 40500 15308 40552 15317
rect 43168 15444 43220 15496
rect 42616 15376 42668 15428
rect 41052 15308 41104 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 14832 15147 14884 15156
rect 14832 15113 14841 15147
rect 14841 15113 14875 15147
rect 14875 15113 14884 15147
rect 14832 15104 14884 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 18052 15104 18104 15156
rect 19984 15104 20036 15156
rect 21456 15104 21508 15156
rect 22836 15104 22888 15156
rect 26056 15147 26108 15156
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 28724 15104 28776 15156
rect 29092 15104 29144 15156
rect 31760 15104 31812 15156
rect 35440 15104 35492 15156
rect 36820 15104 36872 15156
rect 37096 15104 37148 15156
rect 15108 15036 15160 15088
rect 13360 14968 13412 15020
rect 14280 14968 14332 15020
rect 14832 14968 14884 15020
rect 17132 15011 17184 15020
rect 17132 14977 17166 15011
rect 17166 14977 17184 15011
rect 17132 14968 17184 14977
rect 19156 14968 19208 15020
rect 20720 15036 20772 15088
rect 23664 15079 23716 15088
rect 23664 15045 23682 15079
rect 23682 15045 23716 15079
rect 23664 15036 23716 15045
rect 27344 15036 27396 15088
rect 29276 15036 29328 15088
rect 32772 15036 32824 15088
rect 33324 15079 33376 15088
rect 33324 15045 33333 15079
rect 33333 15045 33367 15079
rect 33367 15045 33376 15079
rect 33324 15036 33376 15045
rect 34704 15079 34756 15088
rect 34704 15045 34721 15079
rect 34721 15045 34756 15079
rect 34704 15036 34756 15045
rect 20076 14968 20128 15020
rect 24952 15011 25004 15020
rect 24952 14977 24986 15011
rect 24986 14977 25004 15011
rect 24952 14968 25004 14977
rect 27620 14968 27672 15020
rect 15016 14900 15068 14952
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 15476 14764 15528 14816
rect 19340 14832 19392 14884
rect 19432 14764 19484 14816
rect 23940 14943 23992 14952
rect 23940 14909 23949 14943
rect 23949 14909 23983 14943
rect 23983 14909 23992 14943
rect 23940 14900 23992 14909
rect 29000 15011 29052 15020
rect 29000 14977 29009 15011
rect 29009 14977 29043 15011
rect 29043 14977 29052 15011
rect 29000 14968 29052 14977
rect 29184 14968 29236 15020
rect 31484 14968 31536 15020
rect 33232 14968 33284 15020
rect 35072 15036 35124 15088
rect 35900 15036 35952 15088
rect 37924 15036 37976 15088
rect 34888 15011 34940 15020
rect 34888 14977 34897 15011
rect 34897 14977 34931 15011
rect 34931 14977 34940 15011
rect 34888 14968 34940 14977
rect 29092 14900 29144 14952
rect 34520 14943 34572 14952
rect 34520 14909 34529 14943
rect 34529 14909 34563 14943
rect 34563 14909 34572 14943
rect 34520 14900 34572 14909
rect 34612 14832 34664 14884
rect 36360 14968 36412 15020
rect 36452 15011 36504 15020
rect 36452 14977 36461 15011
rect 36461 14977 36495 15011
rect 36495 14977 36504 15011
rect 36452 14968 36504 14977
rect 36728 15011 36780 15020
rect 36728 14977 36737 15011
rect 36737 14977 36771 15011
rect 36771 14977 36780 15011
rect 36728 14968 36780 14977
rect 35532 14832 35584 14884
rect 37280 14900 37332 14952
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 37648 15011 37700 15020
rect 37648 14977 37657 15011
rect 37657 14977 37691 15011
rect 37691 14977 37700 15011
rect 37648 14968 37700 14977
rect 38384 15104 38436 15156
rect 41236 15104 41288 15156
rect 41880 15104 41932 15156
rect 42616 15147 42668 15156
rect 42616 15113 42625 15147
rect 42625 15113 42659 15147
rect 42659 15113 42668 15147
rect 42616 15104 42668 15113
rect 43352 15147 43404 15156
rect 43352 15113 43361 15147
rect 43361 15113 43395 15147
rect 43395 15113 43404 15147
rect 43352 15104 43404 15113
rect 38108 15036 38160 15088
rect 38752 15036 38804 15088
rect 40132 15036 40184 15088
rect 39764 15011 39816 15020
rect 39764 14977 39773 15011
rect 39773 14977 39807 15011
rect 39807 14977 39816 15011
rect 39764 14968 39816 14977
rect 41052 14968 41104 15020
rect 41604 14968 41656 15020
rect 42800 15011 42852 15020
rect 42800 14977 42809 15011
rect 42809 14977 42843 15011
rect 42843 14977 42852 15011
rect 42800 14968 42852 14977
rect 39856 14900 39908 14952
rect 36728 14832 36780 14884
rect 20168 14764 20220 14816
rect 27528 14807 27580 14816
rect 27528 14773 27537 14807
rect 27537 14773 27571 14807
rect 27571 14773 27580 14807
rect 27528 14764 27580 14773
rect 28724 14764 28776 14816
rect 29092 14764 29144 14816
rect 29736 14807 29788 14816
rect 29736 14773 29745 14807
rect 29745 14773 29779 14807
rect 29779 14773 29788 14807
rect 29736 14764 29788 14773
rect 30288 14764 30340 14816
rect 33416 14764 33468 14816
rect 33784 14764 33836 14816
rect 36268 14764 36320 14816
rect 36452 14807 36504 14816
rect 36452 14773 36461 14807
rect 36461 14773 36495 14807
rect 36495 14773 36504 14807
rect 39028 14832 39080 14884
rect 36452 14764 36504 14773
rect 37832 14764 37884 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 16948 14560 17000 14612
rect 15936 14492 15988 14544
rect 20076 14560 20128 14612
rect 20352 14560 20404 14612
rect 20812 14603 20864 14612
rect 20812 14569 20821 14603
rect 20821 14569 20855 14603
rect 20855 14569 20864 14603
rect 20812 14560 20864 14569
rect 22376 14603 22428 14612
rect 22376 14569 22385 14603
rect 22385 14569 22419 14603
rect 22419 14569 22428 14603
rect 22376 14560 22428 14569
rect 24952 14560 25004 14612
rect 27436 14560 27488 14612
rect 27712 14560 27764 14612
rect 29184 14603 29236 14612
rect 29184 14569 29193 14603
rect 29193 14569 29227 14603
rect 29227 14569 29236 14603
rect 29184 14560 29236 14569
rect 29736 14603 29788 14612
rect 29736 14569 29745 14603
rect 29745 14569 29779 14603
rect 29779 14569 29788 14603
rect 29736 14560 29788 14569
rect 30012 14560 30064 14612
rect 28908 14492 28960 14544
rect 29000 14492 29052 14544
rect 31300 14492 31352 14544
rect 34520 14560 34572 14612
rect 35072 14603 35124 14612
rect 35072 14569 35081 14603
rect 35081 14569 35115 14603
rect 35115 14569 35124 14603
rect 35072 14560 35124 14569
rect 36544 14560 36596 14612
rect 38108 14560 38160 14612
rect 40132 14560 40184 14612
rect 40224 14560 40276 14612
rect 41788 14603 41840 14612
rect 41788 14569 41797 14603
rect 41797 14569 41831 14603
rect 41831 14569 41840 14603
rect 41788 14560 41840 14569
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 15752 14424 15804 14476
rect 16212 14424 16264 14476
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 17684 14467 17736 14476
rect 17684 14433 17693 14467
rect 17693 14433 17727 14467
rect 17727 14433 17736 14467
rect 17684 14424 17736 14433
rect 19156 14424 19208 14476
rect 23940 14424 23992 14476
rect 25136 14424 25188 14476
rect 15844 14356 15896 14408
rect 18052 14356 18104 14408
rect 20260 14356 20312 14408
rect 25228 14399 25280 14408
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 29828 14424 29880 14476
rect 28816 14399 28868 14408
rect 28816 14365 28825 14399
rect 28825 14365 28859 14399
rect 28859 14365 28868 14399
rect 28816 14356 28868 14365
rect 30564 14424 30616 14476
rect 31668 14467 31720 14476
rect 31668 14433 31678 14467
rect 31678 14433 31712 14467
rect 31712 14433 31720 14467
rect 31668 14424 31720 14433
rect 31760 14467 31812 14476
rect 31760 14433 31769 14467
rect 31769 14433 31803 14467
rect 31803 14433 31812 14467
rect 31760 14424 31812 14433
rect 35900 14492 35952 14544
rect 32588 14424 32640 14476
rect 14832 14220 14884 14272
rect 26792 14288 26844 14340
rect 28632 14288 28684 14340
rect 30104 14399 30156 14408
rect 30104 14365 30113 14399
rect 30113 14365 30147 14399
rect 30147 14365 30156 14399
rect 30104 14356 30156 14365
rect 30932 14356 30984 14408
rect 30472 14288 30524 14340
rect 32496 14399 32548 14408
rect 32496 14365 32505 14399
rect 32505 14365 32539 14399
rect 32539 14365 32548 14399
rect 32496 14356 32548 14365
rect 32772 14356 32824 14408
rect 33508 14356 33560 14408
rect 33048 14288 33100 14340
rect 35808 14356 35860 14408
rect 36360 14467 36412 14476
rect 36360 14433 36369 14467
rect 36369 14433 36403 14467
rect 36403 14433 36412 14467
rect 36360 14424 36412 14433
rect 38108 14424 38160 14476
rect 38200 14424 38252 14476
rect 39764 14424 39816 14476
rect 39856 14424 39908 14476
rect 33876 14331 33928 14340
rect 33876 14297 33885 14331
rect 33885 14297 33919 14331
rect 33919 14297 33928 14331
rect 33876 14288 33928 14297
rect 35348 14288 35400 14340
rect 24400 14220 24452 14272
rect 25228 14220 25280 14272
rect 30748 14263 30800 14272
rect 30748 14229 30757 14263
rect 30757 14229 30791 14263
rect 30791 14229 30800 14263
rect 30748 14220 30800 14229
rect 31484 14263 31536 14272
rect 31484 14229 31493 14263
rect 31493 14229 31527 14263
rect 31527 14229 31536 14263
rect 31484 14220 31536 14229
rect 31576 14220 31628 14272
rect 33784 14220 33836 14272
rect 35164 14220 35216 14272
rect 35808 14220 35860 14272
rect 36820 14331 36872 14340
rect 36820 14297 36829 14331
rect 36829 14297 36863 14331
rect 36863 14297 36872 14331
rect 36820 14288 36872 14297
rect 36176 14220 36228 14272
rect 37188 14399 37240 14408
rect 37188 14365 37197 14399
rect 37197 14365 37231 14399
rect 37231 14365 37240 14399
rect 37188 14356 37240 14365
rect 37556 14356 37608 14408
rect 37740 14399 37792 14408
rect 37740 14365 37749 14399
rect 37749 14365 37783 14399
rect 37783 14365 37792 14399
rect 37740 14356 37792 14365
rect 38292 14288 38344 14340
rect 39120 14356 39172 14408
rect 39580 14356 39632 14408
rect 40132 14356 40184 14408
rect 43352 14399 43404 14408
rect 43352 14365 43361 14399
rect 43361 14365 43395 14399
rect 43395 14365 43404 14399
rect 43352 14356 43404 14365
rect 40316 14288 40368 14340
rect 40592 14288 40644 14340
rect 43076 14331 43128 14340
rect 43076 14297 43085 14331
rect 43085 14297 43119 14331
rect 43119 14297 43128 14331
rect 43076 14288 43128 14297
rect 37924 14263 37976 14272
rect 37924 14229 37933 14263
rect 37933 14229 37967 14263
rect 37967 14229 37976 14263
rect 37924 14220 37976 14229
rect 38568 14220 38620 14272
rect 40500 14220 40552 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 15844 14016 15896 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 17500 14016 17552 14068
rect 19984 14016 20036 14068
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 20812 14016 20864 14068
rect 23756 14016 23808 14068
rect 15108 13948 15160 14000
rect 14464 13923 14516 13932
rect 14464 13889 14498 13923
rect 14498 13889 14516 13923
rect 14464 13880 14516 13889
rect 19156 13948 19208 14000
rect 20168 13948 20220 14000
rect 22192 13948 22244 14000
rect 22468 13948 22520 14000
rect 19524 13880 19576 13932
rect 25228 14059 25280 14068
rect 25228 14025 25237 14059
rect 25237 14025 25271 14059
rect 25271 14025 25280 14059
rect 25228 14016 25280 14025
rect 27344 14016 27396 14068
rect 30012 14016 30064 14068
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 30472 14059 30524 14068
rect 30472 14025 30481 14059
rect 30481 14025 30515 14059
rect 30515 14025 30524 14059
rect 30472 14016 30524 14025
rect 31484 14016 31536 14068
rect 31576 14059 31628 14068
rect 31576 14025 31585 14059
rect 31585 14025 31619 14059
rect 31619 14025 31628 14059
rect 31576 14016 31628 14025
rect 27528 13948 27580 14000
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 29000 13880 29052 13932
rect 29092 13923 29144 13932
rect 29092 13889 29101 13923
rect 29101 13889 29135 13923
rect 29135 13889 29144 13923
rect 29092 13880 29144 13889
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 29644 13948 29696 14000
rect 29736 13948 29788 14000
rect 34152 14016 34204 14068
rect 34428 14016 34480 14068
rect 20168 13744 20220 13796
rect 22376 13744 22428 13796
rect 24860 13812 24912 13864
rect 29184 13812 29236 13864
rect 30288 13923 30340 13932
rect 30288 13889 30297 13923
rect 30297 13889 30331 13923
rect 30331 13889 30340 13923
rect 30288 13880 30340 13889
rect 30380 13880 30432 13932
rect 31760 13991 31812 14000
rect 31760 13957 31769 13991
rect 31769 13957 31803 13991
rect 31803 13957 31812 13991
rect 31760 13948 31812 13957
rect 33048 13948 33100 14000
rect 33416 13991 33468 14000
rect 33416 13957 33425 13991
rect 33425 13957 33459 13991
rect 33459 13957 33468 13991
rect 33416 13948 33468 13957
rect 33508 13948 33560 14000
rect 36084 14016 36136 14068
rect 37096 14016 37148 14068
rect 37372 14016 37424 14068
rect 38292 14059 38344 14068
rect 38292 14025 38301 14059
rect 38301 14025 38335 14059
rect 38335 14025 38344 14059
rect 38292 14016 38344 14025
rect 41236 14016 41288 14068
rect 26240 13744 26292 13796
rect 30748 13812 30800 13864
rect 31668 13880 31720 13932
rect 34888 13923 34940 13932
rect 34888 13889 34897 13923
rect 34897 13889 34931 13923
rect 34931 13889 34940 13923
rect 34888 13880 34940 13889
rect 35624 13948 35676 14000
rect 35532 13923 35584 13932
rect 35532 13889 35535 13923
rect 35535 13889 35569 13923
rect 35569 13889 35584 13923
rect 35532 13880 35584 13889
rect 32772 13812 32824 13864
rect 34704 13812 34756 13864
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 26516 13719 26568 13728
rect 26516 13685 26525 13719
rect 26525 13685 26559 13719
rect 26559 13685 26568 13719
rect 26516 13676 26568 13685
rect 27620 13676 27672 13728
rect 34888 13744 34940 13796
rect 35624 13744 35676 13796
rect 36360 13880 36412 13932
rect 36728 13812 36780 13864
rect 37464 13923 37516 13932
rect 37464 13889 37473 13923
rect 37473 13889 37507 13923
rect 37507 13889 37516 13923
rect 37464 13880 37516 13889
rect 38660 13948 38712 14000
rect 39120 13948 39172 14000
rect 43076 14016 43128 14068
rect 41880 13948 41932 14000
rect 37740 13812 37792 13864
rect 38568 13812 38620 13864
rect 39028 13923 39080 13932
rect 39028 13889 39037 13923
rect 39037 13889 39071 13923
rect 39071 13889 39080 13923
rect 39028 13880 39080 13889
rect 39580 13923 39632 13932
rect 39580 13889 39589 13923
rect 39589 13889 39623 13923
rect 39623 13889 39632 13923
rect 39580 13880 39632 13889
rect 39764 13880 39816 13932
rect 40500 13880 40552 13932
rect 41052 13812 41104 13864
rect 42892 13812 42944 13864
rect 43076 13855 43128 13864
rect 43076 13821 43085 13855
rect 43085 13821 43119 13855
rect 43119 13821 43128 13855
rect 43076 13812 43128 13821
rect 38752 13744 38804 13796
rect 40040 13744 40092 13796
rect 41144 13744 41196 13796
rect 43168 13744 43220 13796
rect 29184 13676 29236 13728
rect 29460 13676 29512 13728
rect 29552 13676 29604 13728
rect 32220 13676 32272 13728
rect 32496 13676 32548 13728
rect 33140 13676 33192 13728
rect 34704 13676 34756 13728
rect 35440 13676 35492 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14464 13472 14516 13524
rect 15476 13472 15528 13524
rect 19524 13472 19576 13524
rect 23756 13472 23808 13524
rect 25228 13472 25280 13524
rect 26792 13515 26844 13524
rect 26792 13481 26801 13515
rect 26801 13481 26835 13515
rect 26835 13481 26844 13515
rect 26792 13472 26844 13481
rect 29092 13472 29144 13524
rect 31852 13472 31904 13524
rect 34796 13472 34848 13524
rect 35716 13515 35768 13524
rect 35716 13481 35725 13515
rect 35725 13481 35759 13515
rect 35759 13481 35768 13515
rect 35716 13472 35768 13481
rect 37464 13515 37516 13524
rect 37464 13481 37473 13515
rect 37473 13481 37507 13515
rect 37507 13481 37516 13515
rect 37464 13472 37516 13481
rect 38660 13515 38712 13524
rect 38660 13481 38669 13515
rect 38669 13481 38703 13515
rect 38703 13481 38712 13515
rect 38660 13472 38712 13481
rect 43076 13472 43128 13524
rect 19340 13404 19392 13456
rect 29276 13404 29328 13456
rect 26516 13336 26568 13388
rect 27436 13379 27488 13388
rect 27436 13345 27445 13379
rect 27445 13345 27479 13379
rect 27479 13345 27488 13379
rect 27436 13336 27488 13345
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 19432 13268 19484 13320
rect 22008 13268 22060 13320
rect 23940 13268 23992 13320
rect 25136 13268 25188 13320
rect 29736 13336 29788 13388
rect 28908 13311 28960 13320
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 30840 13336 30892 13388
rect 31668 13336 31720 13388
rect 33140 13404 33192 13456
rect 33232 13404 33284 13456
rect 34244 13404 34296 13456
rect 35348 13404 35400 13456
rect 36452 13404 36504 13456
rect 40040 13404 40092 13456
rect 30012 13311 30064 13320
rect 30012 13277 30021 13311
rect 30021 13277 30055 13311
rect 30055 13277 30064 13311
rect 30012 13268 30064 13277
rect 30380 13268 30432 13320
rect 31024 13311 31076 13320
rect 31024 13277 31033 13311
rect 31033 13277 31067 13311
rect 31067 13277 31076 13311
rect 31024 13268 31076 13277
rect 21272 13132 21324 13184
rect 22192 13200 22244 13252
rect 22652 13200 22704 13252
rect 24860 13243 24912 13252
rect 24860 13209 24894 13243
rect 24894 13209 24912 13243
rect 24860 13200 24912 13209
rect 27620 13200 27672 13252
rect 31852 13268 31904 13320
rect 34428 13336 34480 13388
rect 23296 13132 23348 13184
rect 29920 13132 29972 13184
rect 31484 13200 31536 13252
rect 32220 13311 32272 13320
rect 32220 13277 32229 13311
rect 32229 13277 32263 13311
rect 32263 13277 32272 13311
rect 32220 13268 32272 13277
rect 30748 13175 30800 13184
rect 30748 13141 30757 13175
rect 30757 13141 30791 13175
rect 30791 13141 30800 13175
rect 30748 13132 30800 13141
rect 31024 13132 31076 13184
rect 33784 13268 33836 13320
rect 35532 13336 35584 13388
rect 35624 13268 35676 13320
rect 35808 13268 35860 13320
rect 34520 13200 34572 13252
rect 37372 13268 37424 13320
rect 37556 13268 37608 13320
rect 32956 13132 33008 13184
rect 37280 13243 37332 13252
rect 37280 13209 37289 13243
rect 37289 13209 37323 13243
rect 37323 13209 37332 13243
rect 38568 13311 38620 13320
rect 38568 13277 38577 13311
rect 38577 13277 38611 13311
rect 38611 13277 38620 13311
rect 38568 13268 38620 13277
rect 38752 13311 38804 13320
rect 38752 13277 38761 13311
rect 38761 13277 38795 13311
rect 38795 13277 38804 13311
rect 38752 13268 38804 13277
rect 41328 13268 41380 13320
rect 41972 13268 42024 13320
rect 37280 13200 37332 13209
rect 40408 13200 40460 13252
rect 42156 13243 42208 13252
rect 42156 13209 42190 13243
rect 42190 13209 42208 13243
rect 42156 13200 42208 13209
rect 41052 13132 41104 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 20168 12971 20220 12980
rect 20168 12937 20177 12971
rect 20177 12937 20211 12971
rect 20211 12937 20220 12971
rect 20168 12928 20220 12937
rect 23296 12928 23348 12980
rect 26240 12928 26292 12980
rect 26608 12928 26660 12980
rect 29644 12928 29696 12980
rect 31668 12971 31720 12980
rect 31668 12937 31677 12971
rect 31677 12937 31711 12971
rect 31711 12937 31720 12971
rect 31668 12928 31720 12937
rect 31760 12928 31812 12980
rect 31852 12928 31904 12980
rect 32404 12928 32456 12980
rect 32956 12971 33008 12980
rect 32956 12937 32965 12971
rect 32965 12937 32999 12971
rect 32999 12937 33008 12971
rect 32956 12928 33008 12937
rect 33324 12928 33376 12980
rect 29184 12860 29236 12912
rect 21272 12835 21324 12844
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 27344 12792 27396 12844
rect 29552 12835 29604 12844
rect 29552 12801 29570 12835
rect 29570 12801 29604 12835
rect 29552 12792 29604 12801
rect 30012 12792 30064 12844
rect 29828 12767 29880 12776
rect 29828 12733 29837 12767
rect 29837 12733 29871 12767
rect 29871 12733 29880 12767
rect 29828 12724 29880 12733
rect 30564 12724 30616 12776
rect 31024 12792 31076 12844
rect 31760 12835 31812 12844
rect 31760 12801 31769 12835
rect 31769 12801 31803 12835
rect 31803 12801 31812 12835
rect 31760 12792 31812 12801
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 35624 12903 35676 12912
rect 35624 12869 35633 12903
rect 35633 12869 35667 12903
rect 35667 12869 35676 12903
rect 35624 12860 35676 12869
rect 36820 12928 36872 12980
rect 38752 12928 38804 12980
rect 41052 12928 41104 12980
rect 41420 12971 41472 12980
rect 41420 12937 41429 12971
rect 41429 12937 41463 12971
rect 41463 12937 41472 12971
rect 41420 12928 41472 12937
rect 41880 12928 41932 12980
rect 42156 12928 42208 12980
rect 32864 12724 32916 12776
rect 34428 12835 34480 12844
rect 34428 12801 34437 12835
rect 34437 12801 34471 12835
rect 34471 12801 34480 12835
rect 34428 12792 34480 12801
rect 34888 12792 34940 12844
rect 35348 12792 35400 12844
rect 34612 12767 34664 12776
rect 34612 12733 34621 12767
rect 34621 12733 34655 12767
rect 34655 12733 34664 12767
rect 34612 12724 34664 12733
rect 35992 12724 36044 12776
rect 37464 12792 37516 12844
rect 38568 12792 38620 12844
rect 42524 12860 42576 12912
rect 41236 12792 41288 12844
rect 42984 12971 43036 12980
rect 42984 12937 42993 12971
rect 42993 12937 43027 12971
rect 43027 12937 43036 12971
rect 42984 12928 43036 12937
rect 43076 12971 43128 12980
rect 43076 12937 43085 12971
rect 43085 12937 43119 12971
rect 43119 12937 43128 12971
rect 43076 12928 43128 12937
rect 43352 12860 43404 12912
rect 38660 12767 38712 12776
rect 38660 12733 38669 12767
rect 38669 12733 38703 12767
rect 38703 12733 38712 12767
rect 38660 12724 38712 12733
rect 41052 12724 41104 12776
rect 42892 12724 42944 12776
rect 32772 12656 32824 12708
rect 34704 12656 34756 12708
rect 27436 12588 27488 12640
rect 30932 12588 30984 12640
rect 32128 12588 32180 12640
rect 34336 12588 34388 12640
rect 34796 12588 34848 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 26424 12427 26476 12436
rect 26424 12393 26433 12427
rect 26433 12393 26467 12427
rect 26467 12393 26476 12427
rect 26424 12384 26476 12393
rect 27344 12427 27396 12436
rect 27344 12393 27353 12427
rect 27353 12393 27387 12427
rect 27387 12393 27396 12427
rect 27344 12384 27396 12393
rect 30564 12384 30616 12436
rect 31116 12384 31168 12436
rect 32220 12427 32272 12436
rect 32220 12393 32229 12427
rect 32229 12393 32263 12427
rect 32263 12393 32272 12427
rect 32220 12384 32272 12393
rect 37096 12427 37148 12436
rect 37096 12393 37105 12427
rect 37105 12393 37139 12427
rect 37139 12393 37148 12427
rect 37096 12384 37148 12393
rect 38660 12427 38712 12436
rect 38660 12393 38669 12427
rect 38669 12393 38703 12427
rect 38703 12393 38712 12427
rect 38660 12384 38712 12393
rect 40592 12427 40644 12436
rect 40592 12393 40601 12427
rect 40601 12393 40635 12427
rect 40635 12393 40644 12427
rect 40592 12384 40644 12393
rect 41512 12427 41564 12436
rect 41512 12393 41521 12427
rect 41521 12393 41555 12427
rect 41555 12393 41564 12427
rect 41512 12384 41564 12393
rect 28908 12316 28960 12368
rect 29460 12316 29512 12368
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 26608 12248 26660 12300
rect 28816 12180 28868 12232
rect 25412 12087 25464 12096
rect 25412 12053 25421 12087
rect 25421 12053 25455 12087
rect 25455 12053 25464 12087
rect 25412 12044 25464 12053
rect 28448 12044 28500 12096
rect 30472 12248 30524 12300
rect 30656 12223 30708 12232
rect 30656 12189 30665 12223
rect 30665 12189 30699 12223
rect 30699 12189 30708 12223
rect 30656 12180 30708 12189
rect 31760 12316 31812 12368
rect 32128 12248 32180 12300
rect 32312 12291 32364 12300
rect 32312 12257 32321 12291
rect 32321 12257 32355 12291
rect 32355 12257 32364 12291
rect 32312 12248 32364 12257
rect 32864 12248 32916 12300
rect 34060 12291 34112 12300
rect 34060 12257 34069 12291
rect 34069 12257 34103 12291
rect 34103 12257 34112 12291
rect 34060 12248 34112 12257
rect 30932 12223 30984 12232
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 32220 12223 32272 12232
rect 32220 12189 32229 12223
rect 32229 12189 32263 12223
rect 32263 12189 32272 12223
rect 32220 12180 32272 12189
rect 34152 12223 34204 12232
rect 34152 12189 34161 12223
rect 34161 12189 34195 12223
rect 34195 12189 34204 12223
rect 34152 12180 34204 12189
rect 34336 12223 34388 12232
rect 34336 12189 34345 12223
rect 34345 12189 34379 12223
rect 34379 12189 34388 12223
rect 34336 12180 34388 12189
rect 36636 12248 36688 12300
rect 35532 12180 35584 12232
rect 37280 12155 37332 12164
rect 30012 12044 30064 12096
rect 30840 12044 30892 12096
rect 32036 12087 32088 12096
rect 32036 12053 32045 12087
rect 32045 12053 32079 12087
rect 32079 12053 32088 12087
rect 32036 12044 32088 12053
rect 32772 12044 32824 12096
rect 33876 12044 33928 12096
rect 34612 12044 34664 12096
rect 37280 12121 37289 12155
rect 37289 12121 37323 12155
rect 37323 12121 37332 12155
rect 37280 12112 37332 12121
rect 38292 12180 38344 12232
rect 39212 12316 39264 12368
rect 41972 12291 42024 12300
rect 41972 12257 41981 12291
rect 41981 12257 42015 12291
rect 42015 12257 42024 12291
rect 41972 12248 42024 12257
rect 38660 12180 38712 12232
rect 39396 12223 39448 12232
rect 39396 12189 39405 12223
rect 39405 12189 39439 12223
rect 39439 12189 39448 12223
rect 39396 12180 39448 12189
rect 42064 12112 42116 12164
rect 37648 12044 37700 12096
rect 43076 12044 43128 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 26148 11840 26200 11892
rect 28448 11840 28500 11892
rect 29460 11883 29512 11892
rect 29460 11849 29469 11883
rect 29469 11849 29503 11883
rect 29503 11849 29512 11883
rect 29460 11840 29512 11849
rect 30840 11883 30892 11892
rect 30840 11849 30849 11883
rect 30849 11849 30883 11883
rect 30883 11849 30892 11883
rect 30840 11840 30892 11849
rect 32220 11840 32272 11892
rect 32588 11883 32640 11892
rect 32588 11849 32597 11883
rect 32597 11849 32631 11883
rect 32631 11849 32640 11883
rect 32588 11840 32640 11849
rect 25412 11815 25464 11824
rect 25412 11781 25446 11815
rect 25446 11781 25464 11815
rect 25412 11772 25464 11781
rect 27436 11815 27488 11824
rect 27436 11781 27470 11815
rect 27470 11781 27488 11815
rect 27436 11772 27488 11781
rect 27528 11772 27580 11824
rect 32036 11772 32088 11824
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 29368 11747 29420 11756
rect 29368 11713 29377 11747
rect 29377 11713 29411 11747
rect 29411 11713 29420 11747
rect 29368 11704 29420 11713
rect 31760 11704 31812 11756
rect 32680 11704 32732 11756
rect 32772 11747 32824 11756
rect 32772 11713 32781 11747
rect 32781 11713 32815 11747
rect 32815 11713 32824 11747
rect 32772 11704 32824 11713
rect 34520 11840 34572 11892
rect 34980 11840 35032 11892
rect 35900 11840 35952 11892
rect 37372 11840 37424 11892
rect 39396 11840 39448 11892
rect 40868 11883 40920 11892
rect 40868 11849 40877 11883
rect 40877 11849 40911 11883
rect 40911 11849 40920 11883
rect 40868 11840 40920 11849
rect 42064 11883 42116 11892
rect 42064 11849 42073 11883
rect 42073 11849 42107 11883
rect 42107 11849 42116 11883
rect 42064 11840 42116 11849
rect 42616 11883 42668 11892
rect 42616 11849 42625 11883
rect 42625 11849 42659 11883
rect 42659 11849 42668 11883
rect 42616 11840 42668 11849
rect 43076 11883 43128 11892
rect 43076 11849 43085 11883
rect 43085 11849 43119 11883
rect 43119 11849 43128 11883
rect 43076 11840 43128 11849
rect 29184 11568 29236 11620
rect 30012 11636 30064 11688
rect 30564 11636 30616 11688
rect 30932 11679 30984 11688
rect 30932 11645 30941 11679
rect 30941 11645 30975 11679
rect 30975 11645 30984 11679
rect 30932 11636 30984 11645
rect 31024 11636 31076 11688
rect 34060 11704 34112 11756
rect 33324 11636 33376 11688
rect 34796 11747 34848 11756
rect 34796 11713 34805 11747
rect 34805 11713 34839 11747
rect 34839 11713 34848 11747
rect 34796 11704 34848 11713
rect 34980 11747 35032 11756
rect 34980 11713 34989 11747
rect 34989 11713 35023 11747
rect 35023 11713 35032 11747
rect 34980 11704 35032 11713
rect 37280 11772 37332 11824
rect 36176 11704 36228 11756
rect 37648 11747 37700 11756
rect 37648 11713 37657 11747
rect 37657 11713 37691 11747
rect 37691 11713 37700 11747
rect 37648 11704 37700 11713
rect 39672 11815 39724 11824
rect 39672 11781 39681 11815
rect 39681 11781 39715 11815
rect 39715 11781 39724 11815
rect 39672 11772 39724 11781
rect 40040 11772 40092 11824
rect 38660 11747 38712 11756
rect 38660 11713 38669 11747
rect 38669 11713 38703 11747
rect 38703 11713 38712 11747
rect 38660 11704 38712 11713
rect 40132 11704 40184 11756
rect 41144 11704 41196 11756
rect 42340 11704 42392 11756
rect 42984 11747 43036 11756
rect 42984 11713 42993 11747
rect 42993 11713 43027 11747
rect 43027 11713 43036 11747
rect 42984 11704 43036 11713
rect 41052 11679 41104 11688
rect 41052 11645 41061 11679
rect 41061 11645 41095 11679
rect 41095 11645 41104 11679
rect 41052 11636 41104 11645
rect 43168 11679 43220 11688
rect 43168 11645 43177 11679
rect 43177 11645 43211 11679
rect 43211 11645 43220 11679
rect 43168 11636 43220 11645
rect 34980 11568 35032 11620
rect 29000 11543 29052 11552
rect 29000 11509 29009 11543
rect 29009 11509 29043 11543
rect 29043 11509 29052 11543
rect 29000 11500 29052 11509
rect 30380 11543 30432 11552
rect 30380 11509 30389 11543
rect 30389 11509 30423 11543
rect 30423 11509 30432 11543
rect 30380 11500 30432 11509
rect 34428 11543 34480 11552
rect 34428 11509 34437 11543
rect 34437 11509 34471 11543
rect 34471 11509 34480 11543
rect 34428 11500 34480 11509
rect 35440 11543 35492 11552
rect 35440 11509 35449 11543
rect 35449 11509 35483 11543
rect 35483 11509 35492 11543
rect 35440 11500 35492 11509
rect 38384 11500 38436 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 25596 11339 25648 11348
rect 25596 11305 25605 11339
rect 25605 11305 25639 11339
rect 25639 11305 25648 11339
rect 25596 11296 25648 11305
rect 29184 11339 29236 11348
rect 29184 11305 29193 11339
rect 29193 11305 29227 11339
rect 29227 11305 29236 11339
rect 29184 11296 29236 11305
rect 30656 11296 30708 11348
rect 31024 11296 31076 11348
rect 31944 11296 31996 11348
rect 32220 11339 32272 11348
rect 32220 11305 32229 11339
rect 32229 11305 32263 11339
rect 32263 11305 32272 11339
rect 32220 11296 32272 11305
rect 27528 11228 27580 11280
rect 36912 11228 36964 11280
rect 26424 11160 26476 11212
rect 27160 11160 27212 11212
rect 33600 11203 33652 11212
rect 33600 11169 33609 11203
rect 33609 11169 33643 11203
rect 33643 11169 33652 11203
rect 33600 11160 33652 11169
rect 29828 11092 29880 11144
rect 34152 11135 34204 11144
rect 34152 11101 34161 11135
rect 34161 11101 34195 11135
rect 34195 11101 34204 11135
rect 34152 11092 34204 11101
rect 37648 11160 37700 11212
rect 26148 11024 26200 11076
rect 28356 11024 28408 11076
rect 30564 11024 30616 11076
rect 33140 11024 33192 11076
rect 33692 11024 33744 11076
rect 37280 11092 37332 11144
rect 38384 11160 38436 11212
rect 41052 11296 41104 11348
rect 41144 11296 41196 11348
rect 42340 11339 42392 11348
rect 42340 11305 42349 11339
rect 42349 11305 42383 11339
rect 42383 11305 42392 11339
rect 42340 11296 42392 11305
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 40132 11024 40184 11076
rect 40408 11135 40460 11144
rect 40408 11101 40417 11135
rect 40417 11101 40451 11135
rect 40451 11101 40460 11135
rect 40408 11092 40460 11101
rect 42984 11296 43036 11348
rect 43076 11228 43128 11280
rect 42892 11203 42944 11212
rect 42892 11169 42901 11203
rect 42901 11169 42935 11203
rect 42935 11169 42944 11203
rect 42892 11160 42944 11169
rect 37924 10999 37976 11008
rect 37924 10965 37933 10999
rect 37933 10965 37967 10999
rect 37967 10965 37976 10999
rect 37924 10956 37976 10965
rect 39120 10999 39172 11008
rect 39120 10965 39129 10999
rect 39129 10965 39163 10999
rect 39163 10965 39172 10999
rect 39120 10956 39172 10965
rect 39396 10956 39448 11008
rect 40684 11067 40736 11076
rect 40684 11033 40718 11067
rect 40718 11033 40736 11067
rect 40684 11024 40736 11033
rect 41052 11024 41104 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 28356 10795 28408 10804
rect 28356 10761 28365 10795
rect 28365 10761 28399 10795
rect 28399 10761 28408 10795
rect 28356 10752 28408 10761
rect 30012 10752 30064 10804
rect 31760 10795 31812 10804
rect 31760 10761 31769 10795
rect 31769 10761 31803 10795
rect 31803 10761 31812 10795
rect 31760 10752 31812 10761
rect 33140 10752 33192 10804
rect 34152 10752 34204 10804
rect 35440 10752 35492 10804
rect 29000 10616 29052 10668
rect 29828 10616 29880 10668
rect 30932 10616 30984 10668
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 32588 10616 32640 10625
rect 30380 10480 30432 10532
rect 31852 10480 31904 10532
rect 32864 10591 32916 10600
rect 32864 10557 32873 10591
rect 32873 10557 32907 10591
rect 32907 10557 32916 10591
rect 32864 10548 32916 10557
rect 34428 10480 34480 10532
rect 36912 10752 36964 10804
rect 40132 10795 40184 10804
rect 40132 10761 40141 10795
rect 40141 10761 40175 10795
rect 40175 10761 40184 10795
rect 40132 10752 40184 10761
rect 40868 10752 40920 10804
rect 37280 10684 37332 10736
rect 37924 10684 37976 10736
rect 40408 10684 40460 10736
rect 41144 10795 41196 10804
rect 41144 10761 41153 10795
rect 41153 10761 41187 10795
rect 41187 10761 41196 10795
rect 41144 10752 41196 10761
rect 42248 10752 42300 10804
rect 43536 10752 43588 10804
rect 41420 10684 41472 10736
rect 39028 10659 39080 10668
rect 39028 10625 39062 10659
rect 39062 10625 39080 10659
rect 39028 10616 39080 10625
rect 41052 10548 41104 10600
rect 40868 10412 40920 10464
rect 41696 10412 41748 10464
rect 42064 10412 42116 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 30564 10251 30616 10260
rect 30564 10217 30573 10251
rect 30573 10217 30607 10251
rect 30607 10217 30616 10251
rect 30564 10208 30616 10217
rect 30932 10251 30984 10260
rect 30932 10217 30941 10251
rect 30941 10217 30975 10251
rect 30975 10217 30984 10251
rect 30932 10208 30984 10217
rect 38292 10208 38344 10260
rect 39028 10208 39080 10260
rect 40040 10251 40092 10260
rect 40040 10217 40049 10251
rect 40049 10217 40083 10251
rect 40083 10217 40092 10251
rect 40040 10208 40092 10217
rect 40684 10251 40736 10260
rect 40684 10217 40693 10251
rect 40693 10217 40727 10251
rect 40727 10217 40736 10251
rect 40684 10208 40736 10217
rect 42064 10251 42116 10260
rect 42064 10217 42073 10251
rect 42073 10217 42107 10251
rect 42107 10217 42116 10251
rect 42064 10208 42116 10217
rect 31024 10115 31076 10124
rect 31024 10081 31033 10115
rect 31033 10081 31067 10115
rect 31067 10081 31076 10115
rect 31024 10072 31076 10081
rect 42984 10072 43036 10124
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 39396 10047 39448 10056
rect 39396 10013 39405 10047
rect 39405 10013 39439 10047
rect 39439 10013 39448 10047
rect 39396 10004 39448 10013
rect 40868 10047 40920 10056
rect 40868 10013 40877 10047
rect 40877 10013 40911 10047
rect 40911 10013 40920 10047
rect 40868 10004 40920 10013
rect 43996 10004 44048 10056
rect 43260 9868 43312 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 40040 9664 40092 9716
rect 43260 9707 43312 9716
rect 43260 9673 43269 9707
rect 43269 9673 43303 9707
rect 43303 9673 43312 9707
rect 43260 9664 43312 9673
rect 41328 9596 41380 9648
rect 42800 9639 42852 9648
rect 42800 9605 42809 9639
rect 42809 9605 42843 9639
rect 42843 9605 42852 9639
rect 42800 9596 42852 9605
rect 40040 9324 40092 9376
rect 42984 9324 43036 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 41420 9163 41472 9172
rect 41420 9129 41429 9163
rect 41429 9129 41463 9163
rect 41463 9129 41472 9163
rect 41420 9120 41472 9129
rect 43076 9120 43128 9172
rect 43352 9163 43404 9172
rect 43352 9129 43361 9163
rect 43361 9129 43395 9163
rect 43395 9129 43404 9163
rect 43352 9120 43404 9129
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 42892 8576 42944 8628
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 43996 8032 44048 8084
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 43076 6375 43128 6384
rect 43076 6341 43085 6375
rect 43085 6341 43119 6375
rect 43119 6341 43128 6375
rect 43076 6332 43128 6341
rect 43352 6307 43404 6316
rect 43352 6273 43361 6307
rect 43361 6273 43395 6307
rect 43395 6273 43404 6307
rect 43352 6264 43404 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 43352 5899 43404 5908
rect 43352 5865 43361 5899
rect 43361 5865 43395 5899
rect 43395 5865 43404 5899
rect 43352 5856 43404 5865
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 43352 2839 43404 2848
rect 43352 2805 43361 2839
rect 43361 2805 43395 2839
rect 43395 2805 43404 2839
rect 43352 2796 43404 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 42984 2456 43036 2508
rect 43352 2431 43404 2440
rect 43352 2397 43361 2431
rect 43361 2397 43395 2431
rect 43395 2397 43404 2431
rect 43352 2388 43404 2397
rect 43996 2388 44048 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1278 44200 1390 45000
rect 2842 44200 2954 45000
rect 4406 44200 4518 45000
rect 5970 44200 6082 45000
rect 7534 44200 7646 45000
rect 9098 44200 9210 45000
rect 10662 44200 10774 45000
rect 12226 44200 12338 45000
rect 13790 44200 13902 45000
rect 15354 44200 15466 45000
rect 16918 44200 17030 45000
rect 18482 44200 18594 45000
rect 20046 44200 20158 45000
rect 21610 44200 21722 45000
rect 23174 44200 23286 45000
rect 24738 44200 24850 45000
rect 26302 44200 26414 45000
rect 27866 44200 27978 45000
rect 29430 44200 29542 45000
rect 30994 44200 31106 45000
rect 32558 44200 32670 45000
rect 34122 44200 34234 45000
rect 35686 44200 35798 45000
rect 37250 44200 37362 45000
rect 38814 44200 38926 45000
rect 40378 44200 40490 45000
rect 41942 44200 42054 45000
rect 43506 44200 43618 45000
rect 1320 35834 1348 44200
rect 1308 35828 1360 35834
rect 1308 35770 1360 35776
rect 2884 35154 2912 44200
rect 4448 42106 4476 44200
rect 4448 42078 4660 42106
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35222 4660 42078
rect 6012 35290 6040 44200
rect 6000 35284 6052 35290
rect 6000 35226 6052 35232
rect 4620 35216 4672 35222
rect 4620 35158 4672 35164
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 7576 34513 7604 44200
rect 9140 40118 9168 44200
rect 9128 40112 9180 40118
rect 9128 40054 9180 40060
rect 9680 40112 9732 40118
rect 9680 40054 9732 40060
rect 9692 36378 9720 40054
rect 9680 36372 9732 36378
rect 9680 36314 9732 36320
rect 10416 36032 10468 36038
rect 10416 35974 10468 35980
rect 10428 34649 10456 35974
rect 10414 34640 10470 34649
rect 10414 34575 10470 34584
rect 7562 34504 7618 34513
rect 7562 34439 7618 34448
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 10704 33969 10732 44200
rect 12268 35057 12296 44200
rect 13832 42226 13860 44200
rect 15396 42226 15424 44200
rect 13820 42220 13872 42226
rect 13820 42162 13872 42168
rect 15384 42220 15436 42226
rect 15384 42162 15436 42168
rect 16960 40118 16988 44200
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 18328 40044 18380 40050
rect 18328 39986 18380 39992
rect 18340 39642 18368 39986
rect 16120 39636 16172 39642
rect 16120 39578 16172 39584
rect 18328 39636 18380 39642
rect 18328 39578 18380 39584
rect 14464 38208 14516 38214
rect 14464 38150 14516 38156
rect 14476 37466 14504 38150
rect 15200 37936 15252 37942
rect 15198 37904 15200 37913
rect 15252 37904 15254 37913
rect 15198 37839 15254 37848
rect 15566 37632 15622 37641
rect 15566 37567 15622 37576
rect 15580 37466 15608 37567
rect 16132 37466 16160 39578
rect 16580 38956 16632 38962
rect 16580 38898 16632 38904
rect 16212 37664 16264 37670
rect 16212 37606 16264 37612
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 15568 37460 15620 37466
rect 15568 37402 15620 37408
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 14094 36680 14150 36689
rect 14094 36615 14096 36624
rect 14148 36615 14150 36624
rect 14096 36586 14148 36592
rect 12624 36100 12676 36106
rect 12624 36042 12676 36048
rect 12254 35048 12310 35057
rect 12254 34983 12310 34992
rect 10690 33960 10746 33969
rect 10690 33895 10746 33904
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 12636 33114 12664 36042
rect 15580 35834 15608 37402
rect 16132 36854 16160 37402
rect 16224 37330 16252 37606
rect 16592 37398 16620 38898
rect 18052 38888 18104 38894
rect 16946 38856 17002 38865
rect 18052 38830 18104 38836
rect 16946 38791 16948 38800
rect 17000 38791 17002 38800
rect 16948 38762 17000 38768
rect 16670 37496 16726 37505
rect 16670 37431 16672 37440
rect 16724 37431 16726 37440
rect 16672 37402 16724 37408
rect 16580 37392 16632 37398
rect 16580 37334 16632 37340
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 16224 36922 16252 37266
rect 16212 36916 16264 36922
rect 16212 36858 16264 36864
rect 16120 36848 16172 36854
rect 16120 36790 16172 36796
rect 16212 36712 16264 36718
rect 16212 36654 16264 36660
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 16120 35828 16172 35834
rect 16120 35770 16172 35776
rect 14004 35692 14056 35698
rect 14004 35634 14056 35640
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 13728 34944 13780 34950
rect 13728 34886 13780 34892
rect 13740 34406 13768 34886
rect 14016 34746 14044 35634
rect 15488 35290 15516 35634
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15476 35284 15528 35290
rect 15476 35226 15528 35232
rect 15016 35148 15068 35154
rect 15016 35090 15068 35096
rect 14556 35080 14608 35086
rect 14608 35040 14688 35068
rect 14556 35022 14608 35028
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 14476 34610 14504 34954
rect 14660 34610 14688 35040
rect 15028 34678 15056 35090
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 14464 34604 14516 34610
rect 14464 34546 14516 34552
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 13728 34400 13780 34406
rect 13728 34342 13780 34348
rect 13832 34202 13860 34546
rect 14476 34202 14504 34546
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 13268 34128 13320 34134
rect 13268 34070 13320 34076
rect 13280 33998 13308 34070
rect 14660 33998 14688 34546
rect 15120 34542 15148 35022
rect 15200 35012 15252 35018
rect 15200 34954 15252 34960
rect 15212 34610 15240 34954
rect 15396 34950 15424 35226
rect 16132 35154 16160 35770
rect 16224 35562 16252 36654
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16500 35834 16528 36110
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16684 35630 16712 37402
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 16868 36242 16896 36722
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16212 35556 16264 35562
rect 16212 35498 16264 35504
rect 16224 35290 16252 35498
rect 16960 35494 16988 38762
rect 17222 38448 17278 38457
rect 17222 38383 17278 38392
rect 17236 37738 17264 38383
rect 18064 38350 18092 38830
rect 17500 38344 17552 38350
rect 17500 38286 17552 38292
rect 18052 38344 18104 38350
rect 18052 38286 18104 38292
rect 17224 37732 17276 37738
rect 17224 37674 17276 37680
rect 17132 37664 17184 37670
rect 17132 37606 17184 37612
rect 17144 36038 17172 37606
rect 17236 37466 17264 37674
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17512 36854 17540 38286
rect 18236 38276 18288 38282
rect 18236 38218 18288 38224
rect 18248 38010 18276 38218
rect 18236 38004 18288 38010
rect 18236 37946 18288 37952
rect 18524 37806 18552 44200
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 20088 41698 20116 44200
rect 20720 42220 20772 42226
rect 20720 42162 20772 42168
rect 20444 42016 20496 42022
rect 20444 41958 20496 41964
rect 20088 41670 20208 41698
rect 20076 41608 20128 41614
rect 20076 41550 20128 41556
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 18880 41064 18932 41070
rect 18880 41006 18932 41012
rect 18788 40384 18840 40390
rect 18788 40326 18840 40332
rect 18800 39438 18828 40326
rect 18892 39642 18920 41006
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19156 40112 19208 40118
rect 19156 40054 19208 40060
rect 18880 39636 18932 39642
rect 18880 39578 18932 39584
rect 18788 39432 18840 39438
rect 18788 39374 18840 39380
rect 18892 39386 18920 39578
rect 18800 38554 18828 39374
rect 18892 39358 19012 39386
rect 18880 39296 18932 39302
rect 18880 39238 18932 39244
rect 18892 39030 18920 39238
rect 18880 39024 18932 39030
rect 18880 38966 18932 38972
rect 18788 38548 18840 38554
rect 18788 38490 18840 38496
rect 18984 38418 19012 39358
rect 18972 38412 19024 38418
rect 18972 38354 19024 38360
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 17776 37460 17828 37466
rect 17776 37402 17828 37408
rect 17500 36848 17552 36854
rect 17500 36790 17552 36796
rect 17788 36378 17816 37402
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 19168 36242 19196 40054
rect 19892 40044 19944 40050
rect 19892 39986 19944 39992
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19904 39386 19932 39986
rect 20088 39982 20116 41550
rect 20076 39976 20128 39982
rect 20076 39918 20128 39924
rect 19444 38554 19472 39374
rect 19904 39358 20024 39386
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19996 39098 20024 39358
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 19800 38820 19852 38826
rect 19800 38762 19852 38768
rect 19432 38548 19484 38554
rect 19432 38490 19484 38496
rect 19432 38412 19484 38418
rect 19432 38354 19484 38360
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19260 38010 19288 38150
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 19444 37806 19472 38354
rect 19812 38350 19840 38762
rect 20180 38350 20208 41670
rect 20456 41546 20484 41958
rect 20444 41540 20496 41546
rect 20444 41482 20496 41488
rect 20732 41002 20760 42162
rect 21456 42084 21508 42090
rect 21456 42026 21508 42032
rect 21364 41472 21416 41478
rect 21364 41414 21416 41420
rect 21376 41206 21404 41414
rect 21468 41274 21496 42026
rect 21456 41268 21508 41274
rect 21456 41210 21508 41216
rect 21364 41200 21416 41206
rect 21364 41142 21416 41148
rect 21548 41200 21600 41206
rect 21548 41142 21600 41148
rect 20720 40996 20772 41002
rect 20720 40938 20772 40944
rect 20628 40520 20680 40526
rect 20628 40462 20680 40468
rect 20640 40118 20668 40462
rect 21088 40384 21140 40390
rect 21088 40326 21140 40332
rect 21272 40384 21324 40390
rect 21272 40326 21324 40332
rect 20628 40112 20680 40118
rect 20628 40054 20680 40060
rect 20640 39642 20668 40054
rect 20720 39840 20772 39846
rect 20720 39782 20772 39788
rect 20628 39636 20680 39642
rect 20628 39578 20680 39584
rect 20732 39438 20760 39782
rect 20812 39568 20864 39574
rect 20812 39510 20864 39516
rect 20720 39432 20772 39438
rect 20720 39374 20772 39380
rect 20536 39364 20588 39370
rect 20536 39306 20588 39312
rect 20548 38826 20576 39306
rect 20536 38820 20588 38826
rect 20536 38762 20588 38768
rect 20260 38752 20312 38758
rect 20260 38694 20312 38700
rect 19800 38344 19852 38350
rect 19800 38286 19852 38292
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 20180 37942 20208 38286
rect 20168 37936 20220 37942
rect 20168 37878 20220 37884
rect 19248 37800 19300 37806
rect 19248 37742 19300 37748
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19260 37194 19288 37742
rect 19444 37398 19472 37742
rect 19432 37392 19484 37398
rect 19432 37334 19484 37340
rect 20076 37392 20128 37398
rect 20076 37334 20128 37340
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19248 37188 19300 37194
rect 19248 37130 19300 37136
rect 19352 36378 19380 37198
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19444 36786 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 19156 36236 19208 36242
rect 19156 36178 19208 36184
rect 17132 36032 17184 36038
rect 17132 35974 17184 35980
rect 18788 36032 18840 36038
rect 18788 35974 18840 35980
rect 17960 35760 18012 35766
rect 17960 35702 18012 35708
rect 17132 35692 17184 35698
rect 17132 35634 17184 35640
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16212 35284 16264 35290
rect 16212 35226 16264 35232
rect 16120 35148 16172 35154
rect 16120 35090 16172 35096
rect 17144 35086 17172 35634
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 15384 34944 15436 34950
rect 15384 34886 15436 34892
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13268 33992 13320 33998
rect 13268 33934 13320 33940
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 14648 33992 14700 33998
rect 14648 33934 14700 33940
rect 12624 33108 12676 33114
rect 12624 33050 12676 33056
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 12636 32026 12664 32846
rect 13084 32836 13136 32842
rect 13084 32778 13136 32784
rect 13096 32230 13124 32778
rect 13188 32502 13216 33934
rect 13280 33114 13308 33934
rect 13556 33658 13584 33934
rect 13820 33856 13872 33862
rect 13820 33798 13872 33804
rect 13832 33658 13860 33798
rect 13544 33652 13596 33658
rect 13544 33594 13596 33600
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13268 33108 13320 33114
rect 13268 33050 13320 33056
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13176 32496 13228 32502
rect 13176 32438 13228 32444
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 13280 32026 13308 32710
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 13268 32020 13320 32026
rect 13268 31962 13320 31968
rect 12716 31952 12768 31958
rect 12636 31900 12716 31906
rect 12636 31894 12768 31900
rect 12636 31878 12756 31894
rect 12636 31822 12664 31878
rect 13372 31822 13400 32846
rect 13924 32434 13952 32846
rect 14096 32768 14148 32774
rect 14096 32710 14148 32716
rect 14108 32434 14136 32710
rect 14292 32502 14320 33934
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15120 33658 15148 33866
rect 15580 33658 15608 34546
rect 15948 33998 15976 34546
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 15752 33856 15804 33862
rect 15752 33798 15804 33804
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14384 33114 14412 33254
rect 14372 33108 14424 33114
rect 14372 33050 14424 33056
rect 14556 32836 14608 32842
rect 14556 32778 14608 32784
rect 14280 32496 14332 32502
rect 14280 32438 14332 32444
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 12624 31816 12676 31822
rect 12624 31758 12676 31764
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 12636 30938 12664 31758
rect 13268 31408 13320 31414
rect 13268 31350 13320 31356
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 11888 30864 11940 30870
rect 11888 30806 11940 30812
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 11900 29646 11928 30806
rect 12912 30734 12940 31078
rect 13280 30938 13308 31350
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11992 29850 12020 30534
rect 12912 30326 12940 30670
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 12820 29306 12848 29582
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12912 29170 12940 30262
rect 13004 30258 13032 30670
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 13004 29850 13032 30194
rect 13084 30116 13136 30122
rect 13084 30058 13136 30064
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 13004 29510 13032 29582
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 13004 29034 13032 29446
rect 12992 29028 13044 29034
rect 12992 28970 13044 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 13004 28014 13032 28970
rect 13096 28966 13124 30058
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13188 29034 13216 29582
rect 13176 29028 13228 29034
rect 13176 28970 13228 28976
rect 13084 28960 13136 28966
rect 13084 28902 13136 28908
rect 13188 28082 13216 28970
rect 13372 28694 13400 31758
rect 13464 31754 13492 32166
rect 14108 31958 14136 32370
rect 14292 32026 14320 32438
rect 14464 32292 14516 32298
rect 14464 32234 14516 32240
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14096 31952 14148 31958
rect 14096 31894 14148 31900
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 14200 31754 14228 31826
rect 14476 31822 14504 32234
rect 14568 32026 14596 32778
rect 15016 32428 15068 32434
rect 15120 32416 15148 33594
rect 15764 33522 15792 33798
rect 15948 33658 15976 33934
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15752 33516 15804 33522
rect 15752 33458 15804 33464
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15936 32768 15988 32774
rect 15936 32710 15988 32716
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15068 32388 15148 32416
rect 15016 32370 15068 32376
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 14464 31816 14516 31822
rect 14464 31758 14516 31764
rect 13452 31748 13504 31754
rect 14200 31726 14412 31754
rect 13452 31690 13504 31696
rect 13452 31204 13504 31210
rect 13452 31146 13504 31152
rect 13464 30734 13492 31146
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 13912 30592 13964 30598
rect 13912 30534 13964 30540
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 13556 29646 13584 29990
rect 13636 29776 13688 29782
rect 13636 29718 13688 29724
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13648 29170 13676 29718
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13360 28688 13412 28694
rect 13360 28630 13412 28636
rect 13464 28558 13492 28902
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 13832 27538 13860 30126
rect 13924 29238 13952 30534
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 14108 29850 14136 30126
rect 14096 29844 14148 29850
rect 14096 29786 14148 29792
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14292 29306 14320 29582
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 13912 29232 13964 29238
rect 13912 29174 13964 29180
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13924 27878 13952 28358
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 14292 26382 14320 26862
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14384 26314 14412 31726
rect 15028 31414 15056 32370
rect 15212 32230 15240 32506
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15212 31822 15240 32166
rect 15396 31958 15424 32710
rect 15948 32366 15976 32710
rect 15936 32360 15988 32366
rect 15936 32302 15988 32308
rect 15384 31952 15436 31958
rect 15384 31894 15436 31900
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 15396 31482 15424 31894
rect 15948 31686 15976 32302
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15016 31408 15068 31414
rect 15016 31350 15068 31356
rect 15028 30938 15056 31350
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 15672 30598 15700 31418
rect 15948 31346 15976 31622
rect 15936 31340 15988 31346
rect 15936 31282 15988 31288
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15856 30734 15884 31214
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 15948 30598 15976 31282
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15936 30592 15988 30598
rect 15936 30534 15988 30540
rect 15948 29646 15976 30534
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 14832 29164 14884 29170
rect 14832 29106 14884 29112
rect 14844 28762 14872 29106
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 14752 28218 14780 28426
rect 15212 28422 15240 29174
rect 15856 29170 15884 29446
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15304 28558 15332 29106
rect 15856 28558 15884 29106
rect 16040 28694 16068 34954
rect 16316 34746 16344 35022
rect 16304 34740 16356 34746
rect 16304 34682 16356 34688
rect 16580 34604 16632 34610
rect 16580 34546 16632 34552
rect 16592 33930 16620 34546
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16776 33998 16804 34478
rect 16868 34202 16896 35022
rect 17236 34950 17264 35430
rect 17972 35086 18000 35702
rect 18420 35624 18472 35630
rect 18420 35566 18472 35572
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 18052 35080 18104 35086
rect 18052 35022 18104 35028
rect 18144 35080 18196 35086
rect 18328 35080 18380 35086
rect 18144 35022 18196 35028
rect 18248 35040 18328 35068
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 17408 34944 17460 34950
rect 17408 34886 17460 34892
rect 17144 34610 17172 34886
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 17236 34082 17264 34886
rect 17420 34610 17448 34886
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17592 34604 17644 34610
rect 17592 34546 17644 34552
rect 17328 34202 17356 34546
rect 17316 34196 17368 34202
rect 17316 34138 17368 34144
rect 17040 34060 17092 34066
rect 17236 34054 17356 34082
rect 17040 34002 17092 34008
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16764 33992 16816 33998
rect 16764 33934 16816 33940
rect 16396 33924 16448 33930
rect 16396 33866 16448 33872
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 16224 32366 16252 32914
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16316 31890 16344 32914
rect 16408 32910 16436 33866
rect 16592 33658 16620 33866
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16488 33448 16540 33454
rect 16488 33390 16540 33396
rect 16500 33114 16528 33390
rect 16684 33114 16712 33934
rect 16856 33856 16908 33862
rect 16856 33798 16908 33804
rect 16868 33504 16896 33798
rect 16948 33516 17000 33522
rect 16868 33476 16948 33504
rect 16948 33458 17000 33464
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16408 32570 16436 32846
rect 16396 32564 16448 32570
rect 16396 32506 16448 32512
rect 16500 32298 16528 33050
rect 16488 32292 16540 32298
rect 16488 32234 16540 32240
rect 16960 32230 16988 33458
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16132 29714 16160 30194
rect 16316 30122 16344 31826
rect 16486 31784 16542 31793
rect 16486 31719 16542 31728
rect 16500 30326 16528 31719
rect 16960 31328 16988 32166
rect 17052 32026 17080 34002
rect 17224 33312 17276 33318
rect 17224 33254 17276 33260
rect 17236 32910 17264 33254
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 17236 31958 17264 32846
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 17236 31414 17264 31894
rect 17328 31754 17356 34054
rect 17604 31793 17632 34546
rect 17972 33998 18000 35022
rect 18064 33998 18092 35022
rect 18156 34066 18184 35022
rect 18144 34060 18196 34066
rect 18144 34002 18196 34008
rect 18248 33998 18276 35040
rect 18328 35022 18380 35028
rect 18432 34610 18460 35566
rect 18800 35494 18828 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 36518
rect 20088 36242 20116 37334
rect 20272 37126 20300 38694
rect 20260 37120 20312 37126
rect 20260 37062 20312 37068
rect 20272 36786 20300 37062
rect 20732 36854 20760 39374
rect 20824 39030 20852 39510
rect 21100 39438 21128 40326
rect 21180 39908 21232 39914
rect 21180 39850 21232 39856
rect 21088 39432 21140 39438
rect 21088 39374 21140 39380
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 21192 38962 21220 39850
rect 21180 38956 21232 38962
rect 21180 38898 21232 38904
rect 21284 38842 21312 40326
rect 20996 38820 21048 38826
rect 20996 38762 21048 38768
rect 21100 38814 21312 38842
rect 20812 38344 20864 38350
rect 20812 38286 20864 38292
rect 20824 37942 20852 38286
rect 20812 37936 20864 37942
rect 20812 37878 20864 37884
rect 20904 37868 20956 37874
rect 20904 37810 20956 37816
rect 20720 36848 20772 36854
rect 20720 36790 20772 36796
rect 20260 36780 20312 36786
rect 20260 36722 20312 36728
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 20180 36174 20208 36518
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20076 36100 20128 36106
rect 20076 36042 20128 36048
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 18788 35488 18840 35494
rect 18788 35430 18840 35436
rect 18800 35154 18828 35430
rect 18788 35148 18840 35154
rect 18788 35090 18840 35096
rect 18512 34944 18564 34950
rect 19996 34921 20024 35770
rect 18512 34886 18564 34892
rect 19982 34912 20038 34921
rect 18524 34610 18552 34886
rect 19574 34844 19882 34853
rect 19982 34847 20038 34856
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 20088 34762 20116 36042
rect 19996 34734 20116 34762
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18064 33522 18092 33934
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17696 32842 17724 33390
rect 18064 33114 18092 33458
rect 18340 33114 18368 33934
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 17684 32836 17736 32842
rect 17684 32778 17736 32784
rect 17590 31784 17646 31793
rect 17328 31726 17448 31754
rect 17224 31408 17276 31414
rect 17224 31350 17276 31356
rect 17040 31340 17092 31346
rect 16960 31300 17040 31328
rect 16960 30598 16988 31300
rect 17040 31282 17092 31288
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16304 30116 16356 30122
rect 16304 30058 16356 30064
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 16316 29646 16344 30058
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16132 29170 16160 29514
rect 16396 29504 16448 29510
rect 16396 29446 16448 29452
rect 16408 29306 16436 29446
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16132 28762 16160 29106
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 16028 28688 16080 28694
rect 16028 28630 16080 28636
rect 16224 28626 16252 29106
rect 16776 29102 16804 30194
rect 16856 29776 16908 29782
rect 16856 29718 16908 29724
rect 16868 29170 16896 29718
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16960 29102 16988 30534
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16776 28762 16804 29038
rect 16764 28756 16816 28762
rect 16764 28698 16816 28704
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16960 28558 16988 29038
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14568 27470 14596 27814
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14752 26874 14780 28154
rect 15120 28014 15148 28358
rect 15212 28082 15240 28358
rect 16960 28218 16988 28494
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 17236 27062 17264 31078
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17328 28626 17356 29446
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17328 28082 17356 28562
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17224 27056 17276 27062
rect 17224 26998 17276 27004
rect 14832 26920 14884 26926
rect 14752 26868 14832 26874
rect 14752 26862 14884 26868
rect 14752 26846 14872 26862
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 13280 25838 13308 26182
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 12912 24410 12940 24754
rect 13280 24750 13308 25774
rect 14292 25498 14320 25842
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 13280 22574 13308 24686
rect 14476 23866 14504 25230
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24070 14688 24550
rect 14648 24064 14700 24070
rect 14648 24006 14700 24012
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14660 23798 14688 24006
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22642 13584 22918
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12544 21486 12572 21830
rect 13280 21622 13308 22510
rect 14292 22234 14320 23054
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14384 22166 14412 22442
rect 14476 22438 14504 22986
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 14384 20806 14412 22102
rect 14476 22030 14504 22374
rect 14752 22098 14780 23802
rect 14844 23730 14872 25638
rect 15304 25362 15332 26318
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15580 25294 15608 25638
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15856 24954 15884 25842
rect 16028 25696 16080 25702
rect 16028 25638 16080 25644
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16040 24818 16068 25638
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24886 17080 25094
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14844 22982 14872 23666
rect 15120 23662 15148 24210
rect 16040 24206 16068 24754
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14936 22098 14964 22442
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 21690 14780 21830
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14752 21554 14780 21626
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 15120 20874 15148 23598
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15212 20942 15240 22374
rect 15304 21690 15332 23666
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15396 23118 15424 23598
rect 15488 23254 15516 23666
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15396 22094 15424 23054
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15488 22234 15516 22714
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15396 22066 15516 22094
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15396 21146 15424 21898
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 13820 20800 13872 20806
rect 13648 20748 13820 20754
rect 13648 20742 13872 20748
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 13648 20726 13860 20742
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 13004 20058 13032 20402
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 13188 19446 13216 20198
rect 13464 19922 13492 20334
rect 13648 19922 13676 20726
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13372 19378 13400 19790
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 13648 17746 13676 19858
rect 13832 19786 13860 20198
rect 14660 20058 14688 20402
rect 15120 20398 15148 20810
rect 15488 20482 15516 22066
rect 15580 21554 15608 22986
rect 15764 21706 15792 23122
rect 16040 22778 16068 24142
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16316 23118 16344 23462
rect 17052 23186 17080 24822
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17236 23118 17264 23598
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15672 21678 15792 21706
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15396 20454 15516 20482
rect 15568 20460 15620 20466
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 15120 19394 15148 20334
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15120 19366 15240 19394
rect 15304 19378 15332 20198
rect 15396 19446 15424 20454
rect 15568 20402 15620 20408
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15212 18970 15240 19366
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14292 17270 14320 17478
rect 14660 17270 14688 17478
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 13004 16182 13032 16934
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 13372 16114 13400 17070
rect 13556 16794 13584 17138
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 14660 16250 14688 17206
rect 14752 16726 14780 17478
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 13372 15026 13400 16050
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15026 14320 15302
rect 14844 15162 14872 18226
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 17338 14964 18158
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 14936 16590 14964 17274
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14844 15026 14872 15098
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 15028 14958 15056 17682
rect 15212 16658 15240 18906
rect 15396 18698 15424 19382
rect 15488 19378 15516 20266
rect 15580 19718 15608 20402
rect 15672 20330 15700 21678
rect 15856 21622 15884 22170
rect 17420 22094 17448 31726
rect 17590 31719 17646 31728
rect 17696 31278 17724 32778
rect 18340 32434 18368 33050
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 17788 31414 17816 32370
rect 17880 31754 17908 32370
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17868 31748 17920 31754
rect 17868 31690 17920 31696
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 31482 18000 31622
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17788 30666 17816 31350
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17500 30116 17552 30122
rect 17500 30058 17552 30064
rect 17512 29646 17540 30058
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17788 26314 17816 30602
rect 17972 30394 18000 31418
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 17880 29646 17908 29990
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17972 29594 18000 30330
rect 18064 30326 18092 31758
rect 18524 31754 18552 34546
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 18696 33448 18748 33454
rect 18696 33390 18748 33396
rect 18708 33046 18736 33390
rect 18696 33040 18748 33046
rect 18696 32982 18748 32988
rect 18604 32564 18656 32570
rect 18708 32552 18736 32982
rect 18656 32524 18736 32552
rect 18604 32506 18656 32512
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18340 31726 18552 31754
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18248 31346 18276 31622
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18142 31240 18198 31249
rect 18142 31175 18198 31184
rect 18156 30938 18184 31175
rect 18234 31104 18290 31113
rect 18234 31039 18290 31048
rect 18144 30932 18196 30938
rect 18144 30874 18196 30880
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 18156 29646 18184 29990
rect 18144 29640 18196 29646
rect 17880 29238 17908 29582
rect 17972 29566 18092 29594
rect 18144 29582 18196 29588
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17868 29232 17920 29238
rect 17868 29174 17920 29180
rect 17972 28626 18000 29446
rect 18064 29306 18092 29566
rect 18156 29306 18184 29582
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18144 29096 18196 29102
rect 18142 29064 18144 29073
rect 18196 29064 18198 29073
rect 18142 28999 18198 29008
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 18052 28552 18104 28558
rect 18248 28506 18276 31039
rect 18052 28494 18104 28500
rect 18064 28150 18092 28494
rect 18156 28478 18276 28506
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 18156 27130 18184 28478
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18248 28082 18276 28358
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 18156 25430 18184 27066
rect 18144 25424 18196 25430
rect 18144 25366 18196 25372
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17512 24886 17540 25094
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17696 24410 17724 25230
rect 18340 24970 18368 31726
rect 18512 31476 18564 31482
rect 18512 31418 18564 31424
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18432 30190 18460 30738
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18432 29209 18460 30126
rect 18418 29200 18474 29209
rect 18418 29135 18474 29144
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28694 18460 28902
rect 18420 28688 18472 28694
rect 18420 28630 18472 28636
rect 18524 28558 18552 31418
rect 18616 31346 18644 32370
rect 18708 32230 18736 32524
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18604 31340 18656 31346
rect 18604 31282 18656 31288
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18800 31113 18828 33934
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19248 33448 19300 33454
rect 19248 33390 19300 33396
rect 19156 33312 19208 33318
rect 19156 33254 19208 33260
rect 19168 32434 19196 33254
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18892 31482 18920 31758
rect 18880 31476 18932 31482
rect 18880 31418 18932 31424
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18786 31104 18842 31113
rect 18786 31039 18842 31048
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18800 30326 18828 30874
rect 18892 30734 18920 31214
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 18604 29844 18656 29850
rect 18604 29786 18656 29792
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18616 29238 18644 29786
rect 18708 29646 18736 29786
rect 18984 29646 19012 32370
rect 19076 31958 19104 32370
rect 19260 32298 19288 33390
rect 19352 33318 19380 33866
rect 19996 33862 20024 34734
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33658 20024 33798
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19430 33552 19486 33561
rect 19430 33487 19486 33496
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 19352 32434 19380 33254
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19248 32292 19300 32298
rect 19248 32234 19300 32240
rect 19064 31952 19116 31958
rect 19064 31894 19116 31900
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 19076 31278 19104 31758
rect 19248 31680 19300 31686
rect 19248 31622 19300 31628
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 19168 31124 19196 31418
rect 19076 31096 19196 31124
rect 18696 29640 18748 29646
rect 18880 29640 18932 29646
rect 18696 29582 18748 29588
rect 18878 29608 18880 29617
rect 18972 29640 19024 29646
rect 18932 29608 18934 29617
rect 18972 29582 19024 29588
rect 18878 29543 18934 29552
rect 18984 29306 19012 29582
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 18604 29232 18656 29238
rect 18604 29174 18656 29180
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 18984 29073 19012 29106
rect 18970 29064 19026 29073
rect 18970 28999 19026 29008
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18984 27470 19012 28999
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18524 25906 18552 26726
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18616 25838 18644 26182
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18248 24942 18368 24970
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23866 18184 24006
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17696 23322 17724 23666
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17880 23186 17908 23734
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17604 22710 17632 23054
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17604 22166 17632 22646
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 17236 22066 17448 22094
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15764 20398 15792 21490
rect 15856 20942 15884 21558
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16132 20942 16160 21286
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19514 15608 19654
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15672 19378 15700 19994
rect 15764 19446 15792 20334
rect 15856 19854 15884 20878
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15948 19514 15976 20402
rect 16316 20058 16344 21490
rect 17144 21146 17172 21490
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16592 19718 16620 20742
rect 17236 20602 17264 22066
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15488 19258 15516 19314
rect 15488 19230 15700 19258
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15304 17202 15332 18362
rect 15396 18358 15424 18634
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15672 18290 15700 19230
rect 15764 18426 15792 19382
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17678 15516 18022
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15580 17338 15608 18226
rect 15672 17678 15700 18226
rect 15764 17678 15792 18226
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15502 15148 16050
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15120 15094 15148 15438
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15304 15162 15332 15370
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 14476 13530 14504 13874
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14844 13326 14872 14214
rect 15120 14006 15148 15030
rect 15488 14822 15516 16594
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16250 15608 16526
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15672 15502 15700 16390
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15764 15162 15792 16118
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14482 15516 14758
rect 15764 14482 15792 15098
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15488 13530 15516 14418
rect 15856 14414 15884 17614
rect 16868 17202 16896 19722
rect 16960 19378 16988 19858
rect 17512 19854 17540 21286
rect 17696 20466 17724 22986
rect 17880 21554 17908 23122
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 18064 22098 18092 22578
rect 18156 22098 18184 23802
rect 18248 23254 18276 24942
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 24274 18368 24754
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18236 23248 18288 23254
rect 18236 23190 18288 23196
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17880 20754 17908 21490
rect 18064 21350 18092 22034
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18248 21010 18276 21354
rect 18340 21010 18368 24210
rect 18432 22710 18460 24550
rect 18616 24138 18644 24550
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18616 23662 18644 24074
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18524 22642 18552 22918
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18616 22166 18644 23054
rect 18984 22778 19012 23666
rect 19076 23050 19104 31096
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19168 30002 19196 30534
rect 19260 30122 19288 31622
rect 19444 30802 19472 33487
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19628 32978 19656 33390
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 31890 20024 32710
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 20088 31754 20116 34546
rect 20272 33561 20300 36722
rect 20628 34536 20680 34542
rect 20534 34504 20590 34513
rect 20628 34478 20680 34484
rect 20534 34439 20536 34448
rect 20588 34439 20590 34448
rect 20536 34410 20588 34416
rect 20536 34128 20588 34134
rect 20536 34070 20588 34076
rect 20444 33856 20496 33862
rect 20444 33798 20496 33804
rect 20258 33552 20314 33561
rect 20168 33516 20220 33522
rect 20258 33487 20314 33496
rect 20168 33458 20220 33464
rect 20180 32570 20208 33458
rect 20260 33448 20312 33454
rect 20260 33390 20312 33396
rect 20272 33114 20300 33390
rect 20352 33312 20404 33318
rect 20352 33254 20404 33260
rect 20260 33108 20312 33114
rect 20260 33050 20312 33056
rect 20364 32858 20392 33254
rect 20456 32978 20484 33798
rect 20444 32972 20496 32978
rect 20444 32914 20496 32920
rect 20364 32830 20484 32858
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20168 32564 20220 32570
rect 20168 32506 20220 32512
rect 20260 32292 20312 32298
rect 20260 32234 20312 32240
rect 20088 31726 20208 31754
rect 19800 31680 19852 31686
rect 20076 31680 20128 31686
rect 19852 31640 20024 31668
rect 19800 31622 19852 31628
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31414 20024 31640
rect 20076 31622 20128 31628
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19524 31340 19576 31346
rect 19576 31300 19748 31328
rect 19524 31282 19576 31288
rect 19720 31260 19748 31300
rect 19984 31272 20036 31278
rect 19720 31232 19840 31260
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19708 30728 19760 30734
rect 19812 30716 19840 31232
rect 19984 31214 20036 31220
rect 19996 31113 20024 31214
rect 19982 31104 20038 31113
rect 19982 31039 20038 31048
rect 19892 30728 19944 30734
rect 19812 30688 19892 30716
rect 19708 30670 19760 30676
rect 19944 30688 20024 30716
rect 19892 30670 19944 30676
rect 19352 30326 19380 30670
rect 19720 30598 19748 30670
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19708 30592 19760 30598
rect 19708 30534 19760 30540
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19444 30274 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 30394 20024 30688
rect 20088 30598 20116 31622
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 19984 30388 20036 30394
rect 19984 30330 20036 30336
rect 19444 30258 19564 30274
rect 19996 30258 20024 30330
rect 19444 30252 19576 30258
rect 19444 30246 19524 30252
rect 19524 30194 19576 30200
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19248 30116 19300 30122
rect 19248 30058 19300 30064
rect 20180 30054 20208 31726
rect 20272 31414 20300 32234
rect 20364 31890 20392 32710
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20260 31408 20312 31414
rect 20260 31350 20312 31356
rect 20272 30190 20300 31350
rect 20456 31278 20484 32830
rect 20548 32609 20576 34070
rect 20640 32881 20668 34478
rect 20732 34474 20760 36790
rect 20916 35290 20944 37810
rect 21008 37806 21036 38762
rect 21100 37942 21128 38814
rect 21364 38752 21416 38758
rect 21364 38694 21416 38700
rect 21088 37936 21140 37942
rect 21088 37878 21140 37884
rect 20996 37800 21048 37806
rect 20996 37742 21048 37748
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 20824 34542 20852 35226
rect 20812 34536 20864 34542
rect 20812 34478 20864 34484
rect 20720 34468 20772 34474
rect 20720 34410 20772 34416
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 20824 34105 20852 34342
rect 20810 34096 20866 34105
rect 21100 34066 21128 37878
rect 21272 37868 21324 37874
rect 21272 37810 21324 37816
rect 21284 37398 21312 37810
rect 21376 37738 21404 38694
rect 21456 38548 21508 38554
rect 21456 38490 21508 38496
rect 21468 38282 21496 38490
rect 21560 38418 21588 41142
rect 21652 41138 21680 44200
rect 22744 42220 22796 42226
rect 22744 42162 22796 42168
rect 22100 42016 22152 42022
rect 22100 41958 22152 41964
rect 22560 42016 22612 42022
rect 22560 41958 22612 41964
rect 21640 41132 21692 41138
rect 21640 41074 21692 41080
rect 21824 41132 21876 41138
rect 21824 41074 21876 41080
rect 21640 38548 21692 38554
rect 21640 38490 21692 38496
rect 21548 38412 21600 38418
rect 21548 38354 21600 38360
rect 21560 38321 21588 38354
rect 21652 38350 21680 38490
rect 21836 38350 21864 41074
rect 22112 41002 22140 41958
rect 22572 41614 22600 41958
rect 22560 41608 22612 41614
rect 22560 41550 22612 41556
rect 22756 41274 22784 42162
rect 23216 41414 23244 44200
rect 24780 44146 24808 44200
rect 24780 44118 24900 44146
rect 23388 42016 23440 42022
rect 23388 41958 23440 41964
rect 23216 41386 23336 41414
rect 22744 41268 22796 41274
rect 22744 41210 22796 41216
rect 23308 41070 23336 41386
rect 23400 41070 23428 41958
rect 24124 41472 24176 41478
rect 24124 41414 24176 41420
rect 24136 41138 24164 41414
rect 24124 41132 24176 41138
rect 24124 41074 24176 41080
rect 23296 41064 23348 41070
rect 23296 41006 23348 41012
rect 23388 41064 23440 41070
rect 23388 41006 23440 41012
rect 22100 40996 22152 41002
rect 22100 40938 22152 40944
rect 22652 40928 22704 40934
rect 22652 40870 22704 40876
rect 22560 40384 22612 40390
rect 22560 40326 22612 40332
rect 22376 40180 22428 40186
rect 22376 40122 22428 40128
rect 22192 39568 22244 39574
rect 22192 39510 22244 39516
rect 22204 39370 22232 39510
rect 22192 39364 22244 39370
rect 22192 39306 22244 39312
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22112 38554 22140 38898
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 21640 38344 21692 38350
rect 21546 38312 21602 38321
rect 21456 38276 21508 38282
rect 21640 38286 21692 38292
rect 21824 38344 21876 38350
rect 21824 38286 21876 38292
rect 21546 38247 21602 38256
rect 21456 38218 21508 38224
rect 22008 38208 22060 38214
rect 22008 38150 22060 38156
rect 21454 38040 21510 38049
rect 21454 37975 21510 37984
rect 21468 37874 21496 37975
rect 21456 37868 21508 37874
rect 21456 37810 21508 37816
rect 21364 37732 21416 37738
rect 21364 37674 21416 37680
rect 21916 37664 21968 37670
rect 21916 37606 21968 37612
rect 21272 37392 21324 37398
rect 21272 37334 21324 37340
rect 21928 37330 21956 37606
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 21548 36644 21600 36650
rect 21548 36586 21600 36592
rect 21560 36378 21588 36586
rect 21548 36372 21600 36378
rect 21548 36314 21600 36320
rect 21560 35834 21588 36314
rect 22020 35873 22048 38150
rect 22112 37874 22140 38490
rect 22284 37936 22336 37942
rect 22284 37878 22336 37884
rect 22100 37868 22152 37874
rect 22100 37810 22152 37816
rect 22006 35864 22062 35873
rect 21548 35828 21600 35834
rect 22006 35799 22062 35808
rect 21548 35770 21600 35776
rect 22020 35766 22048 35799
rect 22112 35766 22140 37810
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 22008 35760 22060 35766
rect 22008 35702 22060 35708
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22098 35320 22154 35329
rect 22098 35255 22154 35264
rect 22112 35086 22140 35255
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22020 34134 22048 35022
rect 22112 34950 22140 35022
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22204 34202 22232 37198
rect 22296 36961 22324 37878
rect 22388 37126 22416 40122
rect 22468 39024 22520 39030
rect 22468 38966 22520 38972
rect 22480 38554 22508 38966
rect 22572 38962 22600 40326
rect 22664 40050 22692 40870
rect 22928 40588 22980 40594
rect 22928 40530 22980 40536
rect 22744 40384 22796 40390
rect 22744 40326 22796 40332
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22664 39846 22692 39986
rect 22652 39840 22704 39846
rect 22652 39782 22704 39788
rect 22664 38962 22692 39782
rect 22756 39030 22784 40326
rect 22940 39438 22968 40530
rect 23112 40180 23164 40186
rect 23112 40122 23164 40128
rect 23124 39642 23152 40122
rect 23112 39636 23164 39642
rect 23112 39578 23164 39584
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22928 39296 22980 39302
rect 22928 39238 22980 39244
rect 22744 39024 22796 39030
rect 22744 38966 22796 38972
rect 22560 38956 22612 38962
rect 22560 38898 22612 38904
rect 22652 38956 22704 38962
rect 22652 38898 22704 38904
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 22468 38344 22520 38350
rect 22468 38286 22520 38292
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22282 36952 22338 36961
rect 22480 36922 22508 38286
rect 22572 37913 22600 38898
rect 22664 38486 22692 38898
rect 22652 38480 22704 38486
rect 22652 38422 22704 38428
rect 22558 37904 22614 37913
rect 22664 37874 22692 38422
rect 22756 38418 22784 38966
rect 22744 38412 22796 38418
rect 22744 38354 22796 38360
rect 22744 38276 22796 38282
rect 22744 38218 22796 38224
rect 22558 37839 22614 37848
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 22560 37664 22612 37670
rect 22560 37606 22612 37612
rect 22282 36887 22338 36896
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 22388 36802 22416 36858
rect 22572 36802 22600 37606
rect 22652 37392 22704 37398
rect 22756 37380 22784 38218
rect 22940 38049 22968 39238
rect 23112 38548 23164 38554
rect 23112 38490 23164 38496
rect 22926 38040 22982 38049
rect 22926 37975 22982 37984
rect 22704 37352 22784 37380
rect 22652 37334 22704 37340
rect 22664 37126 22692 37334
rect 22652 37120 22704 37126
rect 22652 37062 22704 37068
rect 22388 36774 22600 36802
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22284 36712 22336 36718
rect 22284 36654 22336 36660
rect 22560 36712 22612 36718
rect 22560 36654 22612 36660
rect 22296 36417 22324 36654
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22282 36408 22338 36417
rect 22282 36343 22338 36352
rect 22388 35714 22416 36518
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 22480 35834 22508 36110
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22388 35686 22508 35714
rect 22480 35018 22508 35686
rect 22572 35154 22600 36654
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22664 35086 22692 36722
rect 22836 36644 22888 36650
rect 22836 36586 22888 36592
rect 22848 36174 22876 36586
rect 22940 36378 22968 37975
rect 23124 37942 23152 38490
rect 23204 38208 23256 38214
rect 23204 38150 23256 38156
rect 23112 37936 23164 37942
rect 23018 37904 23074 37913
rect 23112 37878 23164 37884
rect 23018 37839 23074 37848
rect 22928 36372 22980 36378
rect 22928 36314 22980 36320
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22928 36168 22980 36174
rect 22928 36110 22980 36116
rect 22940 35766 22968 36110
rect 22928 35760 22980 35766
rect 22928 35702 22980 35708
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22848 35018 22876 35634
rect 22468 35012 22520 35018
rect 22468 34954 22520 34960
rect 22836 35012 22888 35018
rect 22836 34954 22888 34960
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22192 34196 22244 34202
rect 22192 34138 22244 34144
rect 22008 34128 22060 34134
rect 21454 34096 21510 34105
rect 20810 34031 20866 34040
rect 21088 34060 21140 34066
rect 22008 34070 22060 34076
rect 21454 34031 21510 34040
rect 21088 34002 21140 34008
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 20720 33380 20772 33386
rect 20720 33322 20772 33328
rect 20732 32910 20760 33322
rect 20720 32904 20772 32910
rect 20626 32872 20682 32881
rect 20772 32864 20852 32892
rect 20720 32846 20772 32852
rect 20626 32807 20682 32816
rect 20534 32600 20590 32609
rect 20534 32535 20590 32544
rect 20548 32366 20576 32535
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20548 31822 20576 32302
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20536 31816 20588 31822
rect 20536 31758 20588 31764
rect 20444 31272 20496 31278
rect 20364 31232 20444 31260
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20168 30048 20220 30054
rect 19168 29974 19472 30002
rect 20168 29990 20220 29996
rect 19154 29608 19210 29617
rect 19154 29543 19210 29552
rect 19340 29572 19392 29578
rect 19168 29510 19196 29543
rect 19340 29514 19392 29520
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19352 29102 19380 29514
rect 19444 29170 19472 29974
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19982 29336 20038 29345
rect 20088 29306 20116 29582
rect 19982 29271 20038 29280
rect 20076 29300 20128 29306
rect 19996 29238 20024 29271
rect 20076 29242 20128 29248
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 20074 29200 20130 29209
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 19352 28762 19380 29038
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19996 28558 20024 29174
rect 20074 29135 20130 29144
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 27946 20024 28494
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25838 19380 26318
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19444 25498 19472 27338
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 19812 26450 19840 26726
rect 19800 26444 19852 26450
rect 19800 26386 19852 26392
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19444 25226 19472 25434
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19444 24954 19472 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 20088 24698 20116 29135
rect 20180 28762 20208 29582
rect 20272 29102 20300 30126
rect 20364 29850 20392 31232
rect 20444 31214 20496 31220
rect 20640 31210 20668 31894
rect 20628 31204 20680 31210
rect 20628 31146 20680 31152
rect 20732 30938 20760 31962
rect 20824 31278 20852 32864
rect 20916 32842 20944 33866
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21284 33318 21312 33458
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21284 32978 21312 33254
rect 21272 32972 21324 32978
rect 21272 32914 21324 32920
rect 20904 32836 20956 32842
rect 20904 32778 20956 32784
rect 20916 32570 20944 32778
rect 20904 32564 20956 32570
rect 20904 32506 20956 32512
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 20916 31754 20944 31826
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 20904 31748 20956 31754
rect 20904 31690 20956 31696
rect 21100 31482 21128 31758
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20456 30258 20484 30738
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20364 29238 20392 29582
rect 20352 29232 20404 29238
rect 20352 29174 20404 29180
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 28756 20220 28762
rect 20168 28698 20220 28704
rect 20364 28490 20392 29174
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20456 27606 20484 29990
rect 20548 29306 20576 30534
rect 20640 30394 20668 30874
rect 20996 30864 21048 30870
rect 20996 30806 21048 30812
rect 20628 30388 20680 30394
rect 20628 30330 20680 30336
rect 21008 29850 21036 30806
rect 21100 30734 21128 31418
rect 21376 31346 21404 31758
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 21272 31272 21324 31278
rect 21272 31214 21324 31220
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21100 30326 21128 30670
rect 21088 30320 21140 30326
rect 21088 30262 21140 30268
rect 21192 30190 21220 30670
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21284 30122 21312 31214
rect 21376 30870 21404 31282
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 21272 30116 21324 30122
rect 21272 30058 21324 30064
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 21008 29578 21036 29786
rect 21192 29646 21220 29990
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20996 29572 21048 29578
rect 20996 29514 21048 29520
rect 21468 29306 21496 34031
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 21916 33040 21968 33046
rect 21836 32988 21916 32994
rect 21836 32982 21968 32988
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 21836 32966 21956 32982
rect 21652 31278 21680 32914
rect 21732 32836 21784 32842
rect 21836 32824 21864 32966
rect 22100 32904 22152 32910
rect 22100 32846 22152 32852
rect 21784 32796 21864 32824
rect 21732 32778 21784 32784
rect 22112 32570 22140 32846
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 21916 31884 21968 31890
rect 21916 31826 21968 31832
rect 21928 31793 21956 31826
rect 21914 31784 21970 31793
rect 21914 31719 21970 31728
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 21640 31272 21692 31278
rect 21640 31214 21692 31220
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21652 30734 21680 31078
rect 21928 30870 21956 31282
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 21916 30864 21968 30870
rect 21916 30806 21968 30812
rect 21640 30728 21692 30734
rect 21640 30670 21692 30676
rect 22112 30433 22140 30874
rect 22098 30424 22154 30433
rect 22098 30359 22154 30368
rect 22008 30252 22060 30258
rect 22008 30194 22060 30200
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 20536 29300 20588 29306
rect 21456 29300 21508 29306
rect 20536 29242 20588 29248
rect 21376 29260 21456 29288
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20548 28558 20576 29106
rect 20628 29096 20680 29102
rect 20628 29038 20680 29044
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20640 28014 20668 29038
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20260 27600 20312 27606
rect 20260 27542 20312 27548
rect 20444 27600 20496 27606
rect 20444 27542 20496 27548
rect 20272 26926 20300 27542
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 19996 24670 20116 24698
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23118 20024 24670
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 24206 20116 24550
rect 20364 24410 20392 26454
rect 20456 25974 20484 26998
rect 20640 26994 20668 27270
rect 20732 27130 20760 28630
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20916 28150 20944 28562
rect 21376 28150 21404 29260
rect 21456 29242 21508 29248
rect 21928 29034 21956 29786
rect 22020 29510 22048 30194
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 22112 28218 22140 30359
rect 22204 29730 22232 33866
rect 22296 32858 22324 34546
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22572 33930 22600 34342
rect 22560 33924 22612 33930
rect 22560 33866 22612 33872
rect 22560 33516 22612 33522
rect 22560 33458 22612 33464
rect 22468 33312 22520 33318
rect 22468 33254 22520 33260
rect 22480 32910 22508 33254
rect 22572 32910 22600 33458
rect 22652 33380 22704 33386
rect 22652 33322 22704 33328
rect 22664 32910 22692 33322
rect 22468 32904 22520 32910
rect 22296 32830 22416 32858
rect 22468 32846 22520 32852
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22388 32774 22416 32830
rect 22376 32768 22428 32774
rect 22376 32710 22428 32716
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22284 31680 22336 31686
rect 22284 31622 22336 31628
rect 22296 31346 22324 31622
rect 22388 31414 22416 31690
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22388 30734 22416 31350
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22388 29850 22416 30670
rect 22480 30326 22508 32302
rect 22572 32230 22600 32846
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 31210 22600 32166
rect 22652 31272 22704 31278
rect 22652 31214 22704 31220
rect 22560 31204 22612 31210
rect 22560 31146 22612 31152
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22664 30138 22692 31214
rect 22572 30110 22692 30138
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 22204 29702 22324 29730
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22204 29306 22232 29582
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22296 29186 22324 29702
rect 22572 29646 22600 30110
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22664 29646 22692 29990
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22204 29158 22324 29186
rect 22204 28558 22232 29158
rect 22572 29034 22600 29582
rect 22756 29238 22784 34886
rect 22928 34672 22980 34678
rect 22928 34614 22980 34620
rect 22940 34066 22968 34614
rect 22928 34060 22980 34066
rect 22928 34002 22980 34008
rect 23032 33844 23060 37839
rect 23216 37262 23244 38150
rect 23308 37942 23336 41006
rect 23572 40452 23624 40458
rect 23572 40394 23624 40400
rect 23584 39982 23612 40394
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 23756 39976 23808 39982
rect 23756 39918 23808 39924
rect 23664 39432 23716 39438
rect 23664 39374 23716 39380
rect 23676 39098 23704 39374
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 23388 38752 23440 38758
rect 23388 38694 23440 38700
rect 23296 37936 23348 37942
rect 23296 37878 23348 37884
rect 23296 37800 23348 37806
rect 23296 37742 23348 37748
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 23124 36854 23152 37198
rect 23112 36848 23164 36854
rect 23112 36790 23164 36796
rect 23204 36576 23256 36582
rect 23202 36544 23204 36553
rect 23256 36544 23258 36553
rect 23202 36479 23258 36488
rect 23308 36281 23336 37742
rect 23400 36718 23428 38694
rect 23570 38312 23626 38321
rect 23570 38247 23626 38256
rect 23584 38214 23612 38247
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23572 37800 23624 37806
rect 23572 37742 23624 37748
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23388 36712 23440 36718
rect 23388 36654 23440 36660
rect 23400 36582 23428 36654
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23294 36272 23350 36281
rect 23294 36207 23350 36216
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23112 35148 23164 35154
rect 23112 35090 23164 35096
rect 22940 33816 23060 33844
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22848 32570 22876 32846
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22940 31686 22968 33816
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 23032 29170 23060 31758
rect 23124 31278 23152 35090
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23216 33930 23244 35022
rect 23308 35018 23336 35566
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23308 34542 23336 34682
rect 23296 34536 23348 34542
rect 23296 34478 23348 34484
rect 23296 34400 23348 34406
rect 23296 34342 23348 34348
rect 23308 33930 23336 34342
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23204 33924 23256 33930
rect 23204 33866 23256 33872
rect 23296 33924 23348 33930
rect 23296 33866 23348 33872
rect 23400 33318 23428 34002
rect 23492 33386 23520 37198
rect 23584 37194 23612 37742
rect 23572 37188 23624 37194
rect 23572 37130 23624 37136
rect 23584 37097 23612 37130
rect 23570 37088 23626 37097
rect 23570 37023 23626 37032
rect 23584 36310 23612 37023
rect 23676 36922 23704 39034
rect 23768 38282 23796 39918
rect 23756 38276 23808 38282
rect 23756 38218 23808 38224
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 36304 23624 36310
rect 23572 36246 23624 36252
rect 23584 35630 23612 36246
rect 23676 36174 23704 36518
rect 23768 36417 23796 38218
rect 23940 38004 23992 38010
rect 23940 37946 23992 37952
rect 23952 37466 23980 37946
rect 24032 37800 24084 37806
rect 24032 37742 24084 37748
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 24044 37330 24072 37742
rect 24136 37466 24164 41074
rect 24872 41070 24900 44118
rect 25412 42220 25464 42226
rect 25412 42162 25464 42168
rect 25044 42016 25096 42022
rect 25044 41958 25096 41964
rect 25228 42016 25280 42022
rect 25228 41958 25280 41964
rect 24952 41608 25004 41614
rect 24952 41550 25004 41556
rect 24860 41064 24912 41070
rect 24860 41006 24912 41012
rect 24308 40724 24360 40730
rect 24308 40666 24360 40672
rect 24216 39908 24268 39914
rect 24216 39850 24268 39856
rect 24228 38826 24256 39850
rect 24216 38820 24268 38826
rect 24216 38762 24268 38768
rect 24320 38185 24348 40666
rect 24964 40594 24992 41550
rect 24952 40588 25004 40594
rect 24952 40530 25004 40536
rect 25056 40526 25084 41958
rect 25240 41546 25268 41958
rect 25228 41540 25280 41546
rect 25228 41482 25280 41488
rect 25424 41274 25452 42162
rect 25412 41268 25464 41274
rect 25412 41210 25464 41216
rect 26344 41070 26372 44200
rect 27068 42356 27120 42362
rect 27068 42298 27120 42304
rect 27080 42022 27108 42298
rect 27528 42288 27580 42294
rect 27528 42230 27580 42236
rect 27344 42220 27396 42226
rect 27344 42162 27396 42168
rect 27436 42220 27488 42226
rect 27436 42162 27488 42168
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 27068 42016 27120 42022
rect 27068 41958 27120 41964
rect 27160 42016 27212 42022
rect 27160 41958 27212 41964
rect 25780 41064 25832 41070
rect 25780 41006 25832 41012
rect 26332 41064 26384 41070
rect 26332 41006 26384 41012
rect 25228 40928 25280 40934
rect 25228 40870 25280 40876
rect 25044 40520 25096 40526
rect 25044 40462 25096 40468
rect 24860 40452 24912 40458
rect 24860 40394 24912 40400
rect 24872 39982 24900 40394
rect 25044 40112 25096 40118
rect 25044 40054 25096 40060
rect 24584 39976 24636 39982
rect 24584 39918 24636 39924
rect 24860 39976 24912 39982
rect 24860 39918 24912 39924
rect 24596 39438 24624 39918
rect 25056 39846 25084 40054
rect 25044 39840 25096 39846
rect 25044 39782 25096 39788
rect 24952 39500 25004 39506
rect 24952 39442 25004 39448
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 24596 39098 24624 39374
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 24412 38554 24440 38898
rect 24400 38548 24452 38554
rect 24400 38490 24452 38496
rect 24306 38176 24362 38185
rect 24306 38111 24362 38120
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24124 37460 24176 37466
rect 24124 37402 24176 37408
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23754 36408 23810 36417
rect 23754 36343 23810 36352
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23676 35766 23704 36110
rect 23664 35760 23716 35766
rect 23664 35702 23716 35708
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23676 35290 23704 35702
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23572 34944 23624 34950
rect 23572 34886 23624 34892
rect 23584 34610 23612 34886
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23676 34542 23704 35226
rect 23768 35034 23796 36343
rect 23860 36242 23888 37198
rect 24136 37194 24164 37402
rect 24124 37188 24176 37194
rect 24124 37130 24176 37136
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24136 36417 24164 36722
rect 24122 36408 24178 36417
rect 24122 36343 24178 36352
rect 24032 36304 24084 36310
rect 24032 36246 24084 36252
rect 23848 36236 23900 36242
rect 23848 36178 23900 36184
rect 23860 35154 23888 36178
rect 23940 36032 23992 36038
rect 23938 36000 23940 36009
rect 23992 36000 23994 36009
rect 23938 35935 23994 35944
rect 24044 35737 24072 36246
rect 24030 35728 24086 35737
rect 23940 35692 23992 35698
rect 24030 35663 24086 35672
rect 23940 35634 23992 35640
rect 23848 35148 23900 35154
rect 23848 35090 23900 35096
rect 23952 35086 23980 35634
rect 23940 35080 23992 35086
rect 23768 35006 23888 35034
rect 23940 35022 23992 35028
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23860 33930 23888 35006
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 23848 33924 23900 33930
rect 23848 33866 23900 33872
rect 23584 33658 23612 33866
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23584 33153 23612 33458
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23570 33144 23626 33153
rect 23570 33079 23626 33088
rect 23768 32978 23796 33390
rect 23846 33008 23902 33017
rect 23756 32972 23808 32978
rect 23676 32932 23756 32960
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23308 31822 23336 32166
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23676 31754 23704 32932
rect 23846 32943 23902 32952
rect 23756 32914 23808 32920
rect 23860 32910 23888 32943
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 24044 32434 24072 35663
rect 24124 34536 24176 34542
rect 24124 34478 24176 34484
rect 24136 33640 24164 34478
rect 24228 34202 24256 37810
rect 24308 37324 24360 37330
rect 24308 37266 24360 37272
rect 24320 36786 24348 37266
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24412 36156 24440 36790
rect 24504 36310 24532 39034
rect 24860 38820 24912 38826
rect 24860 38762 24912 38768
rect 24676 38548 24728 38554
rect 24676 38490 24728 38496
rect 24584 38412 24636 38418
rect 24584 38354 24636 38360
rect 24596 37330 24624 38354
rect 24688 38010 24716 38490
rect 24768 38344 24820 38350
rect 24766 38312 24768 38321
rect 24820 38312 24822 38321
rect 24766 38247 24822 38256
rect 24676 38004 24728 38010
rect 24676 37946 24728 37952
rect 24676 37868 24728 37874
rect 24676 37810 24728 37816
rect 24768 37868 24820 37874
rect 24768 37810 24820 37816
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24688 37126 24716 37810
rect 24780 37369 24808 37810
rect 24766 37360 24822 37369
rect 24766 37295 24822 37304
rect 24872 37262 24900 38762
rect 24860 37256 24912 37262
rect 24860 37198 24912 37204
rect 24964 37194 24992 39442
rect 25056 39438 25084 39782
rect 25044 39432 25096 39438
rect 25044 39374 25096 39380
rect 25044 39296 25096 39302
rect 25044 39238 25096 39244
rect 24952 37188 25004 37194
rect 24952 37130 25004 37136
rect 24676 37120 24728 37126
rect 24676 37062 24728 37068
rect 24766 36952 24822 36961
rect 24766 36887 24822 36896
rect 24780 36854 24808 36887
rect 24768 36848 24820 36854
rect 24768 36790 24820 36796
rect 25056 36786 25084 39238
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25148 38010 25176 38898
rect 25136 38004 25188 38010
rect 25136 37946 25188 37952
rect 25240 37890 25268 40870
rect 25320 38820 25372 38826
rect 25320 38762 25372 38768
rect 25148 37874 25268 37890
rect 25148 37868 25280 37874
rect 25148 37862 25228 37868
rect 25148 37210 25176 37862
rect 25228 37810 25280 37816
rect 25226 37768 25282 37777
rect 25226 37703 25282 37712
rect 25240 37330 25268 37703
rect 25332 37369 25360 38762
rect 25596 38752 25648 38758
rect 25596 38694 25648 38700
rect 25502 38448 25558 38457
rect 25502 38383 25558 38392
rect 25318 37360 25374 37369
rect 25228 37324 25280 37330
rect 25318 37295 25374 37304
rect 25228 37266 25280 37272
rect 25148 37182 25268 37210
rect 24676 36780 24728 36786
rect 24676 36722 24728 36728
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 24492 36304 24544 36310
rect 24492 36246 24544 36252
rect 24584 36168 24636 36174
rect 24412 36128 24532 36156
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24308 35624 24360 35630
rect 24308 35566 24360 35572
rect 24216 34196 24268 34202
rect 24216 34138 24268 34144
rect 24216 33652 24268 33658
rect 24136 33612 24216 33640
rect 24216 33594 24268 33600
rect 24124 33108 24176 33114
rect 24124 33050 24176 33056
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23584 31748 23716 31754
rect 23584 31726 23664 31748
rect 23584 31278 23612 31726
rect 23664 31690 23716 31696
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23572 31272 23624 31278
rect 23572 31214 23624 31220
rect 23400 30938 23428 31214
rect 23388 30932 23440 30938
rect 23388 30874 23440 30880
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23124 30598 23152 30670
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23400 29730 23428 30126
rect 23296 29708 23348 29714
rect 23296 29650 23348 29656
rect 23400 29702 23520 29730
rect 23308 29170 23336 29650
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 21456 28212 21508 28218
rect 21456 28154 21508 28160
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21468 27470 21496 28154
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20640 26518 20668 26930
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20534 26072 20590 26081
rect 20534 26007 20536 26016
rect 20588 26007 20590 26016
rect 20536 25978 20588 25984
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 21284 25906 21312 26250
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20628 24336 20680 24342
rect 20628 24278 20680 24284
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20640 23730 20668 24278
rect 20732 24206 20760 25094
rect 20824 24818 20852 25230
rect 20916 24954 20944 25366
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20916 24818 20944 24890
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 24070 20760 24142
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19352 22778 19380 23054
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18984 22030 19012 22714
rect 19996 22710 20024 23054
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18144 20800 18196 20806
rect 17788 20466 17816 20742
rect 17880 20726 18000 20754
rect 18144 20742 18196 20748
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17696 19530 17724 20402
rect 17972 20398 18000 20726
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 19530 17908 19722
rect 17696 19502 17908 19530
rect 17972 19514 18000 20334
rect 18156 20330 18184 20742
rect 18248 20534 18276 20946
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18248 19718 18276 20470
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17880 19394 17908 19502
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 16948 19372 17000 19378
rect 17880 19366 18000 19394
rect 18340 19378 18368 20198
rect 18800 20058 18828 20266
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 16948 19314 17000 19320
rect 17866 19272 17922 19281
rect 17866 19207 17922 19216
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16960 16182 16988 16458
rect 17052 16454 17080 18702
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 17202 17172 18566
rect 17880 18290 17908 19207
rect 17972 18834 18000 19366
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18290 18000 18770
rect 18236 18760 18288 18766
rect 18340 18748 18368 19314
rect 18288 18720 18368 18748
rect 18236 18702 18288 18708
rect 18616 18290 18644 19450
rect 18984 19310 19012 21286
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 19076 20466 19104 20878
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17224 17672 17276 17678
rect 17222 17640 17224 17649
rect 17276 17640 17278 17649
rect 17222 17575 17278 17584
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17328 16250 17356 17682
rect 17972 17678 18000 18226
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15570 16252 15982
rect 17328 15706 17356 16186
rect 17696 16114 17724 16594
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 14550 15976 14894
rect 16960 14618 16988 15438
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17144 15026 17172 15302
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 17696 14482 17724 16050
rect 17972 15366 18000 16662
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 18064 15162 18092 17614
rect 18156 16250 18184 18158
rect 18616 17678 18644 18226
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18708 17338 18736 18226
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18248 16590 18276 17274
rect 19076 16658 19104 20402
rect 19352 20330 19380 22170
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19444 21622 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19996 21554 20024 21830
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 21490
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19444 20058 19472 20402
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19996 19922 20024 20538
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20088 19666 20116 23462
rect 20824 23322 20852 24550
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20916 23118 20944 24006
rect 21008 23798 21036 25774
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21376 24750 21404 25638
rect 21468 25294 21496 26182
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21468 24614 21496 25230
rect 21916 24948 21968 24954
rect 21916 24890 21968 24896
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21100 24138 21128 24550
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 20996 23792 21048 23798
rect 21048 23752 21128 23780
rect 20996 23734 21048 23740
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 22030 20760 22374
rect 20824 22098 20852 22578
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 19996 19638 20208 19666
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19514 20024 19638
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19168 17202 19196 18702
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19260 18290 19288 18634
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18156 15502 18184 16186
rect 18524 16182 18552 16390
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18616 15706 18644 16526
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 19076 15570 19104 16594
rect 19168 16114 19196 17138
rect 19260 16726 19288 17206
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19352 16114 19380 19110
rect 19996 18630 20024 19314
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19444 16250 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19904 17882 19932 18226
rect 20088 17882 20116 19450
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14074 15884 14350
rect 16224 14074 16252 14418
rect 17512 14074 17540 14418
rect 18064 14414 18092 15098
rect 19168 15026 19196 16050
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 14482 19196 14962
rect 19352 14890 19380 15914
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15162 20024 17546
rect 20180 16726 20208 19638
rect 20272 18358 20300 21898
rect 20916 21622 20944 22442
rect 21008 21690 21036 22918
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 21100 21486 21128 23752
rect 21376 23730 21404 24006
rect 21744 23866 21772 24346
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21836 24206 21864 24278
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21836 23798 21864 24142
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21284 22778 21312 23598
rect 21928 23322 21956 24890
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22020 22114 22048 22170
rect 21928 22098 22048 22114
rect 21916 22092 22048 22098
rect 21968 22086 22048 22092
rect 21916 22034 21968 22040
rect 22020 21486 22048 22086
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 19168 14006 19196 14418
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 19352 13462 19380 14826
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19444 13326 19472 14758
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 15098
rect 20088 15026 20116 15302
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20180 14822 20208 16662
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 15570 20300 15846
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19536 13530 19564 13874
rect 20088 13784 20116 14554
rect 20180 14006 20208 14758
rect 20364 14618 20392 21286
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20456 20602 20484 20810
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20916 20534 20944 20742
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20732 19446 20760 20470
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 19786 20944 20198
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 18766 20760 19246
rect 21100 18970 21128 20402
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21652 20058 21680 20334
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17746 20576 18022
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 17338 20576 17546
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20548 16658 20576 17274
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20732 15094 20760 15506
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20824 14618 20852 18226
rect 20916 17882 20944 18226
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 21008 17762 21036 18090
rect 20916 17734 21036 17762
rect 20916 17542 20944 17734
rect 21100 17542 21128 18226
rect 21192 18086 21220 19382
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21284 18834 21312 19178
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20916 16794 20944 17138
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 21284 16046 21312 18770
rect 21652 18766 21680 19994
rect 22020 19854 22048 21422
rect 22112 21146 22140 21966
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22204 20058 22232 28494
rect 23032 28218 23060 29106
rect 23400 29034 23428 29702
rect 23492 29646 23520 29702
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23480 29504 23532 29510
rect 23480 29446 23532 29452
rect 23492 29306 23520 29446
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23400 28626 23428 28970
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23584 28558 23612 31214
rect 23768 30734 23796 32166
rect 23952 31414 23980 32370
rect 23940 31408 23992 31414
rect 23940 31350 23992 31356
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 24044 29782 24072 31078
rect 24032 29776 24084 29782
rect 24032 29718 24084 29724
rect 23848 29096 23900 29102
rect 23848 29038 23900 29044
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 22928 27872 22980 27878
rect 22928 27814 22980 27820
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22388 26314 22416 26862
rect 22468 26376 22520 26382
rect 22468 26318 22520 26324
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22388 25702 22416 26250
rect 22480 26042 22508 26318
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 23798 22416 24550
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22572 24206 22600 24278
rect 22560 24200 22612 24206
rect 22560 24142 22612 24148
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 22572 23730 22600 24006
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21622 22324 21830
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22296 20942 22324 21082
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 22020 18698 22048 19314
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22296 17882 22324 19314
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 16250 21496 17478
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16794 22232 16934
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21468 15162 21496 16186
rect 21652 15978 21680 16662
rect 22388 16522 22416 22374
rect 22572 20874 22600 23462
rect 22664 22642 22692 27270
rect 22848 27062 22876 27270
rect 22940 27062 22968 27814
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 23676 26994 23704 27542
rect 23768 27470 23796 27950
rect 23860 27606 23888 29038
rect 24032 28416 24084 28422
rect 24032 28358 24084 28364
rect 24044 28150 24072 28358
rect 24032 28144 24084 28150
rect 24032 28086 24084 28092
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 23952 27470 23980 28018
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22756 26382 22784 26726
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22756 25226 22784 26318
rect 22848 25906 22876 26522
rect 23400 26450 23428 26930
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22744 25220 22796 25226
rect 22744 25162 22796 25168
rect 22848 25158 22876 25842
rect 23400 25838 23428 26386
rect 23492 25906 23520 26726
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 23032 25498 23060 25638
rect 23492 25498 23520 25842
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 22836 25152 22888 25158
rect 22836 25094 22888 25100
rect 22848 23322 22876 25094
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22664 22438 22692 22578
rect 22940 22574 22968 24074
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 23032 21894 23060 25434
rect 23492 25294 23520 25434
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 23124 24818 23152 25162
rect 23492 24886 23520 25230
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23124 24342 23152 24754
rect 23584 24750 23612 26522
rect 23676 25906 23704 26930
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23756 25696 23808 25702
rect 23756 25638 23808 25644
rect 23768 25362 23796 25638
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23676 24410 23704 24550
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 23768 24206 23796 25298
rect 23860 25294 23888 25434
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23860 24410 23888 24686
rect 23848 24404 23900 24410
rect 23848 24346 23900 24352
rect 23952 24206 23980 25162
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24044 24682 24072 24890
rect 24032 24676 24084 24682
rect 24032 24618 24084 24624
rect 24044 24206 24072 24618
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23492 23118 23520 23462
rect 23768 23186 23796 23598
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23768 22166 23796 23122
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 23756 22160 23808 22166
rect 23756 22102 23808 22108
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23860 21690 23888 21898
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23400 20942 23428 21286
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19854 22508 20198
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22572 19802 22600 20810
rect 22756 20602 22784 20878
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 23296 19848 23348 19854
rect 22572 19774 22692 19802
rect 23296 19790 23348 19796
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 18426 22600 19654
rect 22664 18766 22692 19774
rect 22742 19544 22798 19553
rect 22742 19479 22744 19488
rect 22796 19479 22798 19488
rect 22744 19450 22796 19456
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22020 15502 22048 15846
rect 22204 15706 22232 16186
rect 22388 16114 22416 16458
rect 22664 16182 22692 18702
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22756 16250 22784 18226
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 22376 16108 22428 16114
rect 22428 16068 22508 16096
rect 22376 16050 22428 16056
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 22388 14618 22416 15506
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20272 14074 20300 14350
rect 20824 14074 20852 14554
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 20168 13796 20220 13802
rect 20088 13756 20168 13784
rect 20168 13738 20220 13744
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20180 12986 20208 13738
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 21284 12850 21312 13126
rect 22020 12850 22048 13262
rect 22204 13258 22232 13942
rect 22388 13802 22416 14554
rect 22480 14006 22508 16068
rect 22664 15434 22692 16118
rect 22848 15502 22876 18158
rect 22940 17678 22968 18158
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22848 15162 22876 15438
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 22480 12238 22508 13670
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22664 12442 22692 13194
rect 23308 13190 23336 19790
rect 23492 18358 23520 20878
rect 23584 20330 23612 20878
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23572 20324 23624 20330
rect 23572 20266 23624 20272
rect 23676 20058 23704 20470
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23584 17882 23612 19858
rect 23768 19854 23796 20402
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19514 23704 19654
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23768 18290 23796 19790
rect 23860 18970 23888 21626
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23952 19310 23980 19994
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 23952 17678 23980 17750
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 23400 16998 23428 17546
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16590 23428 16934
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23400 15706 23428 16050
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23676 15094 23704 15846
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23768 14074 23796 17614
rect 24044 17338 24072 22918
rect 24136 19514 24164 33050
rect 24228 32314 24256 33594
rect 24320 33522 24348 35566
rect 24412 35018 24440 35634
rect 24400 35012 24452 35018
rect 24400 34954 24452 34960
rect 24412 33998 24440 34954
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24308 33516 24360 33522
rect 24308 33458 24360 33464
rect 24320 33114 24348 33458
rect 24308 33108 24360 33114
rect 24308 33050 24360 33056
rect 24306 32464 24362 32473
rect 24412 32450 24440 33798
rect 24504 33386 24532 36128
rect 24582 36136 24584 36145
rect 24636 36136 24638 36145
rect 24582 36071 24638 36080
rect 24582 35864 24638 35873
rect 24582 35799 24638 35808
rect 24596 35766 24624 35799
rect 24584 35760 24636 35766
rect 24584 35702 24636 35708
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24596 35154 24624 35430
rect 24688 35193 24716 36722
rect 24952 36372 25004 36378
rect 24952 36314 25004 36320
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24780 35306 24808 35974
rect 24780 35278 24900 35306
rect 24872 35222 24900 35278
rect 24768 35216 24820 35222
rect 24674 35184 24730 35193
rect 24584 35148 24636 35154
rect 24768 35158 24820 35164
rect 24860 35216 24912 35222
rect 24860 35158 24912 35164
rect 24674 35119 24730 35128
rect 24584 35090 24636 35096
rect 24780 34610 24808 35158
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24872 33658 24900 35022
rect 24860 33652 24912 33658
rect 24860 33594 24912 33600
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24492 33380 24544 33386
rect 24492 33322 24544 33328
rect 24596 32552 24624 33390
rect 24362 32422 24440 32450
rect 24504 32524 24624 32552
rect 24306 32399 24308 32408
rect 24360 32399 24362 32408
rect 24308 32370 24360 32376
rect 24228 32286 24348 32314
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24228 29578 24256 31758
rect 24320 31260 24348 32286
rect 24400 31408 24452 31414
rect 24504 31396 24532 32524
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24596 31754 24624 32370
rect 24688 32337 24716 32438
rect 24674 32328 24730 32337
rect 24674 32263 24730 32272
rect 24780 31958 24808 33526
rect 24964 33454 24992 36314
rect 25056 35329 25084 36722
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 25042 35320 25098 35329
rect 25042 35255 25098 35264
rect 25056 33674 25084 35255
rect 25148 34610 25176 36518
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 25240 34542 25268 37182
rect 25516 36825 25544 38383
rect 25502 36816 25558 36825
rect 25412 36780 25464 36786
rect 25502 36751 25558 36760
rect 25412 36722 25464 36728
rect 25318 36136 25374 36145
rect 25318 36071 25320 36080
rect 25372 36071 25374 36080
rect 25320 36042 25372 36048
rect 25332 35630 25360 36042
rect 25320 35624 25372 35630
rect 25320 35566 25372 35572
rect 25424 35086 25452 36722
rect 25608 36666 25636 38694
rect 25688 38208 25740 38214
rect 25686 38176 25688 38185
rect 25740 38176 25742 38185
rect 25686 38111 25742 38120
rect 25688 37868 25740 37874
rect 25688 37810 25740 37816
rect 25700 37466 25728 37810
rect 25688 37460 25740 37466
rect 25688 37402 25740 37408
rect 25792 37194 25820 41006
rect 26620 40934 26648 41958
rect 27172 41614 27200 41958
rect 26884 41608 26936 41614
rect 26884 41550 26936 41556
rect 27160 41608 27212 41614
rect 27160 41550 27212 41556
rect 26700 41472 26752 41478
rect 26700 41414 26752 41420
rect 26712 41138 26740 41414
rect 26700 41132 26752 41138
rect 26700 41074 26752 41080
rect 26608 40928 26660 40934
rect 26608 40870 26660 40876
rect 25964 40452 26016 40458
rect 25964 40394 26016 40400
rect 26240 40452 26292 40458
rect 26240 40394 26292 40400
rect 25872 38344 25924 38350
rect 25872 38286 25924 38292
rect 25884 38049 25912 38286
rect 25870 38040 25926 38049
rect 25870 37975 25926 37984
rect 25884 37874 25912 37975
rect 25872 37868 25924 37874
rect 25872 37810 25924 37816
rect 25872 37460 25924 37466
rect 25872 37402 25924 37408
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 25884 37097 25912 37402
rect 25870 37088 25926 37097
rect 25870 37023 25926 37032
rect 25884 36922 25912 37023
rect 25872 36916 25924 36922
rect 25872 36858 25924 36864
rect 25870 36816 25926 36825
rect 25780 36780 25832 36786
rect 25870 36751 25872 36760
rect 25780 36722 25832 36728
rect 25924 36751 25926 36760
rect 25872 36722 25924 36728
rect 25516 36638 25636 36666
rect 25516 36174 25544 36638
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25516 36009 25544 36110
rect 25502 36000 25558 36009
rect 25502 35935 25558 35944
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25516 34762 25544 35935
rect 25792 35873 25820 36722
rect 25778 35864 25834 35873
rect 25778 35799 25834 35808
rect 25780 35624 25832 35630
rect 25780 35566 25832 35572
rect 25424 34734 25544 34762
rect 25594 34776 25650 34785
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 25240 34377 25268 34478
rect 25226 34368 25282 34377
rect 25226 34303 25282 34312
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25424 33946 25452 34734
rect 25594 34711 25650 34720
rect 25608 34610 25636 34711
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 25516 34066 25544 34478
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25228 33924 25280 33930
rect 25228 33866 25280 33872
rect 25240 33833 25268 33866
rect 25226 33824 25282 33833
rect 25226 33759 25282 33768
rect 25056 33646 25268 33674
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 25044 33380 25096 33386
rect 25044 33322 25096 33328
rect 25056 32774 25084 33322
rect 25148 32978 25176 33458
rect 25240 33114 25268 33646
rect 25332 33522 25360 33934
rect 25424 33918 25544 33946
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25240 32858 25268 33050
rect 25148 32830 25268 32858
rect 25332 32842 25360 33458
rect 25412 33312 25464 33318
rect 25412 33254 25464 33260
rect 25320 32836 25372 32842
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 24950 32600 25006 32609
rect 24860 32564 24912 32570
rect 24950 32535 24952 32544
rect 24860 32506 24912 32512
rect 25004 32535 25006 32544
rect 24952 32506 25004 32512
rect 24872 32450 24900 32506
rect 24872 32434 24992 32450
rect 24872 32428 25004 32434
rect 24872 32422 24952 32428
rect 24952 32370 25004 32376
rect 24964 32298 24992 32370
rect 24952 32292 25004 32298
rect 24952 32234 25004 32240
rect 25056 32178 25084 32710
rect 24872 32150 25084 32178
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24676 31680 24728 31686
rect 24676 31622 24728 31628
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24452 31368 24532 31396
rect 24400 31350 24452 31356
rect 24688 31346 24716 31622
rect 24780 31414 24808 31622
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 24320 31232 24532 31260
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24216 29572 24268 29578
rect 24216 29514 24268 29520
rect 24320 26353 24348 29990
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24412 29073 24440 29106
rect 24398 29064 24454 29073
rect 24398 28999 24454 29008
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24306 26344 24362 26353
rect 24306 26279 24362 26288
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 24228 24614 24256 24686
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 24228 24138 24256 24550
rect 24216 24132 24268 24138
rect 24216 24074 24268 24080
rect 24320 23798 24348 26279
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24320 19990 24348 20878
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23952 14482 23980 14894
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23768 13530 23796 14010
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23952 13326 23980 14418
rect 24412 14278 24440 27474
rect 24504 27334 24532 31232
rect 24596 29646 24624 31282
rect 24688 30054 24716 31282
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24872 29646 24900 32150
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 24964 31142 24992 31758
rect 25056 31482 25084 31826
rect 25148 31822 25176 32830
rect 25320 32778 25372 32784
rect 25226 32600 25282 32609
rect 25226 32535 25282 32544
rect 25240 32434 25268 32535
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25320 32428 25372 32434
rect 25424 32416 25452 33254
rect 25372 32388 25452 32416
rect 25320 32370 25372 32376
rect 25424 32337 25452 32388
rect 25226 32328 25282 32337
rect 25226 32263 25282 32272
rect 25410 32328 25466 32337
rect 25410 32263 25466 32272
rect 25136 31816 25188 31822
rect 25134 31784 25136 31793
rect 25188 31784 25190 31793
rect 25134 31719 25190 31728
rect 25240 31686 25268 32263
rect 25410 31920 25466 31929
rect 25410 31855 25466 31864
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 24952 31136 25004 31142
rect 25056 31113 25084 31282
rect 24952 31078 25004 31084
rect 25042 31104 25098 31113
rect 25042 31039 25098 31048
rect 24950 30832 25006 30841
rect 24950 30767 25006 30776
rect 24964 30734 24992 30767
rect 25240 30734 25268 31622
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 25044 30116 25096 30122
rect 25044 30058 25096 30064
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 29345 24624 29446
rect 24582 29336 24638 29345
rect 24582 29271 24638 29280
rect 24860 29232 24912 29238
rect 24860 29174 24912 29180
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24780 27470 24808 29038
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 24780 26994 24808 27406
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24504 24206 24532 26726
rect 24872 26450 24900 29174
rect 24964 28994 24992 29650
rect 25056 29170 25084 30058
rect 25148 29306 25176 30534
rect 25240 29578 25268 30670
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 25332 29170 25360 30194
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 24964 28966 25176 28994
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 25056 27538 25084 28358
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24964 27130 24992 27338
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 25056 27010 25084 27474
rect 24964 26982 25084 27010
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24596 25906 24624 26182
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24596 24954 24624 25230
rect 24584 24948 24636 24954
rect 24584 24890 24636 24896
rect 24596 24750 24624 24890
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24780 24410 24808 25298
rect 24872 24614 24900 25842
rect 24964 25498 24992 26982
rect 25044 26920 25096 26926
rect 25044 26862 25096 26868
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24964 24954 24992 25298
rect 24952 24948 25004 24954
rect 24952 24890 25004 24896
rect 24860 24608 24912 24614
rect 24860 24550 24912 24556
rect 24872 24410 24900 24550
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24492 24200 24544 24206
rect 24872 24154 24900 24346
rect 24492 24142 24544 24148
rect 24780 24126 24900 24154
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24504 22778 24532 23666
rect 24780 23186 24808 24126
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24964 23594 24992 23734
rect 24952 23588 25004 23594
rect 24952 23530 25004 23536
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24872 22574 24900 23054
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24596 21010 24624 21966
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24688 20942 24716 21286
rect 24872 21146 24900 22170
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24780 19854 24808 20742
rect 24872 19922 24900 21082
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24504 17814 24532 19790
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 18766 24624 19246
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24492 17808 24544 17814
rect 24492 17750 24544 17756
rect 24596 17678 24624 18702
rect 24780 17882 24808 19790
rect 25056 18426 25084 26862
rect 25148 26042 25176 28966
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25136 26036 25188 26042
rect 25136 25978 25188 25984
rect 25240 25974 25268 26318
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 25240 25498 25268 25910
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25148 24682 25176 25230
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 25240 24206 25268 24686
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 23186 25176 24006
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25332 17882 25360 29106
rect 25424 22642 25452 31855
rect 25516 28234 25544 33918
rect 25700 33658 25728 34546
rect 25688 33652 25740 33658
rect 25688 33594 25740 33600
rect 25688 32904 25740 32910
rect 25688 32846 25740 32852
rect 25596 32224 25648 32230
rect 25596 32166 25648 32172
rect 25608 31686 25636 32166
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25608 30734 25636 31350
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25608 29102 25636 30194
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25700 28422 25728 32846
rect 25792 30734 25820 35566
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25884 34610 25912 35022
rect 25872 34604 25924 34610
rect 25872 34546 25924 34552
rect 25884 33998 25912 34546
rect 25872 33992 25924 33998
rect 25872 33934 25924 33940
rect 25884 33590 25912 33934
rect 25872 33584 25924 33590
rect 25872 33526 25924 33532
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25884 32298 25912 32370
rect 25872 32292 25924 32298
rect 25872 32234 25924 32240
rect 25884 31822 25912 32234
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25884 30734 25912 31758
rect 25976 31260 26004 40394
rect 26252 38570 26280 40394
rect 26332 40384 26384 40390
rect 26332 40326 26384 40332
rect 26344 38826 26372 40326
rect 26516 39500 26568 39506
rect 26516 39442 26568 39448
rect 26528 39370 26556 39442
rect 26516 39364 26568 39370
rect 26516 39306 26568 39312
rect 26332 38820 26384 38826
rect 26332 38762 26384 38768
rect 26424 38752 26476 38758
rect 26424 38694 26476 38700
rect 26160 38542 26280 38570
rect 26160 38457 26188 38542
rect 26146 38448 26202 38457
rect 26146 38383 26202 38392
rect 26240 38344 26292 38350
rect 26238 38312 26240 38321
rect 26292 38312 26294 38321
rect 26238 38247 26294 38256
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26068 36310 26096 37198
rect 26160 36718 26188 37810
rect 26252 37806 26280 38247
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 26344 37942 26372 38150
rect 26332 37936 26384 37942
rect 26332 37878 26384 37884
rect 26240 37800 26292 37806
rect 26436 37788 26464 38694
rect 26528 37856 26556 39306
rect 26712 38350 26740 41074
rect 26896 39982 26924 41550
rect 27356 41274 27384 42162
rect 27344 41268 27396 41274
rect 27344 41210 27396 41216
rect 26976 40928 27028 40934
rect 26976 40870 27028 40876
rect 26884 39976 26936 39982
rect 26884 39918 26936 39924
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 26804 39030 26832 39442
rect 26792 39024 26844 39030
rect 26792 38966 26844 38972
rect 26792 38888 26844 38894
rect 26792 38830 26844 38836
rect 26804 38554 26832 38830
rect 26792 38548 26844 38554
rect 26792 38490 26844 38496
rect 26700 38344 26752 38350
rect 26700 38286 26752 38292
rect 26608 38276 26660 38282
rect 26608 38218 26660 38224
rect 26620 38010 26648 38218
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 26528 37828 26648 37856
rect 26240 37742 26292 37748
rect 26390 37760 26464 37788
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 26056 36304 26108 36310
rect 26056 36246 26108 36252
rect 26252 36174 26280 37742
rect 26390 37652 26418 37760
rect 26516 37732 26568 37738
rect 26620 37720 26648 37828
rect 26568 37692 26648 37720
rect 26516 37674 26568 37680
rect 26390 37624 26464 37652
rect 26332 37392 26384 37398
rect 26332 37334 26384 37340
rect 26436 37346 26464 37624
rect 26344 36786 26372 37334
rect 26436 37318 26648 37346
rect 26424 37256 26476 37262
rect 26424 37198 26476 37204
rect 26436 36922 26464 37198
rect 26424 36916 26476 36922
rect 26424 36858 26476 36864
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 26332 36576 26384 36582
rect 26528 36553 26556 36654
rect 26332 36518 26384 36524
rect 26514 36544 26570 36553
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 26056 36100 26108 36106
rect 26056 36042 26108 36048
rect 26068 35086 26096 36042
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26056 35080 26108 35086
rect 26056 35022 26108 35028
rect 26068 34542 26096 35022
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 26056 33924 26108 33930
rect 26056 33866 26108 33872
rect 26068 33697 26096 33866
rect 26054 33688 26110 33697
rect 26054 33623 26110 33632
rect 26160 32978 26188 35974
rect 26240 35692 26292 35698
rect 26240 35634 26292 35640
rect 26252 34678 26280 35634
rect 26344 35154 26372 36518
rect 26620 36530 26648 37318
rect 26712 36854 26740 38286
rect 26804 37874 26832 38490
rect 26988 38350 27016 40870
rect 27160 39976 27212 39982
rect 27160 39918 27212 39924
rect 27068 39840 27120 39846
rect 27068 39782 27120 39788
rect 26976 38344 27028 38350
rect 26976 38286 27028 38292
rect 26884 38208 26936 38214
rect 26884 38150 26936 38156
rect 26792 37868 26844 37874
rect 26792 37810 26844 37816
rect 26896 37670 26924 38150
rect 26988 38049 27016 38286
rect 26974 38040 27030 38049
rect 26974 37975 27030 37984
rect 26884 37664 26936 37670
rect 26884 37606 26936 37612
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26700 36848 26752 36854
rect 26700 36790 26752 36796
rect 26804 36530 26832 37198
rect 26974 36816 27030 36825
rect 26974 36751 27030 36760
rect 26620 36502 26740 36530
rect 26804 36502 26924 36530
rect 26514 36479 26570 36488
rect 26422 36408 26478 36417
rect 26422 36343 26478 36352
rect 26436 36174 26464 36343
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26528 36106 26556 36479
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26620 36174 26648 36314
rect 26712 36174 26740 36502
rect 26792 36372 26844 36378
rect 26792 36314 26844 36320
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26700 36168 26752 36174
rect 26700 36110 26752 36116
rect 26516 36100 26568 36106
rect 26516 36042 26568 36048
rect 26700 36032 26752 36038
rect 26700 35974 26752 35980
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 26620 35562 26648 35634
rect 26608 35556 26660 35562
rect 26608 35498 26660 35504
rect 26608 35284 26660 35290
rect 26608 35226 26660 35232
rect 26332 35148 26384 35154
rect 26332 35090 26384 35096
rect 26620 35086 26648 35226
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26240 34672 26292 34678
rect 26240 34614 26292 34620
rect 26148 32972 26200 32978
rect 26148 32914 26200 32920
rect 26252 32570 26280 34614
rect 26516 34400 26568 34406
rect 26516 34342 26568 34348
rect 26528 34134 26556 34342
rect 26516 34128 26568 34134
rect 26516 34070 26568 34076
rect 26712 34066 26740 35974
rect 26804 35018 26832 36314
rect 26896 35494 26924 36502
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26792 35012 26844 35018
rect 26792 34954 26844 34960
rect 26792 34196 26844 34202
rect 26792 34138 26844 34144
rect 26700 34060 26752 34066
rect 26700 34002 26752 34008
rect 26422 33960 26478 33969
rect 26422 33895 26478 33904
rect 26436 33862 26464 33895
rect 26424 33856 26476 33862
rect 26330 33824 26386 33833
rect 26424 33798 26476 33804
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 26330 33759 26386 33768
rect 26344 33318 26372 33759
rect 26528 33522 26556 33798
rect 26516 33516 26568 33522
rect 26516 33458 26568 33464
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26240 32564 26292 32570
rect 26160 32524 26240 32552
rect 26056 31748 26108 31754
rect 26056 31690 26108 31696
rect 26068 31414 26096 31690
rect 26160 31482 26188 32524
rect 26240 32506 26292 32512
rect 26240 32292 26292 32298
rect 26240 32234 26292 32240
rect 26252 31686 26280 32234
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26148 31476 26200 31482
rect 26148 31418 26200 31424
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 26148 31272 26200 31278
rect 25976 31232 26148 31260
rect 26148 31214 26200 31220
rect 26056 30864 26108 30870
rect 26056 30806 26108 30812
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 25870 30288 25926 30297
rect 25792 28506 25820 30262
rect 25870 30223 25872 30232
rect 25924 30223 25926 30232
rect 25872 30194 25924 30200
rect 25884 29646 25912 30194
rect 26068 29850 26096 30806
rect 26160 30054 26188 31214
rect 26148 30048 26200 30054
rect 26148 29990 26200 29996
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 25884 28694 25912 28902
rect 25872 28688 25924 28694
rect 25872 28630 25924 28636
rect 25792 28478 25912 28506
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25516 28206 25636 28234
rect 25700 28218 25728 28358
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25516 27606 25544 28018
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25608 26382 25636 28206
rect 25688 28212 25740 28218
rect 25688 28154 25740 28160
rect 25700 27554 25728 28154
rect 25884 27878 25912 28478
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 25700 27526 25820 27554
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25700 27130 25728 27406
rect 25792 27130 25820 27526
rect 25688 27124 25740 27130
rect 25688 27066 25740 27072
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25884 26586 25912 27814
rect 25976 27384 26004 28426
rect 26068 27674 26096 29786
rect 26344 28626 26372 32846
rect 26528 31754 26556 33458
rect 26804 32960 26832 34138
rect 26712 32932 26832 32960
rect 26528 31726 26648 31754
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26332 28620 26384 28626
rect 26332 28562 26384 28568
rect 26056 27668 26108 27674
rect 26056 27610 26108 27616
rect 26056 27396 26108 27402
rect 25976 27356 26056 27384
rect 26056 27338 26108 27344
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25884 26314 25912 26522
rect 26068 26518 26096 27338
rect 26344 27146 26372 28562
rect 26436 28218 26464 29106
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 26344 27118 26464 27146
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26160 26586 26188 26862
rect 26148 26580 26200 26586
rect 26148 26522 26200 26528
rect 26056 26512 26108 26518
rect 26056 26454 26108 26460
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25780 26308 25832 26314
rect 25780 26250 25832 26256
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25700 25906 25728 26182
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25792 25242 25820 26250
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25700 25214 25820 25242
rect 25700 25158 25728 25214
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25424 22094 25452 22578
rect 25700 22506 25728 25094
rect 25884 23866 25912 25978
rect 25976 25362 26004 26386
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 26042 26096 26182
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 26068 25430 26096 25774
rect 26056 25424 26108 25430
rect 26056 25366 26108 25372
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 26160 25158 26188 26318
rect 26252 26042 26280 26862
rect 26344 26518 26372 26930
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 26436 23866 26464 27118
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25976 23322 26004 23666
rect 25964 23316 26016 23322
rect 25964 23258 26016 23264
rect 26436 23118 26464 23802
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 25424 22066 25544 22094
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25424 20602 25452 21898
rect 25516 21690 25544 22066
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25516 21146 25544 21626
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25700 20534 25728 21830
rect 26344 21146 26372 22442
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 25688 20528 25740 20534
rect 25688 20470 25740 20476
rect 25976 20466 26004 21082
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26148 19984 26200 19990
rect 26146 19952 26148 19961
rect 26200 19952 26202 19961
rect 26146 19887 26202 19896
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24596 17270 24624 17614
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 25056 17066 25084 17546
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 25044 17060 25096 17066
rect 25044 17002 25096 17008
rect 24582 16824 24638 16833
rect 24582 16759 24584 16768
rect 24636 16759 24638 16768
rect 24584 16730 24636 16736
rect 25148 16590 25176 17206
rect 25792 17202 25820 17818
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25148 16046 25176 16526
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24964 14618 24992 14962
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 25148 14482 25176 15982
rect 25700 15570 25728 17138
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25228 15360 25280 15366
rect 26056 15360 26108 15366
rect 25228 15302 25280 15308
rect 26054 15328 26056 15337
rect 26108 15328 26110 15337
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25240 14414 25268 15302
rect 26054 15263 26110 15272
rect 26068 15162 26096 15263
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 14074 25268 14214
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24872 13258 24900 13806
rect 25240 13530 25268 14010
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 25148 11762 25176 13262
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25424 11830 25452 12038
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 25608 11354 25636 12174
rect 26160 11898 26188 19887
rect 26528 19514 26556 28630
rect 26620 24290 26648 31726
rect 26712 30326 26740 32932
rect 26792 32836 26844 32842
rect 26792 32778 26844 32784
rect 26804 32298 26832 32778
rect 26882 32464 26938 32473
rect 26988 32434 27016 36751
rect 27080 36718 27108 39782
rect 27172 38894 27200 39918
rect 27160 38888 27212 38894
rect 27160 38830 27212 38836
rect 27068 36712 27120 36718
rect 27068 36654 27120 36660
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 27080 35086 27108 36110
rect 27172 35766 27200 38830
rect 27448 37874 27476 42162
rect 27540 41414 27568 42230
rect 27540 41386 27752 41414
rect 27620 41064 27672 41070
rect 27620 41006 27672 41012
rect 27528 39840 27580 39846
rect 27528 39782 27580 39788
rect 27540 39030 27568 39782
rect 27528 39024 27580 39030
rect 27526 38992 27528 39001
rect 27580 38992 27582 39001
rect 27526 38927 27582 38936
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 27528 37868 27580 37874
rect 27528 37810 27580 37816
rect 27252 37732 27304 37738
rect 27252 37674 27304 37680
rect 27344 37732 27396 37738
rect 27344 37674 27396 37680
rect 27264 37398 27292 37674
rect 27252 37392 27304 37398
rect 27252 37334 27304 37340
rect 27264 37262 27292 37334
rect 27252 37256 27304 37262
rect 27252 37198 27304 37204
rect 27160 35760 27212 35766
rect 27160 35702 27212 35708
rect 27158 35456 27214 35465
rect 27158 35391 27214 35400
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 27080 34202 27108 35022
rect 27068 34196 27120 34202
rect 27068 34138 27120 34144
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 27080 33114 27108 33934
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 27172 32722 27200 35391
rect 27080 32694 27200 32722
rect 26882 32399 26938 32408
rect 26976 32428 27028 32434
rect 26792 32292 26844 32298
rect 26792 32234 26844 32240
rect 26792 31816 26844 31822
rect 26790 31784 26792 31793
rect 26844 31784 26846 31793
rect 26790 31719 26846 31728
rect 26700 30320 26752 30326
rect 26700 30262 26752 30268
rect 26792 30048 26844 30054
rect 26792 29990 26844 29996
rect 26804 29646 26832 29990
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26804 29102 26832 29582
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26712 27713 26740 28562
rect 26804 28150 26832 29038
rect 26792 28144 26844 28150
rect 26792 28086 26844 28092
rect 26698 27704 26754 27713
rect 26698 27639 26754 27648
rect 26700 27600 26752 27606
rect 26700 27542 26752 27548
rect 26712 24818 26740 27542
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 26620 24262 26740 24290
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26620 23594 26648 24142
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26712 23526 26740 24262
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26804 22030 26832 28086
rect 26896 26194 26924 32399
rect 26976 32370 27028 32376
rect 27080 32298 27108 32694
rect 27160 32564 27212 32570
rect 27160 32506 27212 32512
rect 27068 32292 27120 32298
rect 27068 32234 27120 32240
rect 26976 32020 27028 32026
rect 26976 31962 27028 31968
rect 26988 31822 27016 31962
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 26988 28422 27016 28494
rect 27080 28422 27108 28494
rect 26976 28416 27028 28422
rect 26976 28358 27028 28364
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 27080 26382 27108 26726
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26896 26166 27108 26194
rect 26976 25696 27028 25702
rect 26976 25638 27028 25644
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 26896 22438 26924 25094
rect 26884 22432 26936 22438
rect 26884 22374 26936 22380
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26712 18222 26740 18702
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26528 16590 26556 16934
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26240 15632 26292 15638
rect 26240 15574 26292 15580
rect 26252 13802 26280 15574
rect 26424 13932 26476 13938
rect 26528 13920 26556 16526
rect 26606 16280 26662 16289
rect 26896 16266 26924 21490
rect 26988 16454 27016 25638
rect 27080 21554 27108 26166
rect 27172 25974 27200 32506
rect 27264 32502 27292 37198
rect 27356 36922 27384 37674
rect 27448 37641 27476 37810
rect 27434 37632 27490 37641
rect 27434 37567 27490 37576
rect 27540 37466 27568 37810
rect 27528 37460 27580 37466
rect 27528 37402 27580 37408
rect 27632 37262 27660 41006
rect 27724 40526 27752 41386
rect 27908 41138 27936 44200
rect 29472 44130 29500 44200
rect 29460 44124 29512 44130
rect 29460 44066 29512 44072
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 29644 42084 29696 42090
rect 29644 42026 29696 42032
rect 29000 42016 29052 42022
rect 29000 41958 29052 41964
rect 28264 41472 28316 41478
rect 28264 41414 28316 41420
rect 28276 41274 28304 41414
rect 28264 41268 28316 41274
rect 28264 41210 28316 41216
rect 27896 41132 27948 41138
rect 27896 41074 27948 41080
rect 27712 40520 27764 40526
rect 27712 40462 27764 40468
rect 27724 39846 27752 40462
rect 27896 40384 27948 40390
rect 27896 40326 27948 40332
rect 27804 40044 27856 40050
rect 27804 39986 27856 39992
rect 27712 39840 27764 39846
rect 27712 39782 27764 39788
rect 27724 37670 27752 39782
rect 27712 37664 27764 37670
rect 27712 37606 27764 37612
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27356 36786 27568 36802
rect 27356 36780 27580 36786
rect 27356 36774 27528 36780
rect 27356 36224 27384 36774
rect 27528 36722 27580 36728
rect 27436 36712 27488 36718
rect 27488 36660 27568 36666
rect 27436 36654 27568 36660
rect 27448 36638 27568 36654
rect 27356 36196 27476 36224
rect 27344 36100 27396 36106
rect 27344 36042 27396 36048
rect 27356 35737 27384 36042
rect 27342 35728 27398 35737
rect 27342 35663 27398 35672
rect 27342 35048 27398 35057
rect 27342 34983 27398 34992
rect 27356 34678 27384 34983
rect 27344 34672 27396 34678
rect 27344 34614 27396 34620
rect 27448 34542 27476 36196
rect 27540 36106 27568 36638
rect 27620 36576 27672 36582
rect 27620 36518 27672 36524
rect 27528 36100 27580 36106
rect 27528 36042 27580 36048
rect 27540 35766 27568 36042
rect 27632 36009 27660 36518
rect 27724 36145 27752 37062
rect 27816 36174 27844 39986
rect 27908 39953 27936 40326
rect 27894 39944 27950 39953
rect 27894 39879 27950 39888
rect 27988 38344 28040 38350
rect 27988 38286 28040 38292
rect 28172 38344 28224 38350
rect 28276 38332 28304 41210
rect 28540 41064 28592 41070
rect 28540 41006 28592 41012
rect 28356 40452 28408 40458
rect 28356 40394 28408 40400
rect 28368 39506 28396 40394
rect 28356 39500 28408 39506
rect 28356 39442 28408 39448
rect 28368 38826 28396 39442
rect 28356 38820 28408 38826
rect 28356 38762 28408 38768
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 28356 38480 28408 38486
rect 28354 38448 28356 38457
rect 28408 38448 28410 38457
rect 28354 38383 28410 38392
rect 28368 38350 28396 38383
rect 28224 38304 28304 38332
rect 28356 38344 28408 38350
rect 28172 38286 28224 38292
rect 28356 38286 28408 38292
rect 27896 38208 27948 38214
rect 27896 38150 27948 38156
rect 27908 37942 27936 38150
rect 27896 37936 27948 37942
rect 27896 37878 27948 37884
rect 28000 37806 28028 38286
rect 28184 38214 28212 38286
rect 28172 38208 28224 38214
rect 28172 38150 28224 38156
rect 28460 37992 28488 38694
rect 28184 37964 28488 37992
rect 27988 37800 28040 37806
rect 27988 37742 28040 37748
rect 28184 37738 28212 37964
rect 28262 37904 28318 37913
rect 28448 37868 28500 37874
rect 28318 37848 28448 37856
rect 28262 37839 28448 37848
rect 28276 37828 28448 37839
rect 28448 37810 28500 37816
rect 28172 37732 28224 37738
rect 28172 37674 28224 37680
rect 27896 37664 27948 37670
rect 27896 37606 27948 37612
rect 27908 37330 27936 37606
rect 28184 37398 28212 37674
rect 28172 37392 28224 37398
rect 28172 37334 28224 37340
rect 27896 37324 27948 37330
rect 27896 37266 27948 37272
rect 28448 37324 28500 37330
rect 28448 37266 28500 37272
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28080 36780 28132 36786
rect 28080 36722 28132 36728
rect 27804 36168 27856 36174
rect 27710 36136 27766 36145
rect 27804 36110 27856 36116
rect 27710 36071 27766 36080
rect 27618 36000 27674 36009
rect 27618 35935 27674 35944
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27712 35760 27764 35766
rect 27712 35702 27764 35708
rect 27528 35624 27580 35630
rect 27526 35592 27528 35601
rect 27620 35624 27672 35630
rect 27580 35592 27582 35601
rect 27620 35566 27672 35572
rect 27526 35527 27582 35536
rect 27436 34536 27488 34542
rect 27342 34504 27398 34513
rect 27436 34478 27488 34484
rect 27342 34439 27398 34448
rect 27356 33318 27384 34439
rect 27344 33312 27396 33318
rect 27344 33254 27396 33260
rect 27252 32496 27304 32502
rect 27252 32438 27304 32444
rect 27252 32292 27304 32298
rect 27252 32234 27304 32240
rect 27264 31822 27292 32234
rect 27252 31816 27304 31822
rect 27356 31793 27384 33254
rect 27448 32774 27476 34478
rect 27540 33590 27568 35527
rect 27632 33862 27660 35566
rect 27724 35290 27752 35702
rect 27712 35284 27764 35290
rect 27712 35226 27764 35232
rect 27724 33998 27752 35226
rect 27896 35148 27948 35154
rect 27896 35090 27948 35096
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27816 34746 27844 35022
rect 27804 34740 27856 34746
rect 27804 34682 27856 34688
rect 27804 34060 27856 34066
rect 27804 34002 27856 34008
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27620 33856 27672 33862
rect 27620 33798 27672 33804
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 27540 33425 27568 33526
rect 27526 33416 27582 33425
rect 27526 33351 27582 33360
rect 27436 32768 27488 32774
rect 27436 32710 27488 32716
rect 27252 31758 27304 31764
rect 27342 31784 27398 31793
rect 27342 31719 27398 31728
rect 27632 30870 27660 33798
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27724 33318 27752 33390
rect 27712 33312 27764 33318
rect 27712 33254 27764 33260
rect 27816 32978 27844 34002
rect 27908 33998 27936 35090
rect 27988 34944 28040 34950
rect 27988 34886 28040 34892
rect 28000 34610 28028 34886
rect 27988 34604 28040 34610
rect 27988 34546 28040 34552
rect 27986 34232 28042 34241
rect 27986 34167 28042 34176
rect 28000 33998 28028 34167
rect 27896 33992 27948 33998
rect 27896 33934 27948 33940
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 28000 33454 28028 33934
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 28000 32978 28028 33390
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 27988 32972 28040 32978
rect 27988 32914 28040 32920
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27620 30864 27672 30870
rect 27620 30806 27672 30812
rect 27344 30660 27396 30666
rect 27344 30602 27396 30608
rect 27252 30592 27304 30598
rect 27252 30534 27304 30540
rect 27264 30394 27292 30534
rect 27356 30394 27384 30602
rect 27252 30388 27304 30394
rect 27252 30330 27304 30336
rect 27344 30388 27396 30394
rect 27344 30330 27396 30336
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27356 28098 27384 30126
rect 27632 29850 27660 30194
rect 27724 30138 27752 32846
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27816 30326 27844 31758
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27908 30569 27936 30670
rect 27894 30560 27950 30569
rect 27894 30495 27950 30504
rect 27804 30320 27856 30326
rect 27804 30262 27856 30268
rect 27724 30110 27844 30138
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27724 29850 27752 29990
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27816 29782 27844 30110
rect 27804 29776 27856 29782
rect 27804 29718 27856 29724
rect 27712 28688 27764 28694
rect 27712 28630 27764 28636
rect 27356 28070 27476 28098
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27356 27674 27384 27950
rect 27344 27668 27396 27674
rect 27344 27610 27396 27616
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27264 26994 27292 27270
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27356 26874 27384 27270
rect 27264 26846 27384 26874
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27264 25906 27292 26846
rect 27344 26444 27396 26450
rect 27344 26386 27396 26392
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27252 25764 27304 25770
rect 27252 25706 27304 25712
rect 27264 24818 27292 25706
rect 27356 25498 27384 26386
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27448 25226 27476 28070
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27540 25906 27568 27406
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27172 24206 27200 24754
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27172 23186 27200 23462
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27264 22642 27292 23462
rect 27356 23118 27384 24006
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27160 20868 27212 20874
rect 27160 20810 27212 20816
rect 27172 20534 27200 20810
rect 27160 20528 27212 20534
rect 27160 20470 27212 20476
rect 27264 19718 27292 22578
rect 27448 22094 27476 23530
rect 27356 22066 27476 22094
rect 27356 20262 27384 22066
rect 27434 20632 27490 20641
rect 27540 20602 27568 25842
rect 27632 25294 27660 27406
rect 27724 25702 27752 28630
rect 27816 27690 27844 29718
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27908 28014 27936 28358
rect 27896 28008 27948 28014
rect 27896 27950 27948 27956
rect 27816 27662 27936 27690
rect 28000 27674 28028 32914
rect 28092 28490 28120 36722
rect 28172 36100 28224 36106
rect 28172 36042 28224 36048
rect 28184 35222 28212 36042
rect 28172 35216 28224 35222
rect 28172 35158 28224 35164
rect 28172 34944 28224 34950
rect 28172 34886 28224 34892
rect 28184 34610 28212 34886
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28172 34128 28224 34134
rect 28172 34070 28224 34076
rect 28184 32609 28212 34070
rect 28276 33658 28304 37198
rect 28356 35080 28408 35086
rect 28354 35048 28356 35057
rect 28408 35048 28410 35057
rect 28354 34983 28410 34992
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28264 33652 28316 33658
rect 28264 33594 28316 33600
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 28170 32600 28226 32609
rect 28170 32535 28226 32544
rect 28276 32502 28304 33390
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 28368 29306 28396 34546
rect 28460 32230 28488 37266
rect 28552 36922 28580 41006
rect 28908 40452 28960 40458
rect 28908 40394 28960 40400
rect 28724 40044 28776 40050
rect 28724 39986 28776 39992
rect 28736 39642 28764 39986
rect 28724 39636 28776 39642
rect 28724 39578 28776 39584
rect 28920 39438 28948 40394
rect 29012 40338 29040 41958
rect 29656 41682 29684 42026
rect 29644 41676 29696 41682
rect 29644 41618 29696 41624
rect 29092 41608 29144 41614
rect 29092 41550 29144 41556
rect 29104 41274 29132 41550
rect 30668 41274 30696 42162
rect 30840 42016 30892 42022
rect 30840 41958 30892 41964
rect 30852 41614 30880 41958
rect 30840 41608 30892 41614
rect 30840 41550 30892 41556
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 31036 41414 31064 44200
rect 31760 44124 31812 44130
rect 31760 44066 31812 44072
rect 31576 42084 31628 42090
rect 31576 42026 31628 42032
rect 31484 41812 31536 41818
rect 31484 41754 31536 41760
rect 29092 41268 29144 41274
rect 29092 41210 29144 41216
rect 30656 41268 30708 41274
rect 30656 41210 30708 41216
rect 30944 41138 30972 41414
rect 31036 41386 31156 41414
rect 30472 41132 30524 41138
rect 30472 41074 30524 41080
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30288 41064 30340 41070
rect 30288 41006 30340 41012
rect 30104 40928 30156 40934
rect 30104 40870 30156 40876
rect 29828 40384 29880 40390
rect 29012 40310 29408 40338
rect 29828 40326 29880 40332
rect 29184 40180 29236 40186
rect 29184 40122 29236 40128
rect 29092 39840 29144 39846
rect 29092 39782 29144 39788
rect 28908 39432 28960 39438
rect 28908 39374 28960 39380
rect 29000 39296 29052 39302
rect 29000 39238 29052 39244
rect 28632 38956 28684 38962
rect 28632 38898 28684 38904
rect 28644 38554 28672 38898
rect 29012 38865 29040 39238
rect 29104 38962 29132 39782
rect 29092 38956 29144 38962
rect 29092 38898 29144 38904
rect 28998 38856 29054 38865
rect 28998 38791 29054 38800
rect 28908 38752 28960 38758
rect 28906 38720 28908 38729
rect 28960 38720 28962 38729
rect 28906 38655 28962 38664
rect 28632 38548 28684 38554
rect 28632 38490 28684 38496
rect 28632 38344 28684 38350
rect 28630 38312 28632 38321
rect 28684 38312 28686 38321
rect 28630 38247 28686 38256
rect 28906 38312 28962 38321
rect 28906 38247 28962 38256
rect 28722 38040 28778 38049
rect 28722 37975 28778 37984
rect 28632 37936 28684 37942
rect 28632 37878 28684 37884
rect 28644 37466 28672 37878
rect 28632 37460 28684 37466
rect 28632 37402 28684 37408
rect 28540 36916 28592 36922
rect 28540 36858 28592 36864
rect 28630 35864 28686 35873
rect 28630 35799 28686 35808
rect 28644 35630 28672 35799
rect 28540 35624 28592 35630
rect 28540 35566 28592 35572
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 28552 35290 28580 35566
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28552 34474 28580 35226
rect 28644 35018 28672 35566
rect 28632 35012 28684 35018
rect 28632 34954 28684 34960
rect 28644 34921 28672 34954
rect 28630 34912 28686 34921
rect 28630 34847 28686 34856
rect 28540 34468 28592 34474
rect 28540 34410 28592 34416
rect 28552 33658 28580 34410
rect 28540 33652 28592 33658
rect 28540 33594 28592 33600
rect 28552 33318 28580 33594
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28540 32972 28592 32978
rect 28540 32914 28592 32920
rect 28552 32502 28580 32914
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28448 32224 28500 32230
rect 28448 32166 28500 32172
rect 28540 31748 28592 31754
rect 28540 31690 28592 31696
rect 28552 31260 28580 31690
rect 28644 31414 28672 34847
rect 28736 33930 28764 37975
rect 28816 37868 28868 37874
rect 28816 37810 28868 37816
rect 28828 37670 28856 37810
rect 28816 37664 28868 37670
rect 28816 37606 28868 37612
rect 28828 36106 28856 37606
rect 28920 36378 28948 38247
rect 29012 38049 29040 38791
rect 28998 38040 29054 38049
rect 28998 37975 29054 37984
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 29012 36718 29040 37606
rect 29104 37330 29132 38898
rect 29196 38554 29224 40122
rect 29276 38820 29328 38826
rect 29276 38762 29328 38768
rect 29184 38548 29236 38554
rect 29184 38490 29236 38496
rect 29288 38486 29316 38762
rect 29276 38480 29328 38486
rect 29276 38422 29328 38428
rect 29380 37913 29408 40310
rect 29736 39568 29788 39574
rect 29736 39510 29788 39516
rect 29644 39364 29696 39370
rect 29644 39306 29696 39312
rect 29460 39296 29512 39302
rect 29460 39238 29512 39244
rect 29366 37904 29422 37913
rect 29288 37862 29366 37890
rect 29184 37800 29236 37806
rect 29184 37742 29236 37748
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 28908 36372 28960 36378
rect 28908 36314 28960 36320
rect 28816 36100 28868 36106
rect 28816 36042 28868 36048
rect 29104 35834 29132 36722
rect 29196 36174 29224 37742
rect 29288 37369 29316 37862
rect 29366 37839 29422 37848
rect 29274 37360 29330 37369
rect 29274 37295 29330 37304
rect 29276 37256 29328 37262
rect 29276 37198 29328 37204
rect 29288 36786 29316 37198
rect 29368 37188 29420 37194
rect 29368 37130 29420 37136
rect 29276 36780 29328 36786
rect 29276 36722 29328 36728
rect 29288 36310 29316 36722
rect 29276 36304 29328 36310
rect 29276 36246 29328 36252
rect 29184 36168 29236 36174
rect 29184 36110 29236 36116
rect 29380 35873 29408 37130
rect 29472 36786 29500 39238
rect 29656 39098 29684 39306
rect 29644 39092 29696 39098
rect 29644 39034 29696 39040
rect 29552 38548 29604 38554
rect 29552 38490 29604 38496
rect 29460 36780 29512 36786
rect 29460 36722 29512 36728
rect 29366 35864 29422 35873
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 29092 35828 29144 35834
rect 29276 35828 29328 35834
rect 29092 35770 29144 35776
rect 29196 35788 29276 35816
rect 29012 35714 29040 35770
rect 28908 35692 28960 35698
rect 29012 35686 29132 35714
rect 28908 35634 28960 35640
rect 28814 34232 28870 34241
rect 28814 34167 28870 34176
rect 28828 34066 28856 34167
rect 28816 34060 28868 34066
rect 28816 34002 28868 34008
rect 28920 33930 28948 35634
rect 29104 35630 29132 35686
rect 29000 35624 29052 35630
rect 29000 35566 29052 35572
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29012 35057 29040 35566
rect 28998 35048 29054 35057
rect 28998 34983 29054 34992
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29012 34649 29040 34682
rect 29092 34672 29144 34678
rect 28998 34640 29054 34649
rect 29092 34614 29144 34620
rect 28998 34575 29054 34584
rect 29104 34202 29132 34614
rect 29092 34196 29144 34202
rect 29092 34138 29144 34144
rect 29104 34066 29132 34138
rect 29092 34060 29144 34066
rect 29092 34002 29144 34008
rect 28724 33924 28776 33930
rect 28724 33866 28776 33872
rect 28816 33924 28868 33930
rect 28816 33866 28868 33872
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28828 33114 28856 33866
rect 28920 33522 28948 33866
rect 28998 33552 29054 33561
rect 28908 33516 28960 33522
rect 28998 33487 29054 33496
rect 28908 33458 28960 33464
rect 29012 33318 29040 33487
rect 29000 33312 29052 33318
rect 29000 33254 29052 33260
rect 28816 33108 28868 33114
rect 28816 33050 28868 33056
rect 28816 32836 28868 32842
rect 28816 32778 28868 32784
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28736 31822 28764 32166
rect 28828 31958 28856 32778
rect 29012 32774 29040 33254
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 29012 32570 29040 32710
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 29196 32450 29224 35788
rect 29366 35799 29422 35808
rect 29276 35770 29328 35776
rect 29276 35692 29328 35698
rect 29276 35634 29328 35640
rect 29288 35086 29316 35634
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29380 34610 29408 35430
rect 29472 35018 29500 36722
rect 29564 35290 29592 38490
rect 29656 38418 29684 39034
rect 29748 38554 29776 39510
rect 29840 39030 29868 40326
rect 30116 40186 30144 40870
rect 30300 40662 30328 41006
rect 30288 40656 30340 40662
rect 30288 40598 30340 40604
rect 30104 40180 30156 40186
rect 30104 40122 30156 40128
rect 30196 40112 30248 40118
rect 30196 40054 30248 40060
rect 30208 39302 30236 40054
rect 30300 39506 30328 40598
rect 30380 40384 30432 40390
rect 30380 40326 30432 40332
rect 30392 40050 30420 40326
rect 30380 40044 30432 40050
rect 30380 39986 30432 39992
rect 30288 39500 30340 39506
rect 30288 39442 30340 39448
rect 30196 39296 30248 39302
rect 30196 39238 30248 39244
rect 29828 39024 29880 39030
rect 29828 38966 29880 38972
rect 29736 38548 29788 38554
rect 29736 38490 29788 38496
rect 29644 38412 29696 38418
rect 29644 38354 29696 38360
rect 29656 36122 29684 38354
rect 29920 38276 29972 38282
rect 29920 38218 29972 38224
rect 30196 38276 30248 38282
rect 30196 38218 30248 38224
rect 29736 37800 29788 37806
rect 29736 37742 29788 37748
rect 29748 37641 29776 37742
rect 29932 37738 29960 38218
rect 30012 38208 30064 38214
rect 30064 38168 30144 38196
rect 30012 38150 30064 38156
rect 29920 37732 29972 37738
rect 29920 37674 29972 37680
rect 29828 37664 29880 37670
rect 29734 37632 29790 37641
rect 29828 37606 29880 37612
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 29734 37567 29790 37576
rect 29656 36094 29776 36122
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29656 35442 29684 35974
rect 29748 35834 29776 36094
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29840 35680 29868 37606
rect 30024 37262 30052 37606
rect 29920 37256 29972 37262
rect 29918 37224 29920 37233
rect 30012 37256 30064 37262
rect 29972 37224 29974 37233
rect 30012 37198 30064 37204
rect 29918 37159 29974 37168
rect 30010 37088 30066 37097
rect 30010 37023 30066 37032
rect 29920 35692 29972 35698
rect 29840 35652 29920 35680
rect 29920 35634 29972 35640
rect 30024 35601 30052 37023
rect 30116 36786 30144 38168
rect 30208 37806 30236 38218
rect 30196 37800 30248 37806
rect 30196 37742 30248 37748
rect 30300 37369 30328 39442
rect 30392 39001 30420 39986
rect 30378 38992 30434 39001
rect 30378 38927 30434 38936
rect 30484 38842 30512 41074
rect 31128 41070 31156 41386
rect 31116 41064 31168 41070
rect 31116 41006 31168 41012
rect 30656 40452 30708 40458
rect 30656 40394 30708 40400
rect 30564 39024 30616 39030
rect 30564 38966 30616 38972
rect 30392 38814 30512 38842
rect 30392 37942 30420 38814
rect 30576 38554 30604 38966
rect 30668 38962 30696 40394
rect 31024 40044 31076 40050
rect 31024 39986 31076 39992
rect 30840 39840 30892 39846
rect 30840 39782 30892 39788
rect 30852 38962 30880 39782
rect 31036 39098 31064 39986
rect 31024 39092 31076 39098
rect 31024 39034 31076 39040
rect 30656 38956 30708 38962
rect 30656 38898 30708 38904
rect 30840 38956 30892 38962
rect 30840 38898 30892 38904
rect 31128 38554 31156 41006
rect 31496 40526 31524 41754
rect 31588 41682 31616 42026
rect 31576 41676 31628 41682
rect 31576 41618 31628 41624
rect 31588 41414 31616 41618
rect 31588 41386 31708 41414
rect 31680 41138 31708 41386
rect 31668 41132 31720 41138
rect 31668 41074 31720 41080
rect 31576 40928 31628 40934
rect 31576 40870 31628 40876
rect 31588 40594 31616 40870
rect 31576 40588 31628 40594
rect 31576 40530 31628 40536
rect 31484 40520 31536 40526
rect 31484 40462 31536 40468
rect 31392 39976 31444 39982
rect 31392 39918 31444 39924
rect 31482 39944 31538 39953
rect 31404 38826 31432 39918
rect 31482 39879 31538 39888
rect 31392 38820 31444 38826
rect 31392 38762 31444 38768
rect 30564 38548 30616 38554
rect 30564 38490 30616 38496
rect 31116 38548 31168 38554
rect 31116 38490 31168 38496
rect 30840 38344 30892 38350
rect 30840 38286 30892 38292
rect 31024 38344 31076 38350
rect 31024 38286 31076 38292
rect 30564 38004 30616 38010
rect 30564 37946 30616 37952
rect 30748 38004 30800 38010
rect 30748 37946 30800 37952
rect 30380 37936 30432 37942
rect 30380 37878 30432 37884
rect 30286 37360 30342 37369
rect 30286 37295 30342 37304
rect 30300 37194 30328 37295
rect 30392 37194 30420 37878
rect 30472 37868 30524 37874
rect 30472 37810 30524 37816
rect 30288 37188 30340 37194
rect 30288 37130 30340 37136
rect 30380 37188 30432 37194
rect 30380 37130 30432 37136
rect 30208 36910 30420 36938
rect 30484 36922 30512 37810
rect 30576 37126 30604 37946
rect 30656 37868 30708 37874
rect 30656 37810 30708 37816
rect 30564 37120 30616 37126
rect 30564 37062 30616 37068
rect 30208 36786 30236 36910
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 30196 36780 30248 36786
rect 30196 36722 30248 36728
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30300 36145 30328 36722
rect 30392 36582 30420 36910
rect 30472 36916 30524 36922
rect 30472 36858 30524 36864
rect 30564 36916 30616 36922
rect 30564 36858 30616 36864
rect 30576 36718 30604 36858
rect 30564 36712 30616 36718
rect 30564 36654 30616 36660
rect 30380 36576 30432 36582
rect 30380 36518 30432 36524
rect 30286 36136 30342 36145
rect 30286 36071 30342 36080
rect 30392 36038 30420 36518
rect 30472 36372 30524 36378
rect 30472 36314 30524 36320
rect 30484 36174 30512 36314
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 30668 36106 30696 37810
rect 30656 36100 30708 36106
rect 30656 36042 30708 36048
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30104 35760 30156 35766
rect 30104 35702 30156 35708
rect 30194 35728 30250 35737
rect 30010 35592 30066 35601
rect 30010 35527 30066 35536
rect 30012 35488 30064 35494
rect 29656 35414 29776 35442
rect 30012 35430 30064 35436
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 29460 35012 29512 35018
rect 29460 34954 29512 34960
rect 29368 34604 29420 34610
rect 29368 34546 29420 34552
rect 29748 34542 29776 35414
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29736 34536 29788 34542
rect 29736 34478 29788 34484
rect 29288 34202 29316 34478
rect 29276 34196 29328 34202
rect 29276 34138 29328 34144
rect 29460 33992 29512 33998
rect 29458 33960 29460 33969
rect 29552 33992 29604 33998
rect 29512 33960 29514 33969
rect 29552 33934 29604 33940
rect 29458 33895 29514 33904
rect 29564 33590 29592 33934
rect 29552 33584 29604 33590
rect 29552 33526 29604 33532
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 29472 32910 29500 33254
rect 29460 32904 29512 32910
rect 29460 32846 29512 32852
rect 29276 32836 29328 32842
rect 29276 32778 29328 32784
rect 29288 32570 29316 32778
rect 29564 32570 29592 33526
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29276 32564 29328 32570
rect 29276 32506 29328 32512
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29196 32434 29316 32450
rect 29656 32434 29684 33458
rect 29748 33454 29776 34478
rect 29736 33448 29788 33454
rect 29736 33390 29788 33396
rect 29748 33318 29776 33390
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29196 32428 29328 32434
rect 29196 32422 29276 32428
rect 29276 32370 29328 32376
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29644 32292 29696 32298
rect 29644 32234 29696 32240
rect 28816 31952 28868 31958
rect 28816 31894 28868 31900
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28632 31408 28684 31414
rect 28632 31350 28684 31356
rect 28552 31232 28672 31260
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28460 30258 28488 30670
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28644 29578 28672 31232
rect 28828 30802 28856 31894
rect 28908 31816 28960 31822
rect 28906 31784 28908 31793
rect 28960 31784 28962 31793
rect 28906 31719 28962 31728
rect 29276 31680 29328 31686
rect 29276 31622 29328 31628
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 28920 30938 28948 31282
rect 28908 30932 28960 30938
rect 28908 30874 28960 30880
rect 28816 30796 28868 30802
rect 28816 30738 28868 30744
rect 28920 30598 28948 30874
rect 29000 30864 29052 30870
rect 29000 30806 29052 30812
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28814 30288 28870 30297
rect 28814 30223 28816 30232
rect 28868 30223 28870 30232
rect 28816 30194 28868 30200
rect 28920 30138 28948 30534
rect 28828 30110 28948 30138
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28540 29504 28592 29510
rect 28540 29446 28592 29452
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28368 28762 28396 29242
rect 28356 28756 28408 28762
rect 28356 28698 28408 28704
rect 28368 28506 28396 28698
rect 28080 28484 28132 28490
rect 28080 28426 28132 28432
rect 28276 28478 28396 28506
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27816 26790 27844 27542
rect 27908 27470 27936 27662
rect 27988 27668 28040 27674
rect 27988 27610 28040 27616
rect 28092 27470 28120 28426
rect 28276 28150 28304 28478
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28368 28218 28396 28358
rect 28356 28212 28408 28218
rect 28356 28154 28408 28160
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 27804 26784 27856 26790
rect 27804 26726 27856 26732
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27632 24954 27660 25230
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 23526 27660 23734
rect 27724 23662 27752 24142
rect 27816 23730 27844 26726
rect 27988 26444 28040 26450
rect 27988 26386 28040 26392
rect 28000 25906 28028 26386
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28000 25498 28028 25842
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 28000 25294 28028 25434
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28092 24682 28120 27406
rect 28552 27062 28580 29446
rect 28644 28422 28672 29514
rect 28828 28422 28856 30110
rect 29012 29170 29040 30806
rect 29104 30326 29132 31282
rect 29184 30592 29236 30598
rect 29184 30534 29236 30540
rect 29092 30320 29144 30326
rect 29092 30262 29144 30268
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 29196 28966 29224 30534
rect 29288 28966 29316 31622
rect 29552 31408 29604 31414
rect 29552 31350 29604 31356
rect 29368 30320 29420 30326
rect 29368 30262 29420 30268
rect 29184 28960 29236 28966
rect 29184 28902 29236 28908
rect 29276 28960 29328 28966
rect 29276 28902 29328 28908
rect 29380 28778 29408 30262
rect 29460 29232 29512 29238
rect 29460 29174 29512 29180
rect 29564 29186 29592 31350
rect 29656 30190 29684 32234
rect 29840 32026 29868 34954
rect 29932 34649 29960 35022
rect 29918 34640 29974 34649
rect 30024 34610 30052 35430
rect 30116 35222 30144 35702
rect 30194 35663 30196 35672
rect 30248 35663 30250 35672
rect 30300 35680 30328 35974
rect 30654 35864 30710 35873
rect 30654 35799 30710 35808
rect 30380 35692 30432 35698
rect 30300 35652 30380 35680
rect 30196 35634 30248 35640
rect 30380 35634 30432 35640
rect 30286 35592 30342 35601
rect 30286 35527 30342 35536
rect 30104 35216 30156 35222
rect 30104 35158 30156 35164
rect 30116 35086 30144 35158
rect 30300 35086 30328 35527
rect 30104 35080 30156 35086
rect 30104 35022 30156 35028
rect 30288 35080 30340 35086
rect 30288 35022 30340 35028
rect 29918 34575 29974 34584
rect 30012 34604 30064 34610
rect 29932 33046 29960 34575
rect 30012 34546 30064 34552
rect 30024 33862 30052 34546
rect 30562 34368 30618 34377
rect 30562 34303 30618 34312
rect 30104 34128 30156 34134
rect 30104 34070 30156 34076
rect 30116 33998 30144 34070
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30012 33856 30064 33862
rect 30012 33798 30064 33804
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30024 33522 30052 33798
rect 30484 33697 30512 33798
rect 30470 33688 30526 33697
rect 30470 33623 30526 33632
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 30104 33516 30156 33522
rect 30104 33458 30156 33464
rect 30288 33516 30340 33522
rect 30288 33458 30340 33464
rect 29920 33040 29972 33046
rect 29920 32982 29972 32988
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29828 32020 29880 32026
rect 29828 31962 29880 31968
rect 29932 31822 29960 32846
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 30024 32298 30052 32370
rect 30116 32298 30144 33458
rect 30300 32910 30328 33458
rect 30378 33144 30434 33153
rect 30378 33079 30380 33088
rect 30432 33079 30434 33088
rect 30380 33050 30432 33056
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 30196 32836 30248 32842
rect 30196 32778 30248 32784
rect 30012 32292 30064 32298
rect 30012 32234 30064 32240
rect 30104 32292 30156 32298
rect 30104 32234 30156 32240
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29920 31816 29972 31822
rect 29920 31758 29972 31764
rect 29932 31346 29960 31758
rect 29920 31340 29972 31346
rect 29840 31300 29920 31328
rect 29736 31136 29788 31142
rect 29734 31104 29736 31113
rect 29788 31104 29790 31113
rect 29734 31039 29790 31048
rect 29734 30968 29790 30977
rect 29734 30903 29736 30912
rect 29788 30903 29790 30912
rect 29736 30874 29788 30880
rect 29644 30184 29696 30190
rect 29840 30172 29868 31300
rect 29920 31282 29972 31288
rect 29920 31136 29972 31142
rect 30012 31136 30064 31142
rect 29920 31078 29972 31084
rect 30010 31104 30012 31113
rect 30064 31104 30066 31113
rect 29932 30734 29960 31078
rect 30010 31039 30066 31048
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 29920 30592 29972 30598
rect 29920 30534 29972 30540
rect 29932 30326 29960 30534
rect 29920 30320 29972 30326
rect 29920 30262 29972 30268
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 29840 30144 29960 30172
rect 29644 30126 29696 30132
rect 29656 29306 29684 30126
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29840 29646 29868 29990
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29104 28750 29408 28778
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28644 27334 28672 28358
rect 28724 28076 28776 28082
rect 28724 28018 28776 28024
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28540 27056 28592 27062
rect 28540 26998 28592 27004
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28448 26988 28500 26994
rect 28448 26930 28500 26936
rect 28184 25838 28212 26930
rect 28460 26450 28488 26930
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 28552 26042 28580 26998
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28172 25832 28224 25838
rect 28172 25774 28224 25780
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28184 24818 28212 25230
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28080 24676 28132 24682
rect 28080 24618 28132 24624
rect 28092 24206 28120 24618
rect 28184 24274 28212 24754
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28172 24268 28224 24274
rect 28172 24210 28224 24216
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 28276 24154 28304 24550
rect 28354 24168 28410 24177
rect 27908 23730 27936 24142
rect 28276 24126 28354 24154
rect 28354 24103 28410 24112
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 27632 22710 27660 23462
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27632 21146 27660 21422
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27434 20567 27436 20576
rect 27488 20567 27490 20576
rect 27528 20596 27580 20602
rect 27436 20538 27488 20544
rect 27528 20538 27580 20544
rect 27632 20466 27660 20878
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 17134 27200 18158
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 26976 16448 27028 16454
rect 26976 16390 27028 16396
rect 26896 16238 27016 16266
rect 26606 16215 26608 16224
rect 26660 16215 26662 16224
rect 26608 16186 26660 16192
rect 26988 14385 27016 16238
rect 26974 14376 27030 14385
rect 26792 14340 26844 14346
rect 26974 14311 27030 14320
rect 26792 14282 26844 14288
rect 26476 13892 26556 13920
rect 26424 13874 26476 13880
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 12986 26280 13738
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26436 12442 26464 13874
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26528 13394 26556 13670
rect 26804 13530 26832 14282
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 26160 11082 26188 11834
rect 26436 11218 26464 12378
rect 26620 12306 26648 12922
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 27172 11762 27200 17070
rect 27264 16046 27292 19654
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27264 15706 27292 15982
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 27356 15094 27384 20198
rect 27448 19854 27476 20402
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27448 17882 27476 18226
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27632 17814 27660 18362
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27448 16794 27476 17138
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27632 16250 27660 16526
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27344 15088 27396 15094
rect 27344 15030 27396 15036
rect 27356 14074 27384 15030
rect 27632 15026 27660 15302
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27344 14068 27396 14074
rect 27344 14010 27396 14016
rect 27448 13394 27476 14554
rect 27540 14006 27568 14758
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27632 13734 27660 14962
rect 27724 14618 27752 23598
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27816 22506 27844 23122
rect 28368 23118 28396 24103
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28172 22976 28224 22982
rect 28172 22918 28224 22924
rect 28184 22642 28212 22918
rect 28368 22778 28396 23054
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 27804 22500 27856 22506
rect 27804 22442 27856 22448
rect 28080 21956 28132 21962
rect 28080 21898 28132 21904
rect 28092 21690 28120 21898
rect 28080 21684 28132 21690
rect 28080 21626 28132 21632
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27816 17762 27844 19314
rect 27908 17882 27936 20334
rect 28000 19786 28028 20334
rect 27988 19780 28040 19786
rect 27988 19722 28040 19728
rect 28000 19514 28028 19722
rect 27988 19508 28040 19514
rect 27988 19450 28040 19456
rect 27896 17876 27948 17882
rect 27896 17818 27948 17824
rect 27986 17776 28042 17785
rect 27816 17734 27936 17762
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27816 16794 27844 17546
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27908 16561 27936 17734
rect 27986 17711 28042 17720
rect 28000 17678 28028 17711
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 27894 16552 27950 16561
rect 27894 16487 27950 16496
rect 27804 16108 27856 16114
rect 27908 16096 27936 16487
rect 27856 16068 27936 16096
rect 27804 16050 27856 16056
rect 27908 15706 27936 16068
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 28000 15366 28028 17478
rect 28092 15910 28120 21626
rect 28172 21412 28224 21418
rect 28172 21354 28224 21360
rect 28184 21146 28212 21354
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28368 20602 28396 20878
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28356 20256 28408 20262
rect 28356 20198 28408 20204
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28172 19780 28224 19786
rect 28172 19722 28224 19728
rect 28184 18086 28212 19722
rect 28276 19446 28304 19994
rect 28368 19514 28396 20198
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28264 19440 28316 19446
rect 28264 19382 28316 19388
rect 28368 18902 28396 19450
rect 28356 18896 28408 18902
rect 28356 18838 28408 18844
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28172 18080 28224 18086
rect 28172 18022 28224 18028
rect 28184 17542 28212 18022
rect 28368 17678 28396 18634
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 28368 17338 28396 17614
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 28092 15570 28120 15846
rect 28080 15564 28132 15570
rect 28080 15506 28132 15512
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27632 13258 27660 13670
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27356 12442 27384 12786
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27344 12436 27396 12442
rect 27344 12378 27396 12384
rect 27448 11830 27476 12582
rect 28460 12102 28488 25774
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28644 24410 28672 25230
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28632 23656 28684 23662
rect 28632 23598 28684 23604
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28552 21486 28580 21966
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28552 21146 28580 21422
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28552 18222 28580 19246
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28644 17796 28672 23598
rect 28736 21894 28764 28018
rect 28828 27402 28856 28358
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 28816 27396 28868 27402
rect 28816 27338 28868 27344
rect 29012 26246 29040 27814
rect 29104 26450 29132 28750
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29380 27674 29408 28018
rect 29368 27668 29420 27674
rect 29368 27610 29420 27616
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29196 27130 29224 27406
rect 29184 27124 29236 27130
rect 29472 27112 29500 29174
rect 29564 29158 29684 29186
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29564 27674 29592 28018
rect 29656 27878 29684 29158
rect 29748 29073 29776 29582
rect 29734 29064 29790 29073
rect 29734 28999 29790 29008
rect 29828 29028 29880 29034
rect 29644 27872 29696 27878
rect 29644 27814 29696 27820
rect 29552 27668 29604 27674
rect 29552 27610 29604 27616
rect 29184 27066 29236 27072
rect 29380 27084 29500 27112
rect 29380 26994 29408 27084
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29092 26444 29144 26450
rect 29092 26386 29144 26392
rect 29104 26314 29132 26386
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29092 26308 29144 26314
rect 29092 26250 29144 26256
rect 29184 26308 29236 26314
rect 29184 26250 29236 26256
rect 29000 26240 29052 26246
rect 29000 26182 29052 26188
rect 29092 25492 29144 25498
rect 29092 25434 29144 25440
rect 29000 25220 29052 25226
rect 29000 25162 29052 25168
rect 28816 25152 28868 25158
rect 28816 25094 28868 25100
rect 28828 24886 28856 25094
rect 28816 24880 28868 24886
rect 28816 24822 28868 24828
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28920 23322 28948 23666
rect 29012 23594 29040 25162
rect 29104 24886 29132 25434
rect 29196 25430 29224 26250
rect 29184 25424 29236 25430
rect 29184 25366 29236 25372
rect 29092 24880 29144 24886
rect 29092 24822 29144 24828
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 28920 23118 28948 23258
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28908 22976 28960 22982
rect 28908 22918 28960 22924
rect 28816 22500 28868 22506
rect 28816 22442 28868 22448
rect 28828 22001 28856 22442
rect 28920 22234 28948 22918
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 29000 22160 29052 22166
rect 28998 22128 29000 22137
rect 29052 22128 29054 22137
rect 28998 22063 29054 22072
rect 28814 21992 28870 22001
rect 28814 21927 28870 21936
rect 28908 21956 28960 21962
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28828 20942 28856 21927
rect 28908 21898 28960 21904
rect 28920 21690 28948 21898
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 29104 21010 29132 24822
rect 29196 24138 29224 25366
rect 29184 24132 29236 24138
rect 29184 24074 29236 24080
rect 29184 23792 29236 23798
rect 29184 23734 29236 23740
rect 29196 22094 29224 23734
rect 29288 22658 29316 26318
rect 29380 25226 29408 26930
rect 29472 25362 29500 26930
rect 29564 26586 29592 26930
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29460 25356 29512 25362
rect 29460 25298 29512 25304
rect 29368 25220 29420 25226
rect 29368 25162 29420 25168
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29380 22778 29408 24754
rect 29472 24682 29500 25298
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29460 24676 29512 24682
rect 29460 24618 29512 24624
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29472 23798 29500 24142
rect 29460 23792 29512 23798
rect 29460 23734 29512 23740
rect 29564 23526 29592 25230
rect 29644 25152 29696 25158
rect 29644 25094 29696 25100
rect 29552 23520 29604 23526
rect 29552 23462 29604 23468
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29288 22630 29500 22658
rect 29472 22094 29500 22630
rect 29196 22066 29408 22094
rect 29472 22066 29592 22094
rect 29380 21554 29408 22066
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 28816 20936 28868 20942
rect 28736 20896 28816 20924
rect 28736 20058 28764 20896
rect 28816 20878 28868 20884
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29104 20534 29132 20742
rect 29092 20528 29144 20534
rect 29092 20470 29144 20476
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 28724 20052 28776 20058
rect 28724 19994 28776 20000
rect 28828 19922 28856 20266
rect 28920 20262 28948 20402
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 28906 19952 28962 19961
rect 28816 19916 28868 19922
rect 28906 19887 28908 19896
rect 28816 19858 28868 19864
rect 28960 19887 28962 19896
rect 28908 19858 28960 19864
rect 28828 18834 28856 19858
rect 29184 19848 29236 19854
rect 29184 19790 29236 19796
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28920 18086 28948 19450
rect 29196 19378 29224 19790
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29380 19446 29408 19722
rect 29368 19440 29420 19446
rect 29368 19382 29420 19388
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 29012 18970 29040 19246
rect 29092 19168 29144 19174
rect 29092 19110 29144 19116
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29012 18358 29040 18906
rect 29104 18630 29132 19110
rect 29196 18766 29224 19314
rect 29380 18986 29408 19382
rect 29288 18958 29408 18986
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 28908 18080 28960 18086
rect 28908 18022 28960 18028
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28552 17768 28672 17796
rect 28552 17338 28580 17768
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28552 16658 28580 17274
rect 28644 16998 28672 17478
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28644 16590 28672 16934
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 28552 14414 28580 15438
rect 28736 15162 28764 17070
rect 28828 16454 28856 17818
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 28920 16590 28948 17478
rect 29092 17264 29144 17270
rect 29092 17206 29144 17212
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29012 16794 29040 17138
rect 29000 16788 29052 16794
rect 29000 16730 29052 16736
rect 29104 16658 29132 17206
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28816 16448 28868 16454
rect 28816 16390 28868 16396
rect 28828 15314 28856 16390
rect 28920 15502 28948 16526
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28828 15286 28948 15314
rect 28814 15192 28870 15201
rect 28724 15156 28776 15162
rect 28644 15116 28724 15144
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28644 14346 28672 15116
rect 28814 15127 28870 15136
rect 28724 15098 28776 15104
rect 28724 14816 28776 14822
rect 28724 14758 28776 14764
rect 28632 14340 28684 14346
rect 28632 14282 28684 14288
rect 28736 14090 28764 14758
rect 28828 14414 28856 15127
rect 28920 14906 28948 15286
rect 29104 15162 29132 16594
rect 29196 16522 29224 16934
rect 29184 16516 29236 16522
rect 29184 16458 29236 16464
rect 29196 16114 29224 16458
rect 29184 16108 29236 16114
rect 29184 16050 29236 16056
rect 29196 15201 29224 16050
rect 29182 15192 29238 15201
rect 29092 15156 29144 15162
rect 29182 15127 29238 15136
rect 29092 15098 29144 15104
rect 29288 15094 29316 18958
rect 29564 18850 29592 22066
rect 29380 18822 29592 18850
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 29012 14906 29040 14962
rect 28920 14878 29040 14906
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 28920 14550 28948 14878
rect 29104 14822 29132 14894
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29196 14618 29224 14962
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 29000 14544 29052 14550
rect 29000 14486 29052 14492
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28736 14062 28856 14090
rect 28828 12238 28856 14062
rect 29012 13938 29040 14486
rect 29288 13938 29316 15030
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29104 13530 29132 13874
rect 29184 13864 29236 13870
rect 29184 13806 29236 13812
rect 29196 13734 29224 13806
rect 29184 13728 29236 13734
rect 29184 13670 29236 13676
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28920 12374 28948 13262
rect 29196 12918 29224 13670
rect 29288 13462 29316 13874
rect 29276 13456 29328 13462
rect 29276 13398 29328 13404
rect 29184 12912 29236 12918
rect 29184 12854 29236 12860
rect 28908 12368 28960 12374
rect 28908 12310 28960 12316
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28460 11898 28488 12038
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 27436 11824 27488 11830
rect 27436 11766 27488 11772
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27172 11218 27200 11698
rect 27540 11286 27568 11766
rect 29380 11762 29408 18822
rect 29460 18760 29512 18766
rect 29460 18702 29512 18708
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29472 17814 29500 18702
rect 29564 18222 29592 18702
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29564 17134 29592 18158
rect 29552 17128 29604 17134
rect 29552 17070 29604 17076
rect 29564 16046 29592 17070
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29564 14226 29592 15982
rect 29472 14198 29592 14226
rect 29472 13734 29500 14198
rect 29656 14006 29684 25094
rect 29748 24818 29776 28999
rect 29828 28970 29880 28976
rect 29840 27062 29868 28970
rect 29932 27946 29960 30144
rect 30024 29306 30052 30194
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30116 28490 30144 31826
rect 30208 31822 30236 32778
rect 30300 32434 30328 32846
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30288 32428 30340 32434
rect 30288 32370 30340 32376
rect 30392 32366 30420 32506
rect 30484 32502 30512 33623
rect 30576 32910 30604 34303
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 30472 32496 30524 32502
rect 30472 32438 30524 32444
rect 30380 32360 30432 32366
rect 30300 32308 30380 32314
rect 30300 32302 30432 32308
rect 30300 32286 30420 32302
rect 30300 32026 30328 32286
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30208 31396 30236 31758
rect 30288 31408 30340 31414
rect 30208 31368 30288 31396
rect 30288 31350 30340 31356
rect 30196 30864 30248 30870
rect 30196 30806 30248 30812
rect 30104 28484 30156 28490
rect 30104 28426 30156 28432
rect 29920 27940 29972 27946
rect 29920 27882 29972 27888
rect 29918 27568 29974 27577
rect 29918 27503 29974 27512
rect 29828 27056 29880 27062
rect 29828 26998 29880 27004
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29748 24274 29776 24550
rect 29736 24268 29788 24274
rect 29736 24210 29788 24216
rect 29736 22160 29788 22166
rect 29736 22102 29788 22108
rect 29748 21622 29776 22102
rect 29840 21690 29868 26862
rect 29932 26382 29960 27503
rect 30208 27402 30236 30806
rect 30300 30666 30328 31350
rect 30392 31210 30420 32166
rect 30380 31204 30432 31210
rect 30380 31146 30432 31152
rect 30288 30660 30340 30666
rect 30288 30602 30340 30608
rect 30668 30598 30696 35799
rect 30760 35290 30788 37946
rect 30852 37210 30880 38286
rect 31036 37466 31064 38286
rect 31208 37664 31260 37670
rect 31208 37606 31260 37612
rect 31024 37460 31076 37466
rect 31024 37402 31076 37408
rect 31024 37324 31076 37330
rect 31024 37266 31076 37272
rect 30932 37256 30984 37262
rect 30852 37204 30932 37210
rect 30852 37198 30984 37204
rect 30852 37182 30972 37198
rect 30852 36378 30880 37182
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30840 36372 30892 36378
rect 30840 36314 30892 36320
rect 30852 36106 30880 36314
rect 30840 36100 30892 36106
rect 30840 36042 30892 36048
rect 30840 35828 30892 35834
rect 30840 35770 30892 35776
rect 30748 35284 30800 35290
rect 30748 35226 30800 35232
rect 30852 34678 30880 35770
rect 30840 34672 30892 34678
rect 30840 34614 30892 34620
rect 30840 34400 30892 34406
rect 30840 34342 30892 34348
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30760 33590 30788 34138
rect 30748 33584 30800 33590
rect 30748 33526 30800 33532
rect 30746 33416 30802 33425
rect 30746 33351 30802 33360
rect 30760 32910 30788 33351
rect 30748 32904 30800 32910
rect 30748 32846 30800 32852
rect 30748 30796 30800 30802
rect 30748 30738 30800 30744
rect 30656 30592 30708 30598
rect 30656 30534 30708 30540
rect 30760 30326 30788 30738
rect 30748 30320 30800 30326
rect 30852 30308 30880 34342
rect 30944 33862 30972 36722
rect 31036 35494 31064 37266
rect 31220 36786 31248 37606
rect 31208 36780 31260 36786
rect 31208 36722 31260 36728
rect 31208 36576 31260 36582
rect 31208 36518 31260 36524
rect 31116 36032 31168 36038
rect 31116 35974 31168 35980
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30932 33856 30984 33862
rect 31128 33810 31156 35974
rect 31220 35562 31248 36518
rect 31404 36378 31432 38762
rect 31496 37874 31524 39879
rect 31576 39840 31628 39846
rect 31576 39782 31628 39788
rect 31588 39438 31616 39782
rect 31680 39438 31708 41074
rect 31772 40458 31800 44066
rect 32312 42220 32364 42226
rect 32312 42162 32364 42168
rect 31852 41472 31904 41478
rect 31852 41414 31904 41420
rect 31864 41206 31892 41414
rect 31852 41200 31904 41206
rect 31852 41142 31904 41148
rect 32324 40730 32352 42162
rect 32600 42106 32628 44200
rect 34164 44130 34192 44200
rect 35728 44146 35756 44200
rect 34152 44124 34204 44130
rect 34152 44066 34204 44072
rect 34612 44124 34664 44130
rect 35728 44118 35940 44146
rect 34612 44066 34664 44072
rect 34336 42152 34388 42158
rect 32600 42078 32720 42106
rect 34336 42094 34388 42100
rect 32588 42016 32640 42022
rect 32588 41958 32640 41964
rect 32496 41472 32548 41478
rect 32496 41414 32548 41420
rect 32312 40724 32364 40730
rect 32312 40666 32364 40672
rect 31760 40452 31812 40458
rect 31760 40394 31812 40400
rect 31852 40112 31904 40118
rect 31852 40054 31904 40060
rect 31760 40044 31812 40050
rect 31760 39986 31812 39992
rect 31772 39506 31800 39986
rect 31760 39500 31812 39506
rect 31760 39442 31812 39448
rect 31576 39432 31628 39438
rect 31576 39374 31628 39380
rect 31668 39432 31720 39438
rect 31668 39374 31720 39380
rect 31574 38312 31630 38321
rect 31574 38247 31576 38256
rect 31628 38247 31630 38256
rect 31576 38218 31628 38224
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 31496 37466 31524 37810
rect 31484 37460 31536 37466
rect 31484 37402 31536 37408
rect 31680 37233 31708 39374
rect 31772 39098 31800 39442
rect 31760 39092 31812 39098
rect 31760 39034 31812 39040
rect 31760 38820 31812 38826
rect 31760 38762 31812 38768
rect 31772 38010 31800 38762
rect 31760 38004 31812 38010
rect 31760 37946 31812 37952
rect 31760 37392 31812 37398
rect 31760 37334 31812 37340
rect 31666 37224 31722 37233
rect 31666 37159 31722 37168
rect 31576 36780 31628 36786
rect 31576 36722 31628 36728
rect 31392 36372 31444 36378
rect 31392 36314 31444 36320
rect 31484 36168 31536 36174
rect 31484 36110 31536 36116
rect 31496 35562 31524 36110
rect 31208 35556 31260 35562
rect 31208 35498 31260 35504
rect 31484 35556 31536 35562
rect 31484 35498 31536 35504
rect 31220 35018 31248 35498
rect 31392 35080 31444 35086
rect 31392 35022 31444 35028
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 30932 33798 30984 33804
rect 31036 33782 31340 33810
rect 31036 33590 31064 33782
rect 31312 33658 31340 33782
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 31300 33652 31352 33658
rect 31300 33594 31352 33600
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 31220 33454 31248 33594
rect 31208 33448 31260 33454
rect 31208 33390 31260 33396
rect 31024 33380 31076 33386
rect 31024 33322 31076 33328
rect 30932 33312 30984 33318
rect 30932 33254 30984 33260
rect 30944 33114 30972 33254
rect 30932 33108 30984 33114
rect 30932 33050 30984 33056
rect 30932 32360 30984 32366
rect 30932 32302 30984 32308
rect 30944 31346 30972 32302
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 30944 30938 30972 31282
rect 30932 30932 30984 30938
rect 30932 30874 30984 30880
rect 30944 30734 30972 30874
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 30852 30280 30972 30308
rect 30748 30262 30800 30268
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30668 29238 30696 30194
rect 30656 29232 30708 29238
rect 30656 29174 30708 29180
rect 30944 29170 30972 30280
rect 31036 29782 31064 33322
rect 31116 33312 31168 33318
rect 31116 33254 31168 33260
rect 31128 33017 31156 33254
rect 31114 33008 31170 33017
rect 31114 32943 31170 32952
rect 31208 32768 31260 32774
rect 31208 32710 31260 32716
rect 31220 32609 31248 32710
rect 31206 32600 31262 32609
rect 31206 32535 31262 32544
rect 31220 30326 31248 32535
rect 31208 30320 31260 30326
rect 31208 30262 31260 30268
rect 31208 30184 31260 30190
rect 31206 30152 31208 30161
rect 31260 30152 31262 30161
rect 31206 30087 31262 30096
rect 31024 29776 31076 29782
rect 31024 29718 31076 29724
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30300 28762 30328 29106
rect 30288 28756 30340 28762
rect 30288 28698 30340 28704
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30840 28620 30892 28626
rect 30840 28562 30892 28568
rect 30564 28416 30616 28422
rect 30286 28384 30342 28393
rect 30564 28358 30616 28364
rect 30286 28319 30342 28328
rect 30300 27878 30328 28319
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30288 27464 30340 27470
rect 30288 27406 30340 27412
rect 30196 27396 30248 27402
rect 30196 27338 30248 27344
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 29932 24410 29960 24754
rect 29920 24404 29972 24410
rect 29920 24346 29972 24352
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29734 20632 29790 20641
rect 29734 20567 29790 20576
rect 29748 17202 29776 20567
rect 30024 19310 30052 25910
rect 30300 25498 30328 27406
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30392 27130 30420 27270
rect 30380 27124 30432 27130
rect 30380 27066 30432 27072
rect 30576 26586 30604 28358
rect 30564 26580 30616 26586
rect 30564 26522 30616 26528
rect 30654 26344 30710 26353
rect 30654 26279 30656 26288
rect 30708 26279 30710 26288
rect 30656 26250 30708 26256
rect 30760 25498 30788 28562
rect 30852 28218 30880 28562
rect 30840 28212 30892 28218
rect 30840 28154 30892 28160
rect 30944 28098 30972 29106
rect 31036 28558 31064 29718
rect 31208 29572 31260 29578
rect 31208 29514 31260 29520
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 31128 29306 31156 29446
rect 31220 29306 31248 29514
rect 31116 29300 31168 29306
rect 31116 29242 31168 29248
rect 31208 29300 31260 29306
rect 31208 29242 31260 29248
rect 31404 28762 31432 35022
rect 31484 33992 31536 33998
rect 31484 33934 31536 33940
rect 31496 33318 31524 33934
rect 31484 33312 31536 33318
rect 31484 33254 31536 33260
rect 31588 31346 31616 36722
rect 31772 35873 31800 37334
rect 31864 37126 31892 40054
rect 32404 39908 32456 39914
rect 32404 39850 32456 39856
rect 32416 38457 32444 39850
rect 32402 38448 32458 38457
rect 32312 38412 32364 38418
rect 32402 38383 32458 38392
rect 32312 38354 32364 38360
rect 32220 38276 32272 38282
rect 32220 38218 32272 38224
rect 32232 37738 32260 38218
rect 32324 38010 32352 38354
rect 32312 38004 32364 38010
rect 32312 37946 32364 37952
rect 32404 37936 32456 37942
rect 32508 37913 32536 41414
rect 32600 41138 32628 41958
rect 32588 41132 32640 41138
rect 32588 41074 32640 41080
rect 32692 40050 32720 42078
rect 33600 42016 33652 42022
rect 33600 41958 33652 41964
rect 34244 42016 34296 42022
rect 34244 41958 34296 41964
rect 33508 41540 33560 41546
rect 33508 41482 33560 41488
rect 32864 41268 32916 41274
rect 32864 41210 32916 41216
rect 32876 40526 32904 41210
rect 33520 41070 33548 41482
rect 33508 41064 33560 41070
rect 33508 41006 33560 41012
rect 32864 40520 32916 40526
rect 32864 40462 32916 40468
rect 32772 40452 32824 40458
rect 32772 40394 32824 40400
rect 32680 40044 32732 40050
rect 32680 39986 32732 39992
rect 32588 39364 32640 39370
rect 32588 39306 32640 39312
rect 32600 39098 32628 39306
rect 32588 39092 32640 39098
rect 32588 39034 32640 39040
rect 32600 38842 32628 39034
rect 32692 39030 32720 39986
rect 32680 39024 32732 39030
rect 32680 38966 32732 38972
rect 32600 38814 32720 38842
rect 32404 37878 32456 37884
rect 32494 37904 32550 37913
rect 32220 37732 32272 37738
rect 32272 37692 32352 37720
rect 32220 37674 32272 37680
rect 32220 37460 32272 37466
rect 32220 37402 32272 37408
rect 32034 37360 32090 37369
rect 32034 37295 32090 37304
rect 32048 37262 32076 37295
rect 32036 37256 32088 37262
rect 32036 37198 32088 37204
rect 31852 37120 31904 37126
rect 31852 37062 31904 37068
rect 31942 36952 31998 36961
rect 31942 36887 31998 36896
rect 31758 35864 31814 35873
rect 31668 35828 31720 35834
rect 31956 35850 31984 36887
rect 32048 36009 32076 37198
rect 32128 37188 32180 37194
rect 32128 37130 32180 37136
rect 32140 36922 32168 37130
rect 32128 36916 32180 36922
rect 32128 36858 32180 36864
rect 32034 36000 32090 36009
rect 32034 35935 32090 35944
rect 31956 35822 32076 35850
rect 32140 35834 32168 36858
rect 31758 35799 31814 35808
rect 31668 35770 31720 35776
rect 31680 35086 31708 35770
rect 31760 35692 31812 35698
rect 31760 35634 31812 35640
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31680 34746 31708 35022
rect 31772 34746 31800 35634
rect 31944 35624 31996 35630
rect 31944 35566 31996 35572
rect 31852 35216 31904 35222
rect 31852 35158 31904 35164
rect 31668 34740 31720 34746
rect 31668 34682 31720 34688
rect 31760 34740 31812 34746
rect 31760 34682 31812 34688
rect 31864 33998 31892 35158
rect 31852 33992 31904 33998
rect 31852 33934 31904 33940
rect 31956 33844 31984 35566
rect 31864 33816 31984 33844
rect 31760 33584 31812 33590
rect 31760 33526 31812 33532
rect 31772 33046 31800 33526
rect 31760 33040 31812 33046
rect 31760 32982 31812 32988
rect 31864 31498 31892 33816
rect 32048 32910 32076 35822
rect 32128 35828 32180 35834
rect 32128 35770 32180 35776
rect 32128 35692 32180 35698
rect 32128 35634 32180 35640
rect 32140 35222 32168 35634
rect 32128 35216 32180 35222
rect 32128 35158 32180 35164
rect 32232 35068 32260 37402
rect 32324 36802 32352 37692
rect 32416 37126 32444 37878
rect 32494 37839 32550 37848
rect 32588 37868 32640 37874
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 32324 36774 32444 36802
rect 32508 36786 32536 37839
rect 32588 37810 32640 37816
rect 32600 37398 32628 37810
rect 32588 37392 32640 37398
rect 32588 37334 32640 37340
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 32312 36712 32364 36718
rect 32312 36654 32364 36660
rect 32140 35057 32260 35068
rect 32140 35048 32274 35057
rect 32140 35040 32218 35048
rect 31944 32904 31996 32910
rect 31944 32846 31996 32852
rect 32036 32904 32088 32910
rect 32036 32846 32088 32852
rect 31956 32756 31984 32846
rect 31956 32728 32076 32756
rect 32048 32570 32076 32728
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 32036 32564 32088 32570
rect 32036 32506 32088 32512
rect 31956 31958 31984 32506
rect 32140 32502 32168 35040
rect 32218 34983 32274 34992
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 32232 34202 32260 34478
rect 32220 34196 32272 34202
rect 32220 34138 32272 34144
rect 32324 32910 32352 36654
rect 32416 35630 32444 36774
rect 32496 36780 32548 36786
rect 32496 36722 32548 36728
rect 32404 35624 32456 35630
rect 32404 35566 32456 35572
rect 32404 35488 32456 35494
rect 32404 35430 32456 35436
rect 32496 35488 32548 35494
rect 32496 35430 32548 35436
rect 32416 35222 32444 35430
rect 32404 35216 32456 35222
rect 32404 35158 32456 35164
rect 32416 33658 32444 35158
rect 32508 34785 32536 35430
rect 32600 35086 32628 37198
rect 32692 36786 32720 38814
rect 32784 38554 32812 40394
rect 32876 39438 32904 40462
rect 33140 40452 33192 40458
rect 33140 40394 33192 40400
rect 32864 39432 32916 39438
rect 32864 39374 32916 39380
rect 32876 38826 32904 39374
rect 33152 38978 33180 40394
rect 33232 40384 33284 40390
rect 33232 40326 33284 40332
rect 33244 40050 33272 40326
rect 33232 40044 33284 40050
rect 33232 39986 33284 39992
rect 33520 39982 33548 41006
rect 33508 39976 33560 39982
rect 33508 39918 33560 39924
rect 33612 39302 33640 41958
rect 33876 41540 33928 41546
rect 33876 41482 33928 41488
rect 33888 41002 33916 41482
rect 33876 40996 33928 41002
rect 33876 40938 33928 40944
rect 34060 40996 34112 41002
rect 34060 40938 34112 40944
rect 34072 40526 34100 40938
rect 34256 40730 34284 41958
rect 34244 40724 34296 40730
rect 34244 40666 34296 40672
rect 34060 40520 34112 40526
rect 34060 40462 34112 40468
rect 33968 40452 34020 40458
rect 33968 40394 34020 40400
rect 33980 40186 34008 40394
rect 33968 40180 34020 40186
rect 33968 40122 34020 40128
rect 33784 40044 33836 40050
rect 33784 39986 33836 39992
rect 33692 39568 33744 39574
rect 33692 39510 33744 39516
rect 33704 39409 33732 39510
rect 33690 39400 33746 39409
rect 33690 39335 33746 39344
rect 33232 39296 33284 39302
rect 33230 39264 33232 39273
rect 33324 39296 33376 39302
rect 33284 39264 33286 39273
rect 33324 39238 33376 39244
rect 33600 39296 33652 39302
rect 33600 39238 33652 39244
rect 33230 39199 33286 39208
rect 33060 38950 33180 38978
rect 32954 38856 33010 38865
rect 32864 38820 32916 38826
rect 32954 38791 33010 38800
rect 32864 38762 32916 38768
rect 32772 38548 32824 38554
rect 32772 38490 32824 38496
rect 32772 38412 32824 38418
rect 32772 38354 32824 38360
rect 32784 37874 32812 38354
rect 32772 37868 32824 37874
rect 32772 37810 32824 37816
rect 32864 37868 32916 37874
rect 32864 37810 32916 37816
rect 32876 36922 32904 37810
rect 32864 36916 32916 36922
rect 32864 36858 32916 36864
rect 32770 36816 32826 36825
rect 32680 36780 32732 36786
rect 32770 36751 32772 36760
rect 32680 36722 32732 36728
rect 32824 36751 32826 36760
rect 32772 36722 32824 36728
rect 32692 36378 32720 36722
rect 32680 36372 32732 36378
rect 32680 36314 32732 36320
rect 32784 36281 32812 36722
rect 32770 36272 32826 36281
rect 32770 36207 32826 36216
rect 32968 35698 32996 38791
rect 33060 38282 33088 38950
rect 33232 38888 33284 38894
rect 33232 38830 33284 38836
rect 33140 38820 33192 38826
rect 33140 38762 33192 38768
rect 33048 38276 33100 38282
rect 33048 38218 33100 38224
rect 33060 37330 33088 38218
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 33046 37224 33102 37233
rect 33046 37159 33102 37168
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32588 35080 32640 35086
rect 32588 35022 32640 35028
rect 32680 35080 32732 35086
rect 32680 35022 32732 35028
rect 32494 34776 32550 34785
rect 32494 34711 32550 34720
rect 32494 34640 32550 34649
rect 32494 34575 32550 34584
rect 32508 34202 32536 34575
rect 32692 34474 32720 35022
rect 32772 35012 32824 35018
rect 32772 34954 32824 34960
rect 32784 34610 32812 34954
rect 32772 34604 32824 34610
rect 32772 34546 32824 34552
rect 33060 34542 33088 37159
rect 33152 36718 33180 38762
rect 33244 38486 33272 38830
rect 33232 38480 33284 38486
rect 33232 38422 33284 38428
rect 33244 38282 33272 38422
rect 33336 38350 33364 39238
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 33612 38865 33640 38898
rect 33598 38856 33654 38865
rect 33598 38791 33654 38800
rect 33324 38344 33376 38350
rect 33324 38286 33376 38292
rect 33416 38344 33468 38350
rect 33416 38286 33468 38292
rect 33232 38276 33284 38282
rect 33232 38218 33284 38224
rect 33232 37188 33284 37194
rect 33232 37130 33284 37136
rect 33244 36922 33272 37130
rect 33232 36916 33284 36922
rect 33232 36858 33284 36864
rect 33140 36712 33192 36718
rect 33140 36654 33192 36660
rect 33140 35760 33192 35766
rect 33140 35702 33192 35708
rect 33152 35154 33180 35702
rect 33140 35148 33192 35154
rect 33140 35090 33192 35096
rect 33048 34536 33100 34542
rect 33048 34478 33100 34484
rect 32680 34468 32732 34474
rect 32680 34410 32732 34416
rect 32496 34196 32548 34202
rect 32496 34138 32548 34144
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32402 33008 32458 33017
rect 32402 32943 32458 32952
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32128 32496 32180 32502
rect 32128 32438 32180 32444
rect 32036 32428 32088 32434
rect 32036 32370 32088 32376
rect 32048 32065 32076 32370
rect 32140 32337 32168 32438
rect 32126 32328 32182 32337
rect 32126 32263 32182 32272
rect 32034 32056 32090 32065
rect 32034 31991 32090 32000
rect 31944 31952 31996 31958
rect 31944 31894 31996 31900
rect 32232 31906 32260 32846
rect 32416 32842 32444 32943
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32404 32564 32456 32570
rect 32404 32506 32456 32512
rect 32416 32434 32444 32506
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32312 32224 32364 32230
rect 32312 32166 32364 32172
rect 32404 32224 32456 32230
rect 32404 32166 32456 32172
rect 32324 32026 32352 32166
rect 32312 32020 32364 32026
rect 32312 31962 32364 31968
rect 32232 31878 32352 31906
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 32220 31816 32272 31822
rect 32220 31758 32272 31764
rect 31772 31470 31892 31498
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 31772 31278 31800 31470
rect 31850 31376 31906 31385
rect 31850 31311 31852 31320
rect 31904 31311 31906 31320
rect 31852 31282 31904 31288
rect 31760 31272 31812 31278
rect 31760 31214 31812 31220
rect 31772 29102 31800 31214
rect 31864 30802 31892 31282
rect 31852 30796 31904 30802
rect 31852 30738 31904 30744
rect 31944 30592 31996 30598
rect 31942 30560 31944 30569
rect 31996 30560 31998 30569
rect 31942 30495 31998 30504
rect 31852 30388 31904 30394
rect 31852 30330 31904 30336
rect 31668 29096 31720 29102
rect 31668 29038 31720 29044
rect 31760 29096 31812 29102
rect 31760 29038 31812 29044
rect 31576 28960 31628 28966
rect 31576 28902 31628 28908
rect 31392 28756 31444 28762
rect 31392 28698 31444 28704
rect 31588 28694 31616 28902
rect 31484 28688 31536 28694
rect 31484 28630 31536 28636
rect 31576 28688 31628 28694
rect 31576 28630 31628 28636
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 31208 28416 31260 28422
rect 31208 28358 31260 28364
rect 30852 28070 30972 28098
rect 31220 28082 31248 28358
rect 31496 28121 31524 28630
rect 31576 28484 31628 28490
rect 31576 28426 31628 28432
rect 31482 28112 31538 28121
rect 31208 28076 31260 28082
rect 30852 27130 30880 28070
rect 31208 28018 31260 28024
rect 31392 28076 31444 28082
rect 31482 28047 31538 28056
rect 31392 28018 31444 28024
rect 31404 27878 31432 28018
rect 31392 27872 31444 27878
rect 31392 27814 31444 27820
rect 31392 27532 31444 27538
rect 31392 27474 31444 27480
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30288 25492 30340 25498
rect 30288 25434 30340 25440
rect 30748 25492 30800 25498
rect 30748 25434 30800 25440
rect 30380 25356 30432 25362
rect 30380 25298 30432 25304
rect 30392 24886 30420 25298
rect 30852 25294 30880 27066
rect 31404 27062 31432 27474
rect 31392 27056 31444 27062
rect 31392 26998 31444 27004
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30380 24880 30432 24886
rect 30380 24822 30432 24828
rect 30104 24812 30156 24818
rect 30104 24754 30156 24760
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30116 23798 30144 24754
rect 30748 24608 30800 24614
rect 30748 24550 30800 24556
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30208 23798 30236 24142
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 30300 23866 30328 24006
rect 30760 23866 30788 24550
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30748 23860 30800 23866
rect 30748 23802 30800 23808
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 30196 23792 30248 23798
rect 30196 23734 30248 23740
rect 30208 23066 30236 23734
rect 30852 23730 30880 24754
rect 30944 24274 30972 26386
rect 31024 26240 31076 26246
rect 31024 26182 31076 26188
rect 31036 26042 31064 26182
rect 31024 26036 31076 26042
rect 31024 25978 31076 25984
rect 31300 26036 31352 26042
rect 31300 25978 31352 25984
rect 31312 25362 31340 25978
rect 31404 25770 31432 26998
rect 31496 26586 31524 28047
rect 31588 26976 31616 28426
rect 31680 27606 31708 29038
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31668 26988 31720 26994
rect 31588 26948 31668 26976
rect 31668 26930 31720 26936
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 31392 25764 31444 25770
rect 31392 25706 31444 25712
rect 31300 25356 31352 25362
rect 31300 25298 31352 25304
rect 31404 25294 31432 25706
rect 31496 25498 31524 25774
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31576 24948 31628 24954
rect 31576 24890 31628 24896
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 30932 24268 30984 24274
rect 30932 24210 30984 24216
rect 31300 24200 31352 24206
rect 31300 24142 31352 24148
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30840 23724 30892 23730
rect 30840 23666 30892 23672
rect 31208 23724 31260 23730
rect 31208 23666 31260 23672
rect 30288 23656 30340 23662
rect 30288 23598 30340 23604
rect 30116 23038 30236 23066
rect 30300 23050 30328 23598
rect 30288 23044 30340 23050
rect 30116 22710 30144 23038
rect 30288 22986 30340 22992
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30104 22704 30156 22710
rect 30104 22646 30156 22652
rect 30104 22092 30156 22098
rect 30104 22034 30156 22040
rect 30116 21690 30144 22034
rect 30208 21962 30236 22918
rect 30300 22778 30328 22986
rect 30392 22778 30420 23666
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30380 22772 30432 22778
rect 30380 22714 30432 22720
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30484 22438 30512 22714
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 30760 22234 30788 22578
rect 30748 22228 30800 22234
rect 30748 22170 30800 22176
rect 30196 21956 30248 21962
rect 30196 21898 30248 21904
rect 30104 21684 30156 21690
rect 30104 21626 30156 21632
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30116 20058 30144 20198
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 30116 19446 30144 19994
rect 30104 19440 30156 19446
rect 30104 19382 30156 19388
rect 30012 19304 30064 19310
rect 30012 19246 30064 19252
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29932 17882 29960 18226
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 30208 16794 30236 21898
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 30392 20058 30420 20810
rect 30576 20602 30604 21490
rect 30852 21418 30880 23666
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31024 22568 31076 22574
rect 31024 22510 31076 22516
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30840 21412 30892 21418
rect 30840 21354 30892 21360
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30748 20392 30800 20398
rect 30852 20380 30880 21354
rect 30800 20352 30880 20380
rect 30748 20334 30800 20340
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30852 19854 30880 20352
rect 30840 19848 30892 19854
rect 30840 19790 30892 19796
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 17678 30420 19314
rect 30748 18352 30800 18358
rect 30748 18294 30800 18300
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30668 17746 30696 18022
rect 30656 17740 30708 17746
rect 30656 17682 30708 17688
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30392 16794 30420 17614
rect 30760 17270 30788 18294
rect 30944 18086 30972 21966
rect 31036 21554 31064 22510
rect 31128 22030 31156 23598
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 31036 20806 31064 21490
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 31036 20262 31064 20742
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31024 20256 31076 20262
rect 31024 20198 31076 20204
rect 31128 19922 31156 20402
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 31036 18698 31064 19790
rect 31220 18970 31248 23666
rect 31312 23254 31340 24142
rect 31404 24138 31432 24754
rect 31588 24274 31616 24890
rect 31680 24614 31708 26930
rect 31772 25906 31800 29038
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31772 24954 31800 25842
rect 31760 24948 31812 24954
rect 31760 24890 31812 24896
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 31484 24268 31536 24274
rect 31484 24210 31536 24216
rect 31576 24268 31628 24274
rect 31576 24210 31628 24216
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31404 23322 31432 24074
rect 31392 23316 31444 23322
rect 31392 23258 31444 23264
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 31312 22710 31340 23190
rect 31300 22704 31352 22710
rect 31300 22646 31352 22652
rect 31390 21992 31446 22001
rect 31390 21927 31446 21936
rect 31404 21894 31432 21927
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31404 20262 31432 21830
rect 31496 21078 31524 24210
rect 31864 23798 31892 30330
rect 32048 30326 32076 31758
rect 32036 30320 32088 30326
rect 32036 30262 32088 30268
rect 31944 30184 31996 30190
rect 31944 30126 31996 30132
rect 31956 29510 31984 30126
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31956 29102 31984 29446
rect 32232 29306 32260 31758
rect 32324 31226 32352 31878
rect 32416 31414 32444 32166
rect 32508 31686 32536 34138
rect 32588 33992 32640 33998
rect 32692 33980 32720 34410
rect 32864 34196 32916 34202
rect 32864 34138 32916 34144
rect 32876 33998 32904 34138
rect 32640 33952 32720 33980
rect 32864 33992 32916 33998
rect 32588 33934 32640 33940
rect 32864 33934 32916 33940
rect 32600 33454 32628 33934
rect 32956 33924 33008 33930
rect 32956 33866 33008 33872
rect 32772 33516 32824 33522
rect 32692 33476 32772 33504
rect 32588 33448 32640 33454
rect 32588 33390 32640 33396
rect 32692 33318 32720 33476
rect 32772 33458 32824 33464
rect 32864 33448 32916 33454
rect 32784 33396 32864 33402
rect 32784 33390 32916 33396
rect 32784 33374 32904 33390
rect 32680 33312 32732 33318
rect 32600 33272 32680 33300
rect 32496 31680 32548 31686
rect 32496 31622 32548 31628
rect 32404 31408 32456 31414
rect 32404 31350 32456 31356
rect 32508 31346 32536 31622
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32324 31198 32444 31226
rect 32312 31136 32364 31142
rect 32312 31078 32364 31084
rect 32324 30734 32352 31078
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32416 30394 32444 31198
rect 32600 30734 32628 33272
rect 32680 33254 32732 33260
rect 32680 32904 32732 32910
rect 32680 32846 32732 32852
rect 32692 31822 32720 32846
rect 32784 32230 32812 33374
rect 32968 33318 32996 33866
rect 32956 33312 33008 33318
rect 32956 33254 33008 33260
rect 32968 33046 32996 33254
rect 32956 33040 33008 33046
rect 32862 33008 32918 33017
rect 32956 32982 33008 32988
rect 32862 32943 32918 32952
rect 32876 32434 32904 32943
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32772 32224 32824 32230
rect 32772 32166 32824 32172
rect 32772 32020 32824 32026
rect 32772 31962 32824 31968
rect 32784 31822 32812 31962
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32784 31142 32812 31758
rect 32864 31340 32916 31346
rect 32864 31282 32916 31288
rect 32772 31136 32824 31142
rect 32772 31078 32824 31084
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32772 30728 32824 30734
rect 32772 30670 32824 30676
rect 32404 30388 32456 30394
rect 32404 30330 32456 30336
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32496 29164 32548 29170
rect 32496 29106 32548 29112
rect 31944 29096 31996 29102
rect 31944 29038 31996 29044
rect 32508 28150 32536 29106
rect 32496 28144 32548 28150
rect 32496 28086 32548 28092
rect 32128 27940 32180 27946
rect 32128 27882 32180 27888
rect 32312 27940 32364 27946
rect 32312 27882 32364 27888
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 31956 27062 31984 27474
rect 32140 27402 32168 27882
rect 32324 27470 32352 27882
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 32036 27396 32088 27402
rect 32036 27338 32088 27344
rect 32128 27396 32180 27402
rect 32128 27338 32180 27344
rect 31944 27056 31996 27062
rect 31944 26998 31996 27004
rect 31944 26036 31996 26042
rect 31944 25978 31996 25984
rect 31852 23792 31904 23798
rect 31850 23760 31852 23769
rect 31904 23760 31906 23769
rect 31850 23695 31906 23704
rect 31956 23186 31984 25978
rect 32048 24721 32076 27338
rect 32140 24970 32168 27338
rect 32220 27328 32272 27334
rect 32220 27270 32272 27276
rect 32232 27130 32260 27270
rect 32220 27124 32272 27130
rect 32220 27066 32272 27072
rect 32404 26852 32456 26858
rect 32404 26794 32456 26800
rect 32312 26240 32364 26246
rect 32312 26182 32364 26188
rect 32324 26042 32352 26182
rect 32312 26036 32364 26042
rect 32312 25978 32364 25984
rect 32416 25906 32444 26794
rect 32508 26042 32536 28086
rect 32600 28014 32628 30670
rect 32784 30138 32812 30670
rect 32876 30666 32904 31282
rect 32864 30660 32916 30666
rect 32864 30602 32916 30608
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 32784 30110 32904 30138
rect 32772 30048 32824 30054
rect 32772 29990 32824 29996
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 32692 27606 32720 29106
rect 32784 28218 32812 29990
rect 32772 28212 32824 28218
rect 32772 28154 32824 28160
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32784 27674 32812 27950
rect 32772 27668 32824 27674
rect 32772 27610 32824 27616
rect 32680 27600 32732 27606
rect 32680 27542 32732 27548
rect 32692 27062 32720 27542
rect 32784 27470 32812 27610
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32680 27056 32732 27062
rect 32680 26998 32732 27004
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 32496 26036 32548 26042
rect 32496 25978 32548 25984
rect 32404 25900 32456 25906
rect 32404 25842 32456 25848
rect 32416 25498 32444 25842
rect 32404 25492 32456 25498
rect 32404 25434 32456 25440
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32404 25288 32456 25294
rect 32404 25230 32456 25236
rect 32140 24942 32260 24970
rect 32324 24954 32352 25230
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32034 24712 32090 24721
rect 32034 24647 32090 24656
rect 32048 23662 32076 24647
rect 32036 23656 32088 23662
rect 32036 23598 32088 23604
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 31956 23050 31984 23122
rect 31944 23044 31996 23050
rect 31944 22986 31996 22992
rect 31668 22976 31720 22982
rect 31668 22918 31720 22924
rect 31576 22432 31628 22438
rect 31576 22374 31628 22380
rect 31588 22166 31616 22374
rect 31576 22160 31628 22166
rect 31576 22102 31628 22108
rect 31588 21706 31616 22102
rect 31680 21894 31708 22918
rect 32036 22160 32088 22166
rect 32034 22128 32036 22137
rect 32088 22128 32090 22137
rect 32034 22063 32090 22072
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31588 21678 31708 21706
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31484 21072 31536 21078
rect 31484 21014 31536 21020
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31208 18964 31260 18970
rect 31208 18906 31260 18912
rect 31024 18692 31076 18698
rect 31024 18634 31076 18640
rect 30932 18080 30984 18086
rect 30932 18022 30984 18028
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 31036 16998 31064 18634
rect 31404 17320 31432 20198
rect 31496 18442 31524 21014
rect 31588 19990 31616 21354
rect 31680 20534 31708 21678
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31668 20528 31720 20534
rect 31668 20470 31720 20476
rect 31576 19984 31628 19990
rect 31576 19926 31628 19932
rect 31680 19700 31708 20470
rect 31772 19854 31800 20878
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31852 19780 31904 19786
rect 31852 19722 31904 19728
rect 31588 19672 31708 19700
rect 31588 19378 31616 19672
rect 31864 19514 31892 19722
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31852 19508 31904 19514
rect 31852 19450 31904 19456
rect 31680 19394 31708 19450
rect 31576 19372 31628 19378
rect 31680 19366 31800 19394
rect 31576 19314 31628 19320
rect 31772 19242 31800 19366
rect 31760 19236 31812 19242
rect 31760 19178 31812 19184
rect 31496 18414 31616 18442
rect 31484 18352 31536 18358
rect 31484 18294 31536 18300
rect 31496 17882 31524 18294
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31404 17292 31524 17320
rect 31392 17196 31444 17202
rect 31128 17156 31392 17184
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30656 16720 30708 16726
rect 30656 16662 30708 16668
rect 30668 16522 30696 16662
rect 30656 16516 30708 16522
rect 30656 16458 30708 16464
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30024 15638 30052 16390
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30116 15706 30144 16050
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 30012 15632 30064 15638
rect 30012 15574 30064 15580
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 29826 14920 29882 14929
rect 29826 14855 29882 14864
rect 29736 14816 29788 14822
rect 29736 14758 29788 14764
rect 29748 14618 29776 14758
rect 29736 14612 29788 14618
rect 29736 14554 29788 14560
rect 29840 14482 29868 14855
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29644 14000 29696 14006
rect 29644 13942 29696 13948
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29564 12850 29592 13670
rect 29656 12986 29684 13942
rect 29748 13394 29776 13942
rect 29736 13388 29788 13394
rect 29736 13330 29788 13336
rect 29932 13190 29960 15506
rect 30288 15496 30340 15502
rect 30340 15456 30420 15484
rect 30288 15438 30340 15444
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30024 14074 30052 14554
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 30300 13938 30328 14758
rect 30392 13938 30420 15456
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30484 14074 30512 14282
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30392 13326 30420 13874
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 30024 12850 30052 13262
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 29460 12368 29512 12374
rect 29460 12310 29512 12316
rect 29472 11898 29500 12310
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 29368 11756 29420 11762
rect 29368 11698 29420 11704
rect 29184 11620 29236 11626
rect 29184 11562 29236 11568
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 27528 11280 27580 11286
rect 27528 11222 27580 11228
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 28368 10810 28396 11018
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 29012 10674 29040 11494
rect 29196 11354 29224 11562
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29840 11150 29868 12718
rect 30484 12306 30512 14010
rect 30576 12782 30604 14418
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30472 12300 30524 12306
rect 30472 12242 30524 12248
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 30024 11694 30052 12038
rect 30576 11694 30604 12378
rect 30668 12238 30696 16458
rect 31128 15502 31156 17156
rect 31392 17138 31444 17144
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 30748 14272 30800 14278
rect 30748 14214 30800 14220
rect 30760 13870 30788 14214
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 30840 13388 30892 13394
rect 30944 13376 30972 14350
rect 30892 13348 30972 13376
rect 30840 13330 30892 13336
rect 30748 13184 30800 13190
rect 30748 13126 30800 13132
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29840 10674 29868 11086
rect 30024 10810 30052 11630
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 30392 10538 30420 11494
rect 30668 11354 30696 12174
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 30576 10266 30604 11018
rect 30564 10260 30616 10266
rect 30564 10202 30616 10208
rect 30760 10062 30788 13126
rect 30944 12832 30972 13348
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 31036 13190 31064 13262
rect 31024 13184 31076 13190
rect 31024 13126 31076 13132
rect 31024 12844 31076 12850
rect 30944 12804 31024 12832
rect 31024 12786 31076 12792
rect 30932 12640 30984 12646
rect 30932 12582 30984 12588
rect 30944 12238 30972 12582
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 30852 11898 30880 12038
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 31036 11694 31064 12786
rect 31128 12442 31156 15438
rect 31312 14550 31340 16458
rect 31496 16454 31524 17292
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31404 15570 31432 15846
rect 31496 15706 31524 16390
rect 31588 15978 31616 18414
rect 31944 18216 31996 18222
rect 31944 18158 31996 18164
rect 31956 17814 31984 18158
rect 31944 17808 31996 17814
rect 31944 17750 31996 17756
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31668 16108 31720 16114
rect 31720 16068 31800 16096
rect 31668 16050 31720 16056
rect 31576 15972 31628 15978
rect 31576 15914 31628 15920
rect 31772 15706 31800 16068
rect 31484 15700 31536 15706
rect 31484 15642 31536 15648
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 31392 15564 31444 15570
rect 31392 15506 31444 15512
rect 31772 15502 31800 15642
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 15162 31800 15438
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 31300 14544 31352 14550
rect 31300 14486 31352 14492
rect 31496 14278 31524 14962
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 31576 14272 31628 14278
rect 31680 14249 31708 14418
rect 31576 14214 31628 14220
rect 31666 14240 31722 14249
rect 31588 14074 31616 14214
rect 31666 14175 31722 14184
rect 31772 14090 31800 14418
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31680 14062 31800 14090
rect 31496 13258 31524 14010
rect 31680 13938 31708 14062
rect 31760 14000 31812 14006
rect 31760 13942 31812 13948
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31668 13388 31720 13394
rect 31668 13330 31720 13336
rect 31484 13252 31536 13258
rect 31484 13194 31536 13200
rect 31680 12986 31708 13330
rect 31772 12986 31800 13942
rect 31864 13530 31892 17274
rect 31944 17060 31996 17066
rect 31944 17002 31996 17008
rect 31956 16522 31984 17002
rect 31944 16516 31996 16522
rect 31944 16458 31996 16464
rect 31956 16046 31984 16458
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 31852 13524 31904 13530
rect 31852 13466 31904 13472
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31864 12986 31892 13262
rect 31668 12980 31720 12986
rect 31668 12922 31720 12928
rect 31760 12980 31812 12986
rect 31760 12922 31812 12928
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31116 12436 31168 12442
rect 31116 12378 31168 12384
rect 31772 12374 31800 12786
rect 31760 12368 31812 12374
rect 31760 12310 31812 12316
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 30932 11688 30984 11694
rect 30932 11630 30984 11636
rect 31024 11688 31076 11694
rect 31024 11630 31076 11636
rect 30944 10674 30972 11630
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30944 10266 30972 10610
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 31036 10130 31064 11290
rect 31772 10810 31800 11698
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31864 10538 31892 12922
rect 32048 12434 32076 21966
rect 32140 20058 32168 24754
rect 32232 22778 32260 24942
rect 32312 24948 32364 24954
rect 32312 24890 32364 24896
rect 32310 24848 32366 24857
rect 32416 24818 32444 25230
rect 32310 24783 32366 24792
rect 32404 24812 32456 24818
rect 32324 23526 32352 24783
rect 32404 24754 32456 24760
rect 32508 24342 32536 25978
rect 32692 25430 32720 26250
rect 32772 25492 32824 25498
rect 32772 25434 32824 25440
rect 32680 25424 32732 25430
rect 32680 25366 32732 25372
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 32692 24750 32720 25230
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 32496 24336 32548 24342
rect 32496 24278 32548 24284
rect 32508 23798 32536 24278
rect 32496 23792 32548 23798
rect 32496 23734 32548 23740
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32416 22681 32444 23462
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32402 22672 32458 22681
rect 32402 22607 32458 22616
rect 32312 22500 32364 22506
rect 32312 22442 32364 22448
rect 32324 22273 32352 22442
rect 32310 22264 32366 22273
rect 32310 22199 32366 22208
rect 32416 21622 32444 22607
rect 32508 22030 32536 22714
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32404 21616 32456 21622
rect 32404 21558 32456 21564
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32232 20602 32260 20878
rect 32220 20596 32272 20602
rect 32220 20538 32272 20544
rect 32600 20466 32628 24618
rect 32784 24206 32812 25434
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32678 23760 32734 23769
rect 32678 23695 32680 23704
rect 32732 23695 32734 23704
rect 32680 23666 32732 23672
rect 32876 23594 32904 30110
rect 32968 28642 32996 30194
rect 33060 29073 33088 34478
rect 33152 33318 33180 35090
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 33244 32434 33272 36858
rect 33324 35624 33376 35630
rect 33324 35566 33376 35572
rect 33336 35086 33364 35566
rect 33428 35290 33456 38286
rect 33600 37868 33652 37874
rect 33600 37810 33652 37816
rect 33508 37664 33560 37670
rect 33508 37606 33560 37612
rect 33520 37126 33548 37606
rect 33612 37262 33640 37810
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33612 37126 33640 37198
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33600 37120 33652 37126
rect 33600 37062 33652 37068
rect 33520 36786 33548 37062
rect 33612 36786 33640 37062
rect 33508 36780 33560 36786
rect 33508 36722 33560 36728
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33600 36644 33652 36650
rect 33600 36586 33652 36592
rect 33612 36242 33640 36586
rect 33704 36582 33732 39335
rect 33796 38758 33824 39986
rect 33876 39296 33928 39302
rect 33876 39238 33928 39244
rect 33784 38752 33836 38758
rect 33784 38694 33836 38700
rect 33796 36922 33824 38694
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 33888 36786 33916 39238
rect 33966 37904 34022 37913
rect 33966 37839 33968 37848
rect 34020 37839 34022 37848
rect 33968 37810 34020 37816
rect 33968 37324 34020 37330
rect 33968 37266 34020 37272
rect 33980 36854 34008 37266
rect 33968 36848 34020 36854
rect 33968 36790 34020 36796
rect 33876 36780 33928 36786
rect 33796 36740 33876 36768
rect 33692 36576 33744 36582
rect 33692 36518 33744 36524
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 33600 36236 33652 36242
rect 33600 36178 33652 36184
rect 33416 35284 33468 35290
rect 33416 35226 33468 35232
rect 33600 35284 33652 35290
rect 33600 35226 33652 35232
rect 33612 35086 33640 35226
rect 33324 35080 33376 35086
rect 33324 35022 33376 35028
rect 33508 35080 33560 35086
rect 33508 35022 33560 35028
rect 33600 35080 33652 35086
rect 33600 35022 33652 35028
rect 33416 35012 33468 35018
rect 33416 34954 33468 34960
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 33140 32224 33192 32230
rect 33140 32166 33192 32172
rect 33152 31890 33180 32166
rect 33230 31920 33286 31929
rect 33140 31884 33192 31890
rect 33230 31855 33232 31864
rect 33140 31826 33192 31832
rect 33284 31855 33286 31864
rect 33232 31826 33284 31832
rect 33046 29064 33102 29073
rect 33046 28999 33102 29008
rect 32968 28614 33088 28642
rect 32956 28552 33008 28558
rect 32956 28494 33008 28500
rect 32968 28218 32996 28494
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 33060 26858 33088 28614
rect 33152 27538 33180 31826
rect 33232 31408 33284 31414
rect 33232 31350 33284 31356
rect 33244 29782 33272 31350
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 33336 30977 33364 31078
rect 33322 30968 33378 30977
rect 33322 30903 33378 30912
rect 33232 29776 33284 29782
rect 33428 29730 33456 34954
rect 33520 34746 33548 35022
rect 33508 34740 33560 34746
rect 33508 34682 33560 34688
rect 33612 34082 33640 35022
rect 33704 34406 33732 36314
rect 33796 35290 33824 36740
rect 33876 36722 33928 36728
rect 33876 36576 33928 36582
rect 33876 36518 33928 36524
rect 33888 36378 33916 36518
rect 33876 36372 33928 36378
rect 33876 36314 33928 36320
rect 33888 35494 33916 36314
rect 33876 35488 33928 35494
rect 33876 35430 33928 35436
rect 33888 35290 33916 35430
rect 33784 35284 33836 35290
rect 33784 35226 33836 35232
rect 33876 35284 33928 35290
rect 33876 35226 33928 35232
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 33692 34400 33744 34406
rect 33692 34342 33744 34348
rect 33612 34054 33732 34082
rect 33598 33960 33654 33969
rect 33598 33895 33600 33904
rect 33652 33895 33654 33904
rect 33600 33866 33652 33872
rect 33508 33856 33560 33862
rect 33508 33798 33560 33804
rect 33520 32502 33548 33798
rect 33704 33658 33732 34054
rect 33796 33658 33824 35022
rect 33888 34728 33916 35226
rect 33968 35216 34020 35222
rect 33968 35158 34020 35164
rect 33980 35086 34008 35158
rect 33968 35080 34020 35086
rect 33968 35022 34020 35028
rect 33968 34740 34020 34746
rect 33888 34700 33968 34728
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 33784 33652 33836 33658
rect 33784 33594 33836 33600
rect 33888 33522 33916 34700
rect 33968 34682 34020 34688
rect 34072 34678 34100 40462
rect 34348 40458 34376 42094
rect 34624 41070 34652 44066
rect 34796 42220 34848 42226
rect 34796 42162 34848 42168
rect 34704 41472 34756 41478
rect 34704 41414 34756 41420
rect 34716 41138 34744 41414
rect 34808 41274 34836 42162
rect 35440 42016 35492 42022
rect 35440 41958 35492 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35452 41614 35480 41958
rect 35440 41608 35492 41614
rect 35440 41550 35492 41556
rect 34796 41268 34848 41274
rect 34796 41210 34848 41216
rect 34704 41132 34756 41138
rect 34704 41074 34756 41080
rect 34428 41064 34480 41070
rect 34428 41006 34480 41012
rect 34612 41064 34664 41070
rect 34612 41006 34664 41012
rect 34440 40730 34468 41006
rect 34428 40724 34480 40730
rect 34428 40666 34480 40672
rect 34336 40452 34388 40458
rect 34336 40394 34388 40400
rect 34152 40180 34204 40186
rect 34152 40122 34204 40128
rect 34164 38418 34192 40122
rect 34612 39840 34664 39846
rect 34612 39782 34664 39788
rect 34520 39432 34572 39438
rect 34520 39374 34572 39380
rect 34244 38956 34296 38962
rect 34244 38898 34296 38904
rect 34428 38956 34480 38962
rect 34428 38898 34480 38904
rect 34256 38758 34284 38898
rect 34244 38752 34296 38758
rect 34244 38694 34296 38700
rect 34152 38412 34204 38418
rect 34204 38372 34376 38400
rect 34152 38354 34204 38360
rect 34152 37868 34204 37874
rect 34152 37810 34204 37816
rect 34164 37398 34192 37810
rect 34152 37392 34204 37398
rect 34152 37334 34204 37340
rect 34152 37256 34204 37262
rect 34152 37198 34204 37204
rect 34242 37224 34298 37233
rect 34164 36786 34192 37198
rect 34242 37159 34298 37168
rect 34256 37126 34284 37159
rect 34244 37120 34296 37126
rect 34244 37062 34296 37068
rect 34348 36854 34376 38372
rect 34440 38350 34468 38898
rect 34428 38344 34480 38350
rect 34428 38286 34480 38292
rect 34532 38282 34560 39374
rect 34520 38276 34572 38282
rect 34520 38218 34572 38224
rect 34428 37868 34480 37874
rect 34428 37810 34480 37816
rect 34440 37482 34468 37810
rect 34532 37670 34560 38218
rect 34520 37664 34572 37670
rect 34520 37606 34572 37612
rect 34440 37454 34560 37482
rect 34532 37262 34560 37454
rect 34520 37256 34572 37262
rect 34624 37233 34652 39782
rect 34716 38894 34744 41074
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 34808 39030 34836 41006
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35716 40520 35768 40526
rect 35716 40462 35768 40468
rect 35440 40044 35492 40050
rect 35440 39986 35492 39992
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35452 39574 35480 39986
rect 35440 39568 35492 39574
rect 35440 39510 35492 39516
rect 35348 39500 35400 39506
rect 35348 39442 35400 39448
rect 34796 39024 34848 39030
rect 34796 38966 34848 38972
rect 34704 38888 34756 38894
rect 34704 38830 34756 38836
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34888 38480 34940 38486
rect 34888 38422 34940 38428
rect 34900 38350 34928 38422
rect 34888 38344 34940 38350
rect 34808 38304 34888 38332
rect 34704 37936 34756 37942
rect 34704 37878 34756 37884
rect 34716 37670 34744 37878
rect 34808 37738 34836 38304
rect 34888 38286 34940 38292
rect 35254 38312 35310 38321
rect 35072 38276 35124 38282
rect 35072 38218 35124 38224
rect 35164 38276 35216 38282
rect 35254 38247 35310 38256
rect 35164 38218 35216 38224
rect 35084 37738 35112 38218
rect 35176 38185 35204 38218
rect 35162 38176 35218 38185
rect 35162 38111 35218 38120
rect 35268 38010 35296 38247
rect 35256 38004 35308 38010
rect 35256 37946 35308 37952
rect 34796 37732 34848 37738
rect 34796 37674 34848 37680
rect 35072 37732 35124 37738
rect 35072 37674 35124 37680
rect 34704 37664 34756 37670
rect 34704 37606 34756 37612
rect 34808 37398 34836 37674
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37392 34848 37398
rect 34796 37334 34848 37340
rect 34796 37256 34848 37262
rect 34520 37198 34572 37204
rect 34610 37224 34666 37233
rect 34428 37188 34480 37194
rect 34666 37182 34744 37210
rect 34796 37198 34848 37204
rect 35072 37256 35124 37262
rect 35072 37198 35124 37204
rect 35164 37256 35216 37262
rect 35216 37216 35296 37244
rect 35164 37198 35216 37204
rect 34610 37159 34666 37168
rect 34428 37130 34480 37136
rect 34336 36848 34388 36854
rect 34336 36790 34388 36796
rect 34152 36780 34204 36786
rect 34152 36722 34204 36728
rect 34152 36644 34204 36650
rect 34152 36586 34204 36592
rect 34164 36258 34192 36586
rect 34440 36378 34468 37130
rect 34612 37120 34664 37126
rect 34612 37062 34664 37068
rect 34428 36372 34480 36378
rect 34428 36314 34480 36320
rect 34624 36258 34652 37062
rect 34164 36230 34652 36258
rect 34244 36168 34296 36174
rect 34244 36110 34296 36116
rect 34152 35692 34204 35698
rect 34152 35634 34204 35640
rect 34060 34672 34112 34678
rect 34060 34614 34112 34620
rect 34164 34377 34192 35634
rect 34256 34542 34284 36110
rect 34624 35494 34652 36230
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 34612 35488 34664 35494
rect 34612 35430 34664 35436
rect 34244 34536 34296 34542
rect 34244 34478 34296 34484
rect 34150 34368 34206 34377
rect 34150 34303 34206 34312
rect 33876 33516 33928 33522
rect 33876 33458 33928 33464
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 33600 33448 33652 33454
rect 33600 33390 33652 33396
rect 33508 32496 33560 32502
rect 33508 32438 33560 32444
rect 33612 32450 33640 33390
rect 33782 32872 33838 32881
rect 33782 32807 33784 32816
rect 33836 32807 33838 32816
rect 33784 32778 33836 32784
rect 33612 32434 33732 32450
rect 33612 32428 33744 32434
rect 33612 32422 33692 32428
rect 33692 32370 33744 32376
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33704 32337 33732 32370
rect 33690 32328 33746 32337
rect 33690 32263 33746 32272
rect 33796 32230 33824 32370
rect 33784 32224 33836 32230
rect 33784 32166 33836 32172
rect 33784 31680 33836 31686
rect 33784 31622 33836 31628
rect 33692 31272 33744 31278
rect 33692 31214 33744 31220
rect 33600 31204 33652 31210
rect 33600 31146 33652 31152
rect 33612 30734 33640 31146
rect 33600 30728 33652 30734
rect 33600 30670 33652 30676
rect 33232 29718 33284 29724
rect 33244 29646 33272 29718
rect 33336 29702 33456 29730
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33230 28248 33286 28257
rect 33230 28183 33232 28192
rect 33284 28183 33286 28192
rect 33232 28154 33284 28160
rect 33140 27532 33192 27538
rect 33140 27474 33192 27480
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 33140 26784 33192 26790
rect 33140 26726 33192 26732
rect 33152 26450 33180 26726
rect 33336 26466 33364 29702
rect 33416 29640 33468 29646
rect 33468 29600 33548 29628
rect 33416 29582 33468 29588
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33428 27470 33456 29106
rect 33520 29034 33548 29600
rect 33612 29170 33640 30670
rect 33704 30190 33732 31214
rect 33796 30938 33824 31622
rect 33784 30932 33836 30938
rect 33784 30874 33836 30880
rect 33888 30818 33916 33458
rect 33968 33312 34020 33318
rect 33968 33254 34020 33260
rect 33980 32910 34008 33254
rect 33968 32904 34020 32910
rect 33968 32846 34020 32852
rect 34072 32774 34100 33458
rect 33968 32768 34020 32774
rect 33968 32710 34020 32716
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 33980 32570 34008 32710
rect 33968 32564 34020 32570
rect 33968 32506 34020 32512
rect 33966 32056 34022 32065
rect 33966 31991 34022 32000
rect 33980 31414 34008 31991
rect 34072 31657 34100 32710
rect 34256 32230 34284 34478
rect 34440 33998 34468 35430
rect 34624 35136 34652 35430
rect 34532 35108 34652 35136
rect 34532 35018 34560 35108
rect 34520 35012 34572 35018
rect 34520 34954 34572 34960
rect 34612 35012 34664 35018
rect 34612 34954 34664 34960
rect 34428 33992 34480 33998
rect 34428 33934 34480 33940
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34336 33108 34388 33114
rect 34336 33050 34388 33056
rect 34348 32570 34376 33050
rect 34336 32564 34388 32570
rect 34336 32506 34388 32512
rect 34428 32292 34480 32298
rect 34428 32234 34480 32240
rect 34244 32224 34296 32230
rect 34244 32166 34296 32172
rect 34256 32026 34284 32166
rect 34244 32020 34296 32026
rect 34244 31962 34296 31968
rect 34256 31890 34284 31962
rect 34244 31884 34296 31890
rect 34244 31826 34296 31832
rect 34440 31822 34468 32234
rect 34428 31816 34480 31822
rect 34428 31758 34480 31764
rect 34058 31648 34114 31657
rect 34058 31583 34114 31592
rect 33968 31408 34020 31414
rect 33968 31350 34020 31356
rect 33796 30790 33916 30818
rect 34152 30796 34204 30802
rect 33692 30184 33744 30190
rect 33692 30126 33744 30132
rect 33600 29164 33652 29170
rect 33600 29106 33652 29112
rect 33508 29028 33560 29034
rect 33796 28994 33824 30790
rect 34152 30738 34204 30744
rect 34164 30258 34192 30738
rect 34440 30734 34468 31758
rect 34428 30728 34480 30734
rect 34428 30670 34480 30676
rect 34440 30546 34468 30670
rect 34348 30518 34468 30546
rect 33968 30252 34020 30258
rect 33888 30212 33968 30240
rect 33888 29646 33916 30212
rect 33968 30194 34020 30200
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 33968 30116 34020 30122
rect 33968 30058 34020 30064
rect 33876 29640 33928 29646
rect 33876 29582 33928 29588
rect 33508 28970 33560 28976
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33140 26444 33192 26450
rect 33140 26386 33192 26392
rect 33244 26438 33364 26466
rect 33046 26072 33102 26081
rect 33046 26007 33102 26016
rect 33060 25974 33088 26007
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 33060 24410 33088 25910
rect 33152 25906 33180 26386
rect 33244 26314 33272 26438
rect 33322 26344 33378 26353
rect 33232 26308 33284 26314
rect 33322 26279 33378 26288
rect 33232 26250 33284 26256
rect 33232 26036 33284 26042
rect 33232 25978 33284 25984
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 33244 24274 33272 25978
rect 33232 24268 33284 24274
rect 33232 24210 33284 24216
rect 32864 23588 32916 23594
rect 32864 23530 32916 23536
rect 33244 23322 33272 24210
rect 33232 23316 33284 23322
rect 33232 23258 33284 23264
rect 33138 23216 33194 23225
rect 33138 23151 33194 23160
rect 33152 23118 33180 23151
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 32956 22704 33008 22710
rect 32956 22646 33008 22652
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32876 21554 32904 22374
rect 32968 22030 32996 22646
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 32864 21548 32916 21554
rect 32864 21490 32916 21496
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32140 19378 32168 19994
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32324 19242 32352 20402
rect 32416 20330 32444 20402
rect 32404 20324 32456 20330
rect 32404 20266 32456 20272
rect 32312 19236 32364 19242
rect 32312 19178 32364 19184
rect 32324 18426 32352 19178
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 32140 17202 32168 17478
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32416 16794 32444 20266
rect 32600 18630 32628 20402
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32404 16788 32456 16794
rect 32404 16730 32456 16736
rect 32508 16658 32536 18090
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32312 16584 32364 16590
rect 32312 16526 32364 16532
rect 32324 16425 32352 16526
rect 32310 16416 32366 16425
rect 32310 16351 32366 16360
rect 32324 16114 32352 16351
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32404 15360 32456 15366
rect 32508 15337 32536 16594
rect 32600 16153 32628 18226
rect 32586 16144 32642 16153
rect 32586 16079 32642 16088
rect 32404 15302 32456 15308
rect 32494 15328 32550 15337
rect 32220 13728 32272 13734
rect 32220 13670 32272 13676
rect 32232 13410 32260 13670
rect 32232 13382 32352 13410
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 32232 12832 32260 13262
rect 32140 12804 32260 12832
rect 32140 12646 32168 12804
rect 32324 12730 32352 13382
rect 32416 12986 32444 15302
rect 32494 15263 32550 15272
rect 32508 14414 32536 15263
rect 32600 14482 32628 16079
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32496 13728 32548 13734
rect 32496 13670 32548 13676
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32508 12850 32536 13670
rect 32496 12844 32548 12850
rect 32232 12702 32352 12730
rect 32416 12804 32496 12832
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 31956 12406 32076 12434
rect 31956 11354 31984 12406
rect 32140 12306 32168 12582
rect 32232 12442 32260 12702
rect 32416 12594 32444 12804
rect 32496 12786 32548 12792
rect 32324 12566 32444 12594
rect 32220 12436 32272 12442
rect 32220 12378 32272 12384
rect 32324 12306 32352 12566
rect 32128 12300 32180 12306
rect 32128 12242 32180 12248
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 32048 11830 32076 12038
rect 32232 11898 32260 12174
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 32588 11892 32640 11898
rect 32588 11834 32640 11840
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 32218 11384 32274 11393
rect 31944 11348 31996 11354
rect 32218 11319 32220 11328
rect 31944 11290 31996 11296
rect 32272 11319 32274 11328
rect 32220 11290 32272 11296
rect 32600 10674 32628 11834
rect 32692 11762 32720 21354
rect 32968 20942 32996 21966
rect 33152 21486 33180 22578
rect 33140 21480 33192 21486
rect 33140 21422 33192 21428
rect 33048 21344 33100 21350
rect 33048 21286 33100 21292
rect 33060 20942 33088 21286
rect 33152 21146 33180 21422
rect 33140 21140 33192 21146
rect 33140 21082 33192 21088
rect 33152 21010 33180 21082
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32784 20466 32812 20742
rect 32772 20460 32824 20466
rect 32772 20402 32824 20408
rect 32772 20256 32824 20262
rect 32772 20198 32824 20204
rect 32784 18766 32812 20198
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32876 17678 32904 20878
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 33060 19854 33088 20402
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33060 19378 33088 19790
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 33336 18850 33364 26279
rect 33428 25786 33456 27406
rect 33520 26994 33548 28970
rect 33704 28966 33824 28994
rect 33876 29028 33928 29034
rect 33876 28970 33928 28976
rect 33600 27396 33652 27402
rect 33600 27338 33652 27344
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33520 26314 33548 26930
rect 33508 26308 33560 26314
rect 33508 26250 33560 26256
rect 33612 25922 33640 27338
rect 33704 26042 33732 28966
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 33796 27878 33824 28698
rect 33888 28558 33916 28970
rect 33980 28558 34008 30058
rect 34060 29776 34112 29782
rect 34060 29718 34112 29724
rect 34072 29646 34100 29718
rect 34060 29640 34112 29646
rect 34060 29582 34112 29588
rect 34060 29504 34112 29510
rect 34060 29446 34112 29452
rect 34072 28762 34100 29446
rect 34164 28966 34192 30194
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 34152 28960 34204 28966
rect 34152 28902 34204 28908
rect 34060 28756 34112 28762
rect 34060 28698 34112 28704
rect 34072 28558 34100 28698
rect 33876 28552 33928 28558
rect 33876 28494 33928 28500
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 34060 28552 34112 28558
rect 34060 28494 34112 28500
rect 34256 28200 34284 29582
rect 34072 28172 34284 28200
rect 33784 27872 33836 27878
rect 33784 27814 33836 27820
rect 34072 27470 34100 28172
rect 34348 28098 34376 30518
rect 34426 30424 34482 30433
rect 34532 30410 34560 33934
rect 34624 33046 34652 34954
rect 34716 34950 34744 37182
rect 34808 36292 34836 37198
rect 35084 37126 35112 37198
rect 35072 37120 35124 37126
rect 35072 37062 35124 37068
rect 35162 36952 35218 36961
rect 35162 36887 35218 36896
rect 35176 36786 35204 36887
rect 35164 36780 35216 36786
rect 35164 36722 35216 36728
rect 35268 36530 35296 37216
rect 35360 36922 35388 39442
rect 35530 38992 35586 39001
rect 35530 38927 35532 38936
rect 35584 38927 35586 38936
rect 35624 38956 35676 38962
rect 35532 38898 35584 38904
rect 35624 38898 35676 38904
rect 35440 38888 35492 38894
rect 35440 38830 35492 38836
rect 35452 37126 35480 38830
rect 35636 38554 35664 38898
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 35530 37904 35586 37913
rect 35530 37839 35532 37848
rect 35584 37839 35586 37848
rect 35532 37810 35584 37816
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 35348 36916 35400 36922
rect 35348 36858 35400 36864
rect 35268 36502 35388 36530
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34888 36304 34940 36310
rect 34808 36264 34888 36292
rect 34888 36246 34940 36252
rect 34900 35698 34928 36246
rect 34992 36230 35296 36258
rect 35360 36242 35388 36502
rect 34992 36106 35020 36230
rect 34980 36100 35032 36106
rect 34980 36042 35032 36048
rect 35164 36100 35216 36106
rect 35164 36042 35216 36048
rect 34888 35692 34940 35698
rect 34888 35634 34940 35640
rect 34992 35630 35020 36042
rect 35072 35760 35124 35766
rect 35072 35702 35124 35708
rect 34980 35624 35032 35630
rect 34980 35566 35032 35572
rect 35084 35494 35112 35702
rect 35176 35698 35204 36042
rect 35268 36038 35296 36230
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 35256 36032 35308 36038
rect 35256 35974 35308 35980
rect 35346 35864 35402 35873
rect 35346 35799 35402 35808
rect 35256 35760 35308 35766
rect 35256 35702 35308 35708
rect 35164 35692 35216 35698
rect 35164 35634 35216 35640
rect 35268 35562 35296 35702
rect 35256 35556 35308 35562
rect 35256 35498 35308 35504
rect 35072 35488 35124 35494
rect 35072 35430 35124 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34888 35216 34940 35222
rect 34886 35184 34888 35193
rect 34940 35184 34942 35193
rect 34886 35119 34942 35128
rect 35360 35086 35388 35799
rect 35348 35080 35400 35086
rect 35348 35022 35400 35028
rect 34704 34944 34756 34950
rect 34704 34886 34756 34892
rect 34716 33522 34744 34886
rect 35348 34740 35400 34746
rect 35348 34682 35400 34688
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 33930 35388 34682
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 34704 33516 34756 33522
rect 34704 33458 34756 33464
rect 35256 33448 35308 33454
rect 35256 33390 35308 33396
rect 35268 33266 35296 33390
rect 35268 33238 35388 33266
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34612 33040 34664 33046
rect 34612 32982 34664 32988
rect 34624 32026 34652 32982
rect 35360 32978 35388 33238
rect 35348 32972 35400 32978
rect 35348 32914 35400 32920
rect 35162 32464 35218 32473
rect 35162 32399 35164 32408
rect 35216 32399 35218 32408
rect 35164 32370 35216 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34612 32020 34664 32026
rect 34612 31962 34664 31968
rect 34704 31952 34756 31958
rect 34610 31920 34666 31929
rect 34704 31894 34756 31900
rect 34610 31855 34666 31864
rect 34624 31754 34652 31855
rect 34716 31754 34744 31894
rect 34612 31748 34664 31754
rect 34716 31726 34836 31754
rect 35072 31748 35124 31754
rect 34612 31690 34664 31696
rect 34482 30382 34560 30410
rect 34426 30359 34482 30368
rect 34518 30288 34574 30297
rect 34518 30223 34520 30232
rect 34572 30223 34574 30232
rect 34520 30194 34572 30200
rect 34532 29646 34560 30194
rect 34520 29640 34572 29646
rect 34518 29608 34520 29617
rect 34572 29608 34574 29617
rect 34428 29572 34480 29578
rect 34518 29543 34574 29552
rect 34428 29514 34480 29520
rect 34440 29170 34468 29514
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34532 29238 34560 29446
rect 34520 29232 34572 29238
rect 34520 29174 34572 29180
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34440 28218 34468 28426
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34164 28070 34376 28098
rect 34532 28082 34560 29174
rect 34624 29152 34652 31690
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34716 30734 34744 31282
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 34716 29306 34744 30670
rect 34704 29300 34756 29306
rect 34704 29242 34756 29248
rect 34704 29164 34756 29170
rect 34624 29124 34704 29152
rect 34704 29106 34756 29112
rect 34704 28620 34756 28626
rect 34704 28562 34756 28568
rect 34612 28552 34664 28558
rect 34612 28494 34664 28500
rect 34520 28076 34572 28082
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 33968 27056 34020 27062
rect 33968 26998 34020 27004
rect 33876 26852 33928 26858
rect 33876 26794 33928 26800
rect 33888 26518 33916 26794
rect 33876 26512 33928 26518
rect 33876 26454 33928 26460
rect 33784 26376 33836 26382
rect 33782 26344 33784 26353
rect 33836 26344 33838 26353
rect 33782 26279 33838 26288
rect 33692 26036 33744 26042
rect 33692 25978 33744 25984
rect 33612 25894 33732 25922
rect 33428 25758 33548 25786
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 33428 22778 33456 25638
rect 33520 25294 33548 25758
rect 33508 25288 33560 25294
rect 33508 25230 33560 25236
rect 33704 25226 33732 25894
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33692 25220 33744 25226
rect 33692 25162 33744 25168
rect 33600 24744 33652 24750
rect 33600 24686 33652 24692
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33520 23730 33548 24278
rect 33612 24206 33640 24686
rect 33600 24200 33652 24206
rect 33600 24142 33652 24148
rect 33704 23798 33732 25162
rect 33796 24818 33824 25230
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33876 24268 33928 24274
rect 33796 24228 33876 24256
rect 33692 23792 33744 23798
rect 33692 23734 33744 23740
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33428 22030 33456 22714
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33520 21418 33548 23258
rect 33796 23050 33824 24228
rect 33876 24210 33928 24216
rect 33980 23322 34008 26998
rect 34060 26784 34112 26790
rect 34060 26726 34112 26732
rect 34072 26382 34100 26726
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 34058 26208 34114 26217
rect 34058 26143 34114 26152
rect 34072 26042 34100 26143
rect 34060 26036 34112 26042
rect 34060 25978 34112 25984
rect 34072 25498 34100 25978
rect 34164 25770 34192 28070
rect 34520 28018 34572 28024
rect 34244 28008 34296 28014
rect 34244 27950 34296 27956
rect 34336 28008 34388 28014
rect 34336 27950 34388 27956
rect 34428 28008 34480 28014
rect 34518 27976 34574 27985
rect 34480 27956 34518 27962
rect 34428 27950 34518 27956
rect 34256 27538 34284 27950
rect 34348 27656 34376 27950
rect 34440 27934 34518 27950
rect 34518 27911 34574 27920
rect 34428 27668 34480 27674
rect 34348 27628 34428 27656
rect 34428 27610 34480 27616
rect 34532 27577 34560 27911
rect 34624 27606 34652 28494
rect 34612 27600 34664 27606
rect 34518 27568 34574 27577
rect 34244 27532 34296 27538
rect 34612 27542 34664 27548
rect 34518 27503 34574 27512
rect 34244 27474 34296 27480
rect 34256 26994 34284 27474
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34348 26926 34376 27406
rect 34336 26920 34388 26926
rect 34334 26888 34336 26897
rect 34388 26888 34390 26897
rect 34334 26823 34390 26832
rect 34428 26852 34480 26858
rect 34428 26794 34480 26800
rect 34440 26217 34468 26794
rect 34532 26586 34560 27503
rect 34716 27062 34744 28562
rect 34704 27056 34756 27062
rect 34704 26998 34756 27004
rect 34808 26994 34836 31726
rect 34992 31708 35072 31736
rect 34992 31346 35020 31708
rect 35072 31690 35124 31696
rect 34980 31340 35032 31346
rect 34980 31282 35032 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30841 35388 32914
rect 35452 32434 35480 37062
rect 35544 36825 35572 37810
rect 35624 37256 35676 37262
rect 35624 37198 35676 37204
rect 35530 36816 35586 36825
rect 35530 36751 35586 36760
rect 35636 36310 35664 37198
rect 35624 36304 35676 36310
rect 35624 36246 35676 36252
rect 35532 36032 35584 36038
rect 35532 35974 35584 35980
rect 35544 35086 35572 35974
rect 35624 35828 35676 35834
rect 35624 35770 35676 35776
rect 35532 35080 35584 35086
rect 35532 35022 35584 35028
rect 35636 35018 35664 35770
rect 35624 35012 35676 35018
rect 35624 34954 35676 34960
rect 35636 32978 35664 34954
rect 35728 33114 35756 40462
rect 35912 40390 35940 44118
rect 36084 42016 36136 42022
rect 36084 41958 36136 41964
rect 36176 42016 36228 42022
rect 36176 41958 36228 41964
rect 35900 40384 35952 40390
rect 35900 40326 35952 40332
rect 36096 39953 36124 41958
rect 36082 39944 36138 39953
rect 36082 39879 36138 39888
rect 36084 39636 36136 39642
rect 36084 39578 36136 39584
rect 36096 39506 36124 39578
rect 36084 39500 36136 39506
rect 36084 39442 36136 39448
rect 35992 39296 36044 39302
rect 35992 39238 36044 39244
rect 36084 39296 36136 39302
rect 36084 39238 36136 39244
rect 36004 39030 36032 39238
rect 35992 39024 36044 39030
rect 35992 38966 36044 38972
rect 35992 38208 36044 38214
rect 35992 38150 36044 38156
rect 35900 37868 35952 37874
rect 35900 37810 35952 37816
rect 35808 37800 35860 37806
rect 35808 37742 35860 37748
rect 35820 36854 35848 37742
rect 35808 36848 35860 36854
rect 35808 36790 35860 36796
rect 35820 35834 35848 36790
rect 35912 36786 35940 37810
rect 35900 36780 35952 36786
rect 35900 36722 35952 36728
rect 35912 36650 35940 36722
rect 35900 36644 35952 36650
rect 35900 36586 35952 36592
rect 35900 36168 35952 36174
rect 35898 36136 35900 36145
rect 35952 36136 35954 36145
rect 35898 36071 35954 36080
rect 36004 36088 36032 38150
rect 36096 38010 36124 39238
rect 36084 38004 36136 38010
rect 36084 37946 36136 37952
rect 36188 37913 36216 41958
rect 36728 41608 36780 41614
rect 36728 41550 36780 41556
rect 36912 41608 36964 41614
rect 36912 41550 36964 41556
rect 36268 41472 36320 41478
rect 36268 41414 36320 41420
rect 36280 41138 36308 41414
rect 36268 41132 36320 41138
rect 36268 41074 36320 41080
rect 36452 40384 36504 40390
rect 36452 40326 36504 40332
rect 36268 39296 36320 39302
rect 36268 39238 36320 39244
rect 36280 38962 36308 39238
rect 36268 38956 36320 38962
rect 36268 38898 36320 38904
rect 36464 38554 36492 40326
rect 36636 40044 36688 40050
rect 36636 39986 36688 39992
rect 36452 38548 36504 38554
rect 36452 38490 36504 38496
rect 36648 38214 36676 39986
rect 36740 39982 36768 41550
rect 36924 40730 36952 41550
rect 37004 40928 37056 40934
rect 37004 40870 37056 40876
rect 36912 40724 36964 40730
rect 36912 40666 36964 40672
rect 37016 40526 37044 40870
rect 37004 40520 37056 40526
rect 37004 40462 37056 40468
rect 37188 40452 37240 40458
rect 37292 40440 37320 44200
rect 37924 42356 37976 42362
rect 37924 42298 37976 42304
rect 37556 42288 37608 42294
rect 37556 42230 37608 42236
rect 37568 41818 37596 42230
rect 37556 41812 37608 41818
rect 37556 41754 37608 41760
rect 37464 41608 37516 41614
rect 37464 41550 37516 41556
rect 37476 40730 37504 41550
rect 37568 41414 37596 41754
rect 37740 41472 37792 41478
rect 37740 41414 37792 41420
rect 37568 41386 37688 41414
rect 37464 40724 37516 40730
rect 37464 40666 37516 40672
rect 37464 40452 37516 40458
rect 37292 40412 37464 40440
rect 37188 40394 37240 40400
rect 37464 40394 37516 40400
rect 37096 40180 37148 40186
rect 37096 40122 37148 40128
rect 36728 39976 36780 39982
rect 36728 39918 36780 39924
rect 36912 39568 36964 39574
rect 36912 39510 36964 39516
rect 36924 38962 36952 39510
rect 36912 38956 36964 38962
rect 36912 38898 36964 38904
rect 37108 38654 37136 40122
rect 37200 39574 37228 40394
rect 37188 39568 37240 39574
rect 37188 39510 37240 39516
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 36740 38626 37136 38654
rect 36636 38208 36688 38214
rect 36636 38150 36688 38156
rect 36174 37904 36230 37913
rect 36174 37839 36230 37848
rect 36452 37868 36504 37874
rect 36452 37810 36504 37816
rect 36544 37868 36596 37874
rect 36544 37810 36596 37816
rect 36464 37738 36492 37810
rect 36452 37732 36504 37738
rect 36452 37674 36504 37680
rect 36360 37460 36412 37466
rect 36360 37402 36412 37408
rect 36176 37188 36228 37194
rect 36176 37130 36228 37136
rect 36188 36854 36216 37130
rect 36176 36848 36228 36854
rect 36176 36790 36228 36796
rect 36084 36100 36136 36106
rect 35808 35828 35860 35834
rect 35808 35770 35860 35776
rect 35820 35562 35848 35770
rect 35808 35556 35860 35562
rect 35808 35498 35860 35504
rect 35808 35284 35860 35290
rect 35808 35226 35860 35232
rect 35820 34950 35848 35226
rect 35808 34944 35860 34950
rect 35808 34886 35860 34892
rect 35808 33992 35860 33998
rect 35806 33960 35808 33969
rect 35860 33960 35862 33969
rect 35806 33895 35862 33904
rect 35912 33454 35940 36071
rect 36004 36060 36084 36088
rect 36084 36042 36136 36048
rect 35992 35692 36044 35698
rect 35992 35634 36044 35640
rect 36004 34388 36032 35634
rect 36096 34542 36124 36042
rect 36188 35562 36216 36790
rect 36372 36786 36400 37402
rect 36464 37380 36492 37674
rect 36556 37505 36584 37810
rect 36740 37806 36768 38626
rect 36820 38344 36872 38350
rect 36820 38286 36872 38292
rect 37096 38344 37148 38350
rect 37292 38321 37320 38694
rect 37372 38344 37424 38350
rect 37096 38286 37148 38292
rect 37278 38312 37334 38321
rect 36832 37874 36860 38286
rect 37004 38208 37056 38214
rect 37004 38150 37056 38156
rect 37016 37874 37044 38150
rect 36820 37868 36872 37874
rect 36820 37810 36872 37816
rect 37004 37868 37056 37874
rect 37004 37810 37056 37816
rect 36728 37800 36780 37806
rect 36728 37742 36780 37748
rect 36636 37664 36688 37670
rect 36636 37606 36688 37612
rect 36542 37496 36598 37505
rect 36542 37431 36598 37440
rect 36464 37352 36584 37380
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 36360 36780 36412 36786
rect 36360 36722 36412 36728
rect 36372 36582 36400 36722
rect 36360 36576 36412 36582
rect 36360 36518 36412 36524
rect 36268 36236 36320 36242
rect 36268 36178 36320 36184
rect 36176 35556 36228 35562
rect 36176 35498 36228 35504
rect 36188 35222 36216 35498
rect 36280 35290 36308 36178
rect 36268 35284 36320 35290
rect 36268 35226 36320 35232
rect 36176 35216 36228 35222
rect 36176 35158 36228 35164
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 36360 35012 36412 35018
rect 36464 35000 36492 37198
rect 36556 37194 36584 37352
rect 36648 37330 36676 37606
rect 36636 37324 36688 37330
rect 36636 37266 36688 37272
rect 36544 37188 36596 37194
rect 36544 37130 36596 37136
rect 36636 36780 36688 36786
rect 36412 34972 36492 35000
rect 36556 36740 36636 36768
rect 36360 34954 36412 34960
rect 36188 34610 36216 34954
rect 36176 34604 36228 34610
rect 36176 34546 36228 34552
rect 36084 34536 36136 34542
rect 36084 34478 36136 34484
rect 36004 34360 36216 34388
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 35716 33108 35768 33114
rect 35716 33050 35768 33056
rect 35900 33040 35952 33046
rect 35900 32982 35952 32988
rect 35624 32972 35676 32978
rect 35624 32914 35676 32920
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35714 32600 35770 32609
rect 35714 32535 35770 32544
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 35452 31958 35480 32166
rect 35440 31952 35492 31958
rect 35440 31894 35492 31900
rect 35728 31754 35756 32535
rect 35820 32298 35848 32846
rect 35808 32292 35860 32298
rect 35808 32234 35860 32240
rect 35440 31748 35492 31754
rect 35440 31690 35492 31696
rect 35716 31748 35768 31754
rect 35716 31690 35768 31696
rect 35452 31634 35480 31690
rect 35452 31606 35572 31634
rect 35544 31414 35572 31606
rect 35532 31408 35584 31414
rect 35532 31350 35584 31356
rect 35714 31376 35770 31385
rect 35438 31104 35494 31113
rect 35438 31039 35494 31048
rect 35346 30832 35402 30841
rect 35346 30767 35402 30776
rect 35452 30734 35480 31039
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29782 35388 30194
rect 35348 29776 35400 29782
rect 35348 29718 35400 29724
rect 35164 29504 35216 29510
rect 35164 29446 35216 29452
rect 35176 29306 35204 29446
rect 35164 29300 35216 29306
rect 35164 29242 35216 29248
rect 34888 29232 34940 29238
rect 34888 29174 34940 29180
rect 35348 29232 35400 29238
rect 35348 29174 35400 29180
rect 34900 29034 34928 29174
rect 34888 29028 34940 29034
rect 34888 28970 34940 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28762 35388 29174
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35452 28529 35480 30670
rect 35544 30274 35572 31350
rect 35714 31311 35770 31320
rect 35728 31278 35756 31311
rect 35716 31272 35768 31278
rect 35716 31214 35768 31220
rect 35716 31136 35768 31142
rect 35716 31078 35768 31084
rect 35624 30728 35676 30734
rect 35624 30670 35676 30676
rect 35636 30394 35664 30670
rect 35624 30388 35676 30394
rect 35624 30330 35676 30336
rect 35544 30246 35664 30274
rect 35728 30258 35756 31078
rect 35808 30932 35860 30938
rect 35808 30874 35860 30880
rect 35820 30258 35848 30874
rect 35636 29209 35664 30246
rect 35716 30252 35768 30258
rect 35716 30194 35768 30200
rect 35808 30252 35860 30258
rect 35808 30194 35860 30200
rect 35622 29200 35678 29209
rect 35622 29135 35678 29144
rect 35624 29028 35676 29034
rect 35624 28970 35676 28976
rect 35532 28960 35584 28966
rect 35532 28902 35584 28908
rect 35438 28520 35494 28529
rect 35348 28484 35400 28490
rect 35438 28455 35494 28464
rect 35348 28426 35400 28432
rect 35162 28112 35218 28121
rect 35162 28047 35164 28056
rect 35216 28047 35218 28056
rect 35164 28018 35216 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27674 35388 28426
rect 35440 28212 35492 28218
rect 35440 28154 35492 28160
rect 34980 27668 35032 27674
rect 34980 27610 35032 27616
rect 35348 27668 35400 27674
rect 35348 27610 35400 27616
rect 34992 27452 35020 27610
rect 35072 27464 35124 27470
rect 34992 27424 35072 27452
rect 34992 27334 35020 27424
rect 35072 27406 35124 27412
rect 34980 27328 35032 27334
rect 34980 27270 35032 27276
rect 35164 27328 35216 27334
rect 35164 27270 35216 27276
rect 35176 26994 35204 27270
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 35164 26988 35216 26994
rect 35164 26930 35216 26936
rect 34704 26784 34756 26790
rect 34704 26726 34756 26732
rect 34520 26580 34572 26586
rect 34520 26522 34572 26528
rect 34612 26376 34664 26382
rect 34612 26318 34664 26324
rect 34520 26240 34572 26246
rect 34426 26208 34482 26217
rect 34520 26182 34572 26188
rect 34426 26143 34482 26152
rect 34152 25764 34204 25770
rect 34152 25706 34204 25712
rect 34060 25492 34112 25498
rect 34060 25434 34112 25440
rect 34440 24800 34468 26143
rect 34532 25362 34560 26182
rect 34624 25770 34652 26318
rect 34716 25974 34744 26726
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 34612 25764 34664 25770
rect 34612 25706 34664 25712
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 34612 25220 34664 25226
rect 34612 25162 34664 25168
rect 34520 24812 34572 24818
rect 34440 24772 34520 24800
rect 34520 24754 34572 24760
rect 34428 24676 34480 24682
rect 34428 24618 34480 24624
rect 34242 24304 34298 24313
rect 34242 24239 34298 24248
rect 34336 24268 34388 24274
rect 34256 24206 34284 24239
rect 34336 24210 34388 24216
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 34152 24064 34204 24070
rect 34152 24006 34204 24012
rect 34164 23905 34192 24006
rect 34150 23896 34206 23905
rect 34150 23831 34206 23840
rect 34164 23730 34192 23831
rect 34256 23730 34284 24142
rect 34348 23866 34376 24210
rect 34440 24206 34468 24618
rect 34520 24608 34572 24614
rect 34520 24550 34572 24556
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34336 23860 34388 23866
rect 34336 23802 34388 23808
rect 34152 23724 34204 23730
rect 34152 23666 34204 23672
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33600 23044 33652 23050
rect 33600 22986 33652 22992
rect 33784 23044 33836 23050
rect 33784 22986 33836 22992
rect 33612 22506 33640 22986
rect 33796 22710 33824 22986
rect 33784 22704 33836 22710
rect 33784 22646 33836 22652
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33612 21554 33640 22442
rect 33888 22098 33916 23054
rect 34348 22778 34376 23802
rect 34060 22772 34112 22778
rect 34060 22714 34112 22720
rect 34336 22772 34388 22778
rect 34336 22714 34388 22720
rect 33968 22704 34020 22710
rect 33968 22646 34020 22652
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33980 21554 34008 22646
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33968 21548 34020 21554
rect 33968 21490 34020 21496
rect 34072 21418 34100 22714
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 33508 21412 33560 21418
rect 33508 21354 33560 21360
rect 34060 21412 34112 21418
rect 34060 21354 34112 21360
rect 34348 21146 34376 21830
rect 34532 21570 34560 24550
rect 34624 21690 34652 25162
rect 34716 24954 34744 25910
rect 34704 24948 34756 24954
rect 34704 24890 34756 24896
rect 34704 24608 34756 24614
rect 34704 24550 34756 24556
rect 34716 23798 34744 24550
rect 34808 23866 34836 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35254 26344 35310 26353
rect 35254 26279 35256 26288
rect 35308 26279 35310 26288
rect 35256 26250 35308 26256
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35072 25356 35124 25362
rect 35072 25298 35124 25304
rect 34980 25288 35032 25294
rect 34980 25230 35032 25236
rect 34992 24818 35020 25230
rect 34980 24812 35032 24818
rect 34980 24754 35032 24760
rect 35084 24682 35112 25298
rect 35256 25288 35308 25294
rect 35256 25230 35308 25236
rect 35268 24682 35296 25230
rect 35360 25226 35388 25638
rect 35452 25242 35480 28154
rect 35544 27674 35572 28902
rect 35532 27668 35584 27674
rect 35532 27610 35584 27616
rect 35636 27470 35664 28970
rect 35728 27538 35756 30194
rect 35912 29730 35940 32982
rect 36004 32978 36032 34138
rect 36084 33380 36136 33386
rect 36084 33322 36136 33328
rect 35992 32972 36044 32978
rect 35992 32914 36044 32920
rect 36096 32910 36124 33322
rect 36084 32904 36136 32910
rect 36084 32846 36136 32852
rect 36096 32434 36124 32846
rect 36188 32434 36216 34360
rect 36372 33844 36400 34954
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 36464 34513 36492 34546
rect 36450 34504 36506 34513
rect 36450 34439 36506 34448
rect 36452 33856 36504 33862
rect 36372 33816 36452 33844
rect 36452 33798 36504 33804
rect 36266 33144 36322 33153
rect 36266 33079 36322 33088
rect 36084 32428 36136 32434
rect 36084 32370 36136 32376
rect 36176 32428 36228 32434
rect 36176 32370 36228 32376
rect 36096 32337 36124 32370
rect 36082 32328 36138 32337
rect 36082 32263 36138 32272
rect 36188 31906 36216 32370
rect 36004 31878 36216 31906
rect 36004 31822 36032 31878
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 36084 31816 36136 31822
rect 36084 31758 36136 31764
rect 35992 31408 36044 31414
rect 35992 31350 36044 31356
rect 36004 29850 36032 31350
rect 36096 31210 36124 31758
rect 36280 31754 36308 33079
rect 36464 32366 36492 33798
rect 36556 33561 36584 36740
rect 36636 36722 36688 36728
rect 36740 36564 36768 37742
rect 36832 37262 36860 37810
rect 36912 37800 36964 37806
rect 36912 37742 36964 37748
rect 36924 37466 36952 37742
rect 36912 37460 36964 37466
rect 36912 37402 36964 37408
rect 36820 37256 36872 37262
rect 36820 37198 36872 37204
rect 36832 36786 36860 37198
rect 36820 36780 36872 36786
rect 37016 36768 37044 37810
rect 37108 37398 37136 38286
rect 37372 38286 37424 38292
rect 37278 38247 37334 38256
rect 37384 38010 37412 38286
rect 37372 38004 37424 38010
rect 37372 37946 37424 37952
rect 37476 37466 37504 40394
rect 37556 39840 37608 39846
rect 37556 39782 37608 39788
rect 37464 37460 37516 37466
rect 37464 37402 37516 37408
rect 37096 37392 37148 37398
rect 37096 37334 37148 37340
rect 36820 36722 36872 36728
rect 36924 36740 37044 36768
rect 36648 36536 36768 36564
rect 36648 35873 36676 36536
rect 36832 36378 36860 36722
rect 36728 36372 36780 36378
rect 36728 36314 36780 36320
rect 36820 36372 36872 36378
rect 36820 36314 36872 36320
rect 36740 36174 36768 36314
rect 36818 36272 36874 36281
rect 36818 36207 36874 36216
rect 36832 36174 36860 36207
rect 36728 36168 36780 36174
rect 36726 36136 36728 36145
rect 36820 36168 36872 36174
rect 36780 36136 36782 36145
rect 36820 36110 36872 36116
rect 36726 36071 36782 36080
rect 36634 35864 36690 35873
rect 36634 35799 36690 35808
rect 36648 35494 36676 35799
rect 36740 35698 36768 36071
rect 36818 36000 36874 36009
rect 36818 35935 36874 35944
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 36636 35488 36688 35494
rect 36636 35430 36688 35436
rect 36740 35086 36768 35634
rect 36832 35630 36860 35935
rect 36820 35624 36872 35630
rect 36820 35566 36872 35572
rect 36924 35154 36952 36740
rect 37004 36644 37056 36650
rect 37004 36586 37056 36592
rect 37016 35290 37044 36586
rect 37004 35284 37056 35290
rect 37004 35226 37056 35232
rect 36820 35148 36872 35154
rect 36820 35090 36872 35096
rect 36912 35148 36964 35154
rect 36912 35090 36964 35096
rect 36728 35080 36780 35086
rect 36728 35022 36780 35028
rect 36832 34610 36860 35090
rect 36728 34604 36780 34610
rect 36728 34546 36780 34552
rect 36820 34604 36872 34610
rect 36820 34546 36872 34552
rect 36542 33552 36598 33561
rect 36542 33487 36598 33496
rect 36636 33516 36688 33522
rect 36636 33458 36688 33464
rect 36648 33017 36676 33458
rect 36740 33096 36768 34546
rect 36912 33992 36964 33998
rect 36912 33934 36964 33940
rect 36820 33108 36872 33114
rect 36740 33068 36820 33096
rect 36820 33050 36872 33056
rect 36634 33008 36690 33017
rect 36634 32943 36690 32952
rect 36360 32360 36412 32366
rect 36360 32302 36412 32308
rect 36452 32360 36504 32366
rect 36452 32302 36504 32308
rect 36188 31726 36308 31754
rect 36084 31204 36136 31210
rect 36084 31146 36136 31152
rect 35992 29844 36044 29850
rect 35992 29786 36044 29792
rect 35912 29702 36032 29730
rect 35900 29028 35952 29034
rect 35900 28970 35952 28976
rect 35912 28762 35940 28970
rect 35900 28756 35952 28762
rect 35900 28698 35952 28704
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 35532 27396 35584 27402
rect 35532 27338 35584 27344
rect 35544 25430 35572 27338
rect 35532 25424 35584 25430
rect 35532 25366 35584 25372
rect 35348 25220 35400 25226
rect 35452 25214 35572 25242
rect 35348 25162 35400 25168
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 35072 24676 35124 24682
rect 35072 24618 35124 24624
rect 35256 24676 35308 24682
rect 35256 24618 35308 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24410 35388 24754
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 34716 23186 34744 23734
rect 35268 23474 35296 24006
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 35360 23662 35388 23802
rect 35452 23730 35480 25094
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 35348 23656 35400 23662
rect 35348 23598 35400 23604
rect 35440 23588 35492 23594
rect 35440 23530 35492 23536
rect 35268 23446 35388 23474
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34796 23112 34848 23118
rect 34796 23054 34848 23060
rect 34980 23112 35032 23118
rect 34980 23054 35032 23060
rect 34808 22778 34836 23054
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 34808 22234 34836 22714
rect 34900 22438 34928 22714
rect 34992 22438 35020 23054
rect 34888 22432 34940 22438
rect 34888 22374 34940 22380
rect 34980 22432 35032 22438
rect 34980 22374 35032 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 35164 22228 35216 22234
rect 35164 22170 35216 22176
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34532 21542 34652 21570
rect 35176 21554 35204 22170
rect 34336 21140 34388 21146
rect 34336 21082 34388 21088
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33520 19446 33548 20334
rect 33888 20058 33916 20402
rect 34624 20398 34652 21542
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 35164 21548 35216 21554
rect 35164 21490 35216 21496
rect 34808 20602 34836 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 20641 35388 23446
rect 35452 23361 35480 23530
rect 35438 23352 35494 23361
rect 35438 23287 35494 23296
rect 35544 22658 35572 25214
rect 35636 24818 35664 27406
rect 35820 27130 35848 28494
rect 35912 28218 35940 28494
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 36004 28014 36032 29702
rect 36188 29646 36216 31726
rect 36268 31136 36320 31142
rect 36268 31078 36320 31084
rect 36280 30734 36308 31078
rect 36268 30728 36320 30734
rect 36268 30670 36320 30676
rect 36176 29640 36228 29646
rect 36096 29600 36176 29628
rect 35992 28008 36044 28014
rect 35992 27950 36044 27956
rect 36004 27384 36032 27950
rect 35912 27356 36032 27384
rect 35808 27124 35860 27130
rect 35808 27066 35860 27072
rect 35808 26852 35860 26858
rect 35808 26794 35860 26800
rect 35716 26444 35768 26450
rect 35716 26386 35768 26392
rect 35624 24812 35676 24818
rect 35624 24754 35676 24760
rect 35624 24676 35676 24682
rect 35624 24618 35676 24624
rect 35636 23662 35664 24618
rect 35728 24614 35756 26386
rect 35820 26246 35848 26794
rect 35912 26246 35940 27356
rect 35990 27296 36046 27305
rect 35990 27231 36046 27240
rect 35808 26240 35860 26246
rect 35808 26182 35860 26188
rect 35900 26240 35952 26246
rect 35900 26182 35952 26188
rect 35820 25838 35848 26182
rect 36004 25974 36032 27231
rect 35992 25968 36044 25974
rect 35992 25910 36044 25916
rect 35808 25832 35860 25838
rect 35808 25774 35860 25780
rect 35900 25424 35952 25430
rect 35900 25366 35952 25372
rect 35912 24886 35940 25366
rect 35900 24880 35952 24886
rect 36004 24857 36032 25910
rect 35900 24822 35952 24828
rect 35990 24848 36046 24857
rect 35716 24608 35768 24614
rect 35716 24550 35768 24556
rect 35728 24342 35756 24550
rect 35912 24410 35940 24822
rect 35990 24783 36046 24792
rect 35992 24744 36044 24750
rect 35992 24686 36044 24692
rect 35808 24404 35860 24410
rect 35808 24346 35860 24352
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35716 24336 35768 24342
rect 35716 24278 35768 24284
rect 35716 23724 35768 23730
rect 35716 23666 35768 23672
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35624 23044 35676 23050
rect 35624 22986 35676 22992
rect 35452 22630 35572 22658
rect 35636 22642 35664 22986
rect 35624 22636 35676 22642
rect 35452 22234 35480 22630
rect 35624 22578 35676 22584
rect 35636 22522 35664 22578
rect 35544 22494 35664 22522
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35544 22094 35572 22494
rect 35624 22094 35676 22098
rect 35544 22092 35676 22094
rect 35544 22066 35624 22092
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35452 20806 35480 21490
rect 35544 21350 35572 22066
rect 35624 22034 35676 22040
rect 35728 21622 35756 23666
rect 35820 23594 35848 24346
rect 35808 23588 35860 23594
rect 35808 23530 35860 23536
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35912 22642 35940 23462
rect 36004 23118 36032 24686
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 36096 22794 36124 29600
rect 36176 29582 36228 29588
rect 36176 28552 36228 28558
rect 36176 28494 36228 28500
rect 36188 27130 36216 28494
rect 36176 27124 36228 27130
rect 36176 27066 36228 27072
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 36188 26382 36216 26862
rect 36176 26376 36228 26382
rect 36176 26318 36228 26324
rect 36004 22766 36124 22794
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 35808 22568 35860 22574
rect 36004 22522 36032 22766
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35808 22510 35860 22516
rect 35820 22166 35848 22510
rect 35912 22494 36032 22522
rect 35912 22438 35940 22494
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 35808 22160 35860 22166
rect 35808 22102 35860 22108
rect 35716 21616 35768 21622
rect 35716 21558 35768 21564
rect 35808 21548 35860 21554
rect 35808 21490 35860 21496
rect 35716 21480 35768 21486
rect 35716 21422 35768 21428
rect 35532 21344 35584 21350
rect 35532 21286 35584 21292
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35544 20942 35572 21286
rect 35636 21010 35664 21286
rect 35624 21004 35676 21010
rect 35624 20946 35676 20952
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 35440 20800 35492 20806
rect 35440 20742 35492 20748
rect 35346 20632 35402 20641
rect 34796 20596 34848 20602
rect 35346 20567 35402 20576
rect 34796 20538 34848 20544
rect 34612 20392 34664 20398
rect 34612 20334 34664 20340
rect 34612 20256 34664 20262
rect 34612 20198 34664 20204
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 33876 20052 33928 20058
rect 33876 19994 33928 20000
rect 34624 19990 34652 20198
rect 34612 19984 34664 19990
rect 34612 19926 34664 19932
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 33508 19440 33560 19446
rect 33980 19417 34008 19450
rect 33508 19382 33560 19388
rect 33966 19408 34022 19417
rect 33966 19343 34022 19352
rect 34060 19372 34112 19378
rect 33336 18822 33732 18850
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 32968 18222 32996 18702
rect 33048 18352 33100 18358
rect 33048 18294 33100 18300
rect 32956 18216 33008 18222
rect 32956 18158 33008 18164
rect 32968 17762 32996 18158
rect 33060 17882 33088 18294
rect 33612 18222 33640 18702
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33048 17876 33100 17882
rect 33048 17818 33100 17824
rect 32968 17734 33088 17762
rect 33060 17678 33088 17734
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 33048 17672 33100 17678
rect 33048 17614 33100 17620
rect 32876 17338 32904 17614
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 32864 16516 32916 16522
rect 32864 16458 32916 16464
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32784 15570 32812 15846
rect 32876 15706 32904 16458
rect 33428 16114 33456 16730
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 33244 15978 33272 16050
rect 33232 15972 33284 15978
rect 33232 15914 33284 15920
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 32864 15700 32916 15706
rect 32864 15642 32916 15648
rect 33152 15638 33180 15846
rect 33140 15632 33192 15638
rect 33140 15574 33192 15580
rect 32772 15564 32824 15570
rect 32772 15506 32824 15512
rect 32864 15564 32916 15570
rect 32864 15506 32916 15512
rect 32772 15088 32824 15094
rect 32772 15030 32824 15036
rect 32784 14414 32812 15030
rect 32772 14408 32824 14414
rect 32772 14350 32824 14356
rect 32784 13870 32812 14350
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 32876 12782 32904 15506
rect 33244 15026 33272 15914
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33520 15337 33548 15438
rect 33506 15328 33562 15337
rect 33506 15263 33562 15272
rect 33324 15088 33376 15094
rect 33322 15056 33324 15065
rect 33376 15056 33378 15065
rect 33232 15020 33284 15026
rect 33322 14991 33378 15000
rect 33232 14962 33284 14968
rect 33048 14340 33100 14346
rect 33048 14282 33100 14288
rect 33060 14006 33088 14282
rect 33048 14000 33100 14006
rect 33048 13942 33100 13948
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33152 13462 33180 13670
rect 33244 13462 33272 14962
rect 33416 14816 33468 14822
rect 33416 14758 33468 14764
rect 33322 14240 33378 14249
rect 33322 14175 33378 14184
rect 33140 13456 33192 13462
rect 33140 13398 33192 13404
rect 33232 13456 33284 13462
rect 33232 13398 33284 13404
rect 32956 13184 33008 13190
rect 32956 13126 33008 13132
rect 32968 12986 32996 13126
rect 33336 12986 33364 14175
rect 33428 14006 33456 14758
rect 33508 14408 33560 14414
rect 33508 14350 33560 14356
rect 33520 14006 33548 14350
rect 33416 14000 33468 14006
rect 33416 13942 33468 13948
rect 33508 14000 33560 14006
rect 33508 13942 33560 13948
rect 32956 12980 33008 12986
rect 32956 12922 33008 12928
rect 33324 12980 33376 12986
rect 33324 12922 33376 12928
rect 32864 12776 32916 12782
rect 32864 12718 32916 12724
rect 32772 12708 32824 12714
rect 32772 12650 32824 12656
rect 32784 12102 32812 12650
rect 32876 12306 32904 12718
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 32784 11762 32812 12038
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 33336 11694 33364 12922
rect 33324 11688 33376 11694
rect 33324 11630 33376 11636
rect 32862 11384 32918 11393
rect 32862 11319 32918 11328
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 32876 10606 32904 11319
rect 33612 11218 33640 18158
rect 33600 11212 33652 11218
rect 33600 11154 33652 11160
rect 33704 11082 33732 18822
rect 33980 18766 34008 19343
rect 34060 19314 34112 19320
rect 34072 18970 34100 19314
rect 34060 18964 34112 18970
rect 34060 18906 34112 18912
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 34624 18426 34652 19926
rect 34716 19786 34744 20198
rect 34808 19922 34836 20538
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34888 20052 34940 20058
rect 34888 19994 34940 20000
rect 34796 19916 34848 19922
rect 34796 19858 34848 19864
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34900 19258 34928 19994
rect 34808 19230 34928 19258
rect 34808 18698 34836 19230
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18692 34848 18698
rect 34796 18634 34848 18640
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34612 18420 34664 18426
rect 34612 18362 34664 18368
rect 34716 18290 34744 18566
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34440 18154 34468 18226
rect 34428 18148 34480 18154
rect 34428 18090 34480 18096
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34532 17746 34560 18022
rect 34612 17876 34664 17882
rect 34612 17818 34664 17824
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34152 17672 34204 17678
rect 34152 17614 34204 17620
rect 34336 17672 34388 17678
rect 34336 17614 34388 17620
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34164 16561 34192 17614
rect 34348 17134 34376 17614
rect 34440 17202 34468 17614
rect 34532 17270 34560 17682
rect 34520 17264 34572 17270
rect 34520 17206 34572 17212
rect 34624 17202 34652 17818
rect 34428 17196 34480 17202
rect 34428 17138 34480 17144
rect 34612 17196 34664 17202
rect 34612 17138 34664 17144
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34336 16584 34388 16590
rect 34150 16552 34206 16561
rect 33784 16516 33836 16522
rect 34336 16526 34388 16532
rect 34150 16487 34206 16496
rect 33784 16458 33836 16464
rect 33796 14822 33824 16458
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33888 14634 33916 16050
rect 34348 16046 34376 16526
rect 34440 16454 34468 17138
rect 34612 16992 34664 16998
rect 34612 16934 34664 16940
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 34624 16182 34652 16934
rect 34612 16176 34664 16182
rect 34612 16118 34664 16124
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34244 15496 34296 15502
rect 34244 15438 34296 15444
rect 34520 15496 34572 15502
rect 34520 15438 34572 15444
rect 34152 15360 34204 15366
rect 34152 15302 34204 15308
rect 33796 14606 33916 14634
rect 33796 14278 33824 14606
rect 33876 14340 33928 14346
rect 33876 14282 33928 14288
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33796 13326 33824 14214
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 33888 12102 33916 14282
rect 34164 14074 34192 15302
rect 34152 14068 34204 14074
rect 34152 14010 34204 14016
rect 34060 12300 34112 12306
rect 34060 12242 34112 12248
rect 33876 12096 33928 12102
rect 33876 12038 33928 12044
rect 34072 11762 34100 12242
rect 34164 12238 34192 14010
rect 34256 13462 34284 15438
rect 34532 14958 34560 15438
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34532 14618 34560 14894
rect 34624 14890 34652 15846
rect 34716 15502 34744 18226
rect 34808 17542 34836 18634
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35072 16788 35124 16794
rect 35072 16730 35124 16736
rect 35084 16674 35112 16730
rect 34980 16652 35032 16658
rect 35084 16646 35204 16674
rect 34980 16594 35032 16600
rect 34888 16516 34940 16522
rect 34888 16458 34940 16464
rect 34900 16425 34928 16458
rect 34886 16416 34942 16425
rect 34886 16351 34942 16360
rect 34992 16250 35020 16594
rect 35176 16590 35204 16646
rect 35164 16584 35216 16590
rect 35256 16584 35308 16590
rect 35164 16526 35216 16532
rect 35254 16552 35256 16561
rect 35308 16552 35310 16561
rect 34980 16244 35032 16250
rect 34980 16186 35032 16192
rect 34992 15978 35020 16186
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 34980 15972 35032 15978
rect 34980 15914 35032 15920
rect 34808 15688 34836 15914
rect 35176 15910 35204 16526
rect 35254 16487 35310 16496
rect 35164 15904 35216 15910
rect 35164 15846 35216 15852
rect 35268 15858 35296 16487
rect 35360 16454 35388 20402
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 35348 16448 35400 16454
rect 35348 16390 35400 16396
rect 35268 15830 35388 15858
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34808 15660 34928 15688
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 15088 34756 15094
rect 34704 15030 34756 15036
rect 34612 14884 34664 14890
rect 34612 14826 34664 14832
rect 34520 14612 34572 14618
rect 34520 14554 34572 14560
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34244 13456 34296 13462
rect 34244 13398 34296 13404
rect 34440 13394 34468 14010
rect 34716 13870 34744 15030
rect 34704 13864 34756 13870
rect 34704 13806 34756 13812
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 34440 12850 34468 13330
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34336 12640 34388 12646
rect 34336 12582 34388 12588
rect 34348 12238 34376 12582
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34532 11898 34560 13194
rect 34716 12832 34744 13670
rect 34808 13530 34836 15370
rect 34900 15026 34928 15660
rect 35360 15570 35388 15830
rect 35348 15564 35400 15570
rect 35348 15506 35400 15512
rect 35072 15088 35124 15094
rect 35072 15030 35124 15036
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 35084 14929 35112 15030
rect 35070 14920 35126 14929
rect 35070 14855 35126 14864
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35072 14612 35124 14618
rect 35072 14554 35124 14560
rect 35084 14521 35112 14554
rect 35070 14512 35126 14521
rect 35070 14447 35126 14456
rect 35360 14346 35388 15506
rect 35452 15162 35480 19654
rect 35544 18970 35572 20878
rect 35624 20256 35676 20262
rect 35624 20198 35676 20204
rect 35636 18970 35664 20198
rect 35532 18964 35584 18970
rect 35532 18906 35584 18912
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35624 18760 35676 18766
rect 35624 18702 35676 18708
rect 35636 18358 35664 18702
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 35532 16788 35584 16794
rect 35532 16730 35584 16736
rect 35544 15502 35572 16730
rect 35636 16454 35664 18294
rect 35728 18154 35756 21422
rect 35820 21146 35848 21490
rect 35912 21350 35940 22374
rect 36004 21554 36032 22374
rect 36096 22098 36124 22578
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 36084 21956 36136 21962
rect 36084 21898 36136 21904
rect 36096 21690 36124 21898
rect 36084 21684 36136 21690
rect 36084 21626 36136 21632
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35912 20874 35940 21082
rect 36004 21010 36032 21490
rect 35992 21004 36044 21010
rect 35992 20946 36044 20952
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35820 19666 35848 20742
rect 36188 20398 36216 26318
rect 36280 25294 36308 30670
rect 36372 30161 36400 32302
rect 36648 31346 36676 32943
rect 36832 31929 36860 33050
rect 36818 31920 36874 31929
rect 36818 31855 36874 31864
rect 36636 31340 36688 31346
rect 36636 31282 36688 31288
rect 36452 31272 36504 31278
rect 36452 31214 36504 31220
rect 36464 31113 36492 31214
rect 36450 31104 36506 31113
rect 36450 31039 36506 31048
rect 36648 30938 36676 31282
rect 36728 31136 36780 31142
rect 36728 31078 36780 31084
rect 36636 30932 36688 30938
rect 36636 30874 36688 30880
rect 36544 30796 36596 30802
rect 36544 30738 36596 30744
rect 36452 30184 36504 30190
rect 36358 30152 36414 30161
rect 36452 30126 36504 30132
rect 36358 30087 36414 30096
rect 36464 30025 36492 30126
rect 36450 30016 36506 30025
rect 36450 29951 36506 29960
rect 36358 29064 36414 29073
rect 36358 28999 36414 29008
rect 36372 28218 36400 28999
rect 36556 28422 36584 30738
rect 36636 30660 36688 30666
rect 36636 30602 36688 30608
rect 36544 28416 36596 28422
rect 36544 28358 36596 28364
rect 36360 28212 36412 28218
rect 36360 28154 36412 28160
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36360 27668 36412 27674
rect 36360 27610 36412 27616
rect 36372 27577 36400 27610
rect 36358 27568 36414 27577
rect 36358 27503 36360 27512
rect 36412 27503 36414 27512
rect 36360 27474 36412 27480
rect 36464 27334 36492 28018
rect 36556 27554 36584 28358
rect 36648 27674 36676 30602
rect 36740 29578 36768 31078
rect 36820 30932 36872 30938
rect 36820 30874 36872 30880
rect 36728 29572 36780 29578
rect 36728 29514 36780 29520
rect 36636 27668 36688 27674
rect 36636 27610 36688 27616
rect 36556 27526 36768 27554
rect 36544 27464 36596 27470
rect 36544 27406 36596 27412
rect 36360 27328 36412 27334
rect 36360 27270 36412 27276
rect 36452 27328 36504 27334
rect 36452 27270 36504 27276
rect 36372 26994 36400 27270
rect 36360 26988 36412 26994
rect 36360 26930 36412 26936
rect 36464 26874 36492 27270
rect 36556 27130 36584 27406
rect 36544 27124 36596 27130
rect 36544 27066 36596 27072
rect 36636 26920 36688 26926
rect 36464 26846 36584 26874
rect 36636 26862 36688 26868
rect 36452 26784 36504 26790
rect 36452 26726 36504 26732
rect 36464 25974 36492 26726
rect 36452 25968 36504 25974
rect 36452 25910 36504 25916
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 36372 24426 36400 25638
rect 36464 24614 36492 25910
rect 36556 24818 36584 26846
rect 36648 26382 36676 26862
rect 36636 26376 36688 26382
rect 36636 26318 36688 26324
rect 36636 25288 36688 25294
rect 36636 25230 36688 25236
rect 36648 24818 36676 25230
rect 36740 25226 36768 27526
rect 36832 25362 36860 30874
rect 36924 29850 36952 33934
rect 37016 33522 37044 35226
rect 37108 33930 37136 37334
rect 37188 37188 37240 37194
rect 37188 37130 37240 37136
rect 37200 35873 37228 37130
rect 37280 36304 37332 36310
rect 37280 36246 37332 36252
rect 37292 36174 37320 36246
rect 37280 36168 37332 36174
rect 37280 36110 37332 36116
rect 37186 35864 37242 35873
rect 37186 35799 37242 35808
rect 37188 35760 37240 35766
rect 37188 35702 37240 35708
rect 37200 35222 37228 35702
rect 37292 35494 37320 36110
rect 37464 36032 37516 36038
rect 37462 36000 37464 36009
rect 37516 36000 37518 36009
rect 37462 35935 37518 35944
rect 37568 35680 37596 39782
rect 37660 39250 37688 41386
rect 37752 41138 37780 41414
rect 37740 41132 37792 41138
rect 37740 41074 37792 41080
rect 37936 40526 37964 42298
rect 38384 42220 38436 42226
rect 38384 42162 38436 42168
rect 38200 42152 38252 42158
rect 38200 42094 38252 42100
rect 37740 40520 37792 40526
rect 37924 40520 37976 40526
rect 37792 40468 37872 40474
rect 37740 40462 37872 40468
rect 37924 40462 37976 40468
rect 37752 40446 37872 40462
rect 37660 39222 37780 39250
rect 37648 39092 37700 39098
rect 37648 39034 37700 39040
rect 37660 38350 37688 39034
rect 37648 38344 37700 38350
rect 37648 38286 37700 38292
rect 37648 36780 37700 36786
rect 37648 36722 37700 36728
rect 37660 35698 37688 36722
rect 37752 36582 37780 39222
rect 37844 38350 37872 40446
rect 37936 40186 37964 40462
rect 37924 40180 37976 40186
rect 37924 40122 37976 40128
rect 38108 39840 38160 39846
rect 38028 39800 38108 39828
rect 38028 39438 38056 39800
rect 38108 39782 38160 39788
rect 38016 39432 38068 39438
rect 38014 39400 38016 39409
rect 38068 39400 38070 39409
rect 38014 39335 38070 39344
rect 37832 38344 37884 38350
rect 37832 38286 37884 38292
rect 37740 36576 37792 36582
rect 37740 36518 37792 36524
rect 37752 36310 37780 36518
rect 37844 36417 37872 38286
rect 37924 38276 37976 38282
rect 37924 38218 37976 38224
rect 37936 37233 37964 38218
rect 38212 37738 38240 42094
rect 38396 42022 38424 42162
rect 38384 42016 38436 42022
rect 38384 41958 38436 41964
rect 38396 41478 38424 41958
rect 38660 41608 38712 41614
rect 38660 41550 38712 41556
rect 38384 41472 38436 41478
rect 38384 41414 38436 41420
rect 38396 41386 38516 41414
rect 38384 40656 38436 40662
rect 38384 40598 38436 40604
rect 38200 37732 38252 37738
rect 38200 37674 38252 37680
rect 38108 37256 38160 37262
rect 37922 37224 37978 37233
rect 38108 37198 38160 37204
rect 38200 37256 38252 37262
rect 38200 37198 38252 37204
rect 38292 37256 38344 37262
rect 38292 37198 38344 37204
rect 37922 37159 37978 37168
rect 37936 36650 37964 37159
rect 37924 36644 37976 36650
rect 37924 36586 37976 36592
rect 38016 36644 38068 36650
rect 38016 36586 38068 36592
rect 37830 36408 37886 36417
rect 37830 36343 37886 36352
rect 37740 36304 37792 36310
rect 37740 36246 37792 36252
rect 38028 36174 38056 36586
rect 38120 36582 38148 37198
rect 38212 36922 38240 37198
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 38304 36854 38332 37198
rect 38292 36848 38344 36854
rect 38292 36790 38344 36796
rect 38396 36786 38424 40598
rect 38488 40050 38516 41386
rect 38672 40730 38700 41550
rect 38856 41154 38884 44200
rect 39304 42084 39356 42090
rect 39304 42026 39356 42032
rect 38936 42016 38988 42022
rect 38936 41958 38988 41964
rect 38948 41414 38976 41958
rect 39316 41478 39344 42026
rect 39396 41744 39448 41750
rect 39396 41686 39448 41692
rect 39304 41472 39356 41478
rect 39304 41414 39356 41420
rect 38948 41386 39252 41414
rect 38856 41126 39068 41154
rect 38844 41064 38896 41070
rect 38844 41006 38896 41012
rect 38752 40928 38804 40934
rect 38752 40870 38804 40876
rect 38660 40724 38712 40730
rect 38660 40666 38712 40672
rect 38764 40390 38792 40870
rect 38752 40384 38804 40390
rect 38752 40326 38804 40332
rect 38476 40044 38528 40050
rect 38476 39986 38528 39992
rect 38568 39296 38620 39302
rect 38568 39238 38620 39244
rect 38476 38208 38528 38214
rect 38476 38150 38528 38156
rect 38488 37874 38516 38150
rect 38476 37868 38528 37874
rect 38476 37810 38528 37816
rect 38488 37262 38516 37810
rect 38476 37256 38528 37262
rect 38476 37198 38528 37204
rect 38384 36780 38436 36786
rect 38384 36722 38436 36728
rect 38108 36576 38160 36582
rect 38108 36518 38160 36524
rect 37740 36168 37792 36174
rect 37738 36136 37740 36145
rect 38016 36168 38068 36174
rect 37792 36136 37794 36145
rect 38016 36110 38068 36116
rect 37738 36071 37794 36080
rect 37476 35652 37596 35680
rect 37648 35692 37700 35698
rect 37280 35488 37332 35494
rect 37280 35430 37332 35436
rect 37188 35216 37240 35222
rect 37188 35158 37240 35164
rect 37188 34400 37240 34406
rect 37188 34342 37240 34348
rect 37280 34400 37332 34406
rect 37280 34342 37332 34348
rect 37200 34134 37228 34342
rect 37188 34128 37240 34134
rect 37188 34070 37240 34076
rect 37096 33924 37148 33930
rect 37096 33866 37148 33872
rect 37188 33856 37240 33862
rect 37188 33798 37240 33804
rect 37004 33516 37056 33522
rect 37004 33458 37056 33464
rect 37200 32502 37228 33798
rect 37188 32496 37240 32502
rect 37188 32438 37240 32444
rect 37096 32360 37148 32366
rect 37096 32302 37148 32308
rect 37002 32056 37058 32065
rect 37108 32026 37136 32302
rect 37002 31991 37058 32000
rect 37096 32020 37148 32026
rect 37016 31822 37044 31991
rect 37096 31962 37148 31968
rect 37188 31952 37240 31958
rect 37188 31894 37240 31900
rect 37004 31816 37056 31822
rect 37002 31784 37004 31793
rect 37056 31784 37058 31793
rect 37002 31719 37058 31728
rect 37004 31408 37056 31414
rect 37002 31376 37004 31385
rect 37056 31376 37058 31385
rect 37002 31311 37058 31320
rect 37004 30320 37056 30326
rect 37004 30262 37056 30268
rect 37016 29850 37044 30262
rect 36912 29844 36964 29850
rect 36912 29786 36964 29792
rect 37004 29844 37056 29850
rect 37004 29786 37056 29792
rect 37200 29730 37228 31894
rect 37292 31482 37320 34342
rect 37476 33386 37504 35652
rect 37700 35652 37964 35680
rect 37648 35634 37700 35640
rect 37832 35556 37884 35562
rect 37832 35498 37884 35504
rect 37844 35018 37872 35498
rect 37832 35012 37884 35018
rect 37832 34954 37884 34960
rect 37738 34912 37794 34921
rect 37738 34847 37794 34856
rect 37752 34610 37780 34847
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 37648 34604 37700 34610
rect 37648 34546 37700 34552
rect 37740 34604 37792 34610
rect 37740 34546 37792 34552
rect 37568 34406 37596 34546
rect 37556 34400 37608 34406
rect 37556 34342 37608 34348
rect 37660 33998 37688 34546
rect 37648 33992 37700 33998
rect 37648 33934 37700 33940
rect 37740 33652 37792 33658
rect 37740 33594 37792 33600
rect 37648 33584 37700 33590
rect 37648 33526 37700 33532
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 37464 33380 37516 33386
rect 37464 33322 37516 33328
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 37384 32337 37412 32846
rect 37462 32736 37518 32745
rect 37462 32671 37518 32680
rect 37476 32570 37504 32671
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37370 32328 37426 32337
rect 37370 32263 37426 32272
rect 37280 31476 37332 31482
rect 37280 31418 37332 31424
rect 37372 31272 37424 31278
rect 37372 31214 37424 31220
rect 37280 31204 37332 31210
rect 37280 31146 37332 31152
rect 37292 30734 37320 31146
rect 37280 30728 37332 30734
rect 37280 30670 37332 30676
rect 37384 30598 37412 31214
rect 37568 30938 37596 33458
rect 37660 33318 37688 33526
rect 37752 33386 37780 33594
rect 37740 33380 37792 33386
rect 37740 33322 37792 33328
rect 37648 33312 37700 33318
rect 37648 33254 37700 33260
rect 37752 33114 37780 33322
rect 37844 33300 37872 34954
rect 37936 34610 37964 35652
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 38028 34134 38056 36110
rect 38120 35737 38148 36518
rect 38382 36408 38438 36417
rect 38382 36343 38438 36352
rect 38200 36304 38252 36310
rect 38200 36246 38252 36252
rect 38212 36174 38240 36246
rect 38200 36168 38252 36174
rect 38200 36110 38252 36116
rect 38292 36168 38344 36174
rect 38292 36110 38344 36116
rect 38106 35728 38162 35737
rect 38106 35663 38162 35672
rect 38200 35488 38252 35494
rect 38304 35476 38332 36110
rect 38252 35448 38332 35476
rect 38200 35430 38252 35436
rect 38212 35086 38240 35430
rect 38292 35148 38344 35154
rect 38292 35090 38344 35096
rect 38200 35080 38252 35086
rect 38200 35022 38252 35028
rect 38108 34672 38160 34678
rect 38108 34614 38160 34620
rect 38016 34128 38068 34134
rect 38016 34070 38068 34076
rect 38016 33924 38068 33930
rect 38016 33866 38068 33872
rect 37924 33856 37976 33862
rect 37924 33798 37976 33804
rect 37936 33425 37964 33798
rect 38028 33697 38056 33866
rect 38120 33862 38148 34614
rect 38108 33856 38160 33862
rect 38108 33798 38160 33804
rect 38014 33688 38070 33697
rect 38212 33674 38240 35022
rect 38304 34542 38332 35090
rect 38292 34536 38344 34542
rect 38292 34478 38344 34484
rect 38014 33623 38070 33632
rect 38120 33646 38240 33674
rect 37922 33416 37978 33425
rect 37922 33351 37978 33360
rect 37844 33272 37964 33300
rect 37648 33108 37700 33114
rect 37648 33050 37700 33056
rect 37740 33108 37792 33114
rect 37740 33050 37792 33056
rect 37660 32978 37688 33050
rect 37648 32972 37700 32978
rect 37648 32914 37700 32920
rect 37648 32768 37700 32774
rect 37648 32710 37700 32716
rect 37660 32026 37688 32710
rect 37832 32428 37884 32434
rect 37832 32370 37884 32376
rect 37844 32026 37872 32370
rect 37648 32020 37700 32026
rect 37648 31962 37700 31968
rect 37832 32020 37884 32026
rect 37832 31962 37884 31968
rect 37740 31884 37792 31890
rect 37740 31826 37792 31832
rect 37648 31136 37700 31142
rect 37648 31078 37700 31084
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37372 30592 37424 30598
rect 37372 30534 37424 30540
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37016 29714 37228 29730
rect 37004 29708 37228 29714
rect 37056 29702 37228 29708
rect 37004 29650 37056 29656
rect 37292 29646 37320 30194
rect 37096 29640 37148 29646
rect 37280 29640 37332 29646
rect 37148 29600 37228 29628
rect 37096 29582 37148 29588
rect 37004 29572 37056 29578
rect 37004 29514 37056 29520
rect 37016 29306 37044 29514
rect 37200 29510 37228 29600
rect 37280 29582 37332 29588
rect 37188 29504 37240 29510
rect 37188 29446 37240 29452
rect 37004 29300 37056 29306
rect 37004 29242 37056 29248
rect 37016 28762 37044 29242
rect 37004 28756 37056 28762
rect 37004 28698 37056 28704
rect 36912 28416 36964 28422
rect 36912 28358 36964 28364
rect 36924 27878 36952 28358
rect 37096 28144 37148 28150
rect 37096 28086 37148 28092
rect 37004 28008 37056 28014
rect 37004 27950 37056 27956
rect 36912 27872 36964 27878
rect 36912 27814 36964 27820
rect 37016 27470 37044 27950
rect 37108 27606 37136 28086
rect 37096 27600 37148 27606
rect 37096 27542 37148 27548
rect 37004 27464 37056 27470
rect 37004 27406 37056 27412
rect 37108 27062 37136 27542
rect 37096 27056 37148 27062
rect 37096 26998 37148 27004
rect 37004 26852 37056 26858
rect 37004 26794 37056 26800
rect 37016 26450 37044 26794
rect 37108 26586 37136 26998
rect 37096 26580 37148 26586
rect 37096 26522 37148 26528
rect 37004 26444 37056 26450
rect 37004 26386 37056 26392
rect 36820 25356 36872 25362
rect 36820 25298 36872 25304
rect 36728 25220 36780 25226
rect 36728 25162 36780 25168
rect 37094 24848 37150 24857
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 36636 24812 36688 24818
rect 37094 24783 37150 24792
rect 36636 24754 36688 24760
rect 37108 24750 37136 24783
rect 37096 24744 37148 24750
rect 37096 24686 37148 24692
rect 36452 24608 36504 24614
rect 36452 24550 36504 24556
rect 36912 24608 36964 24614
rect 36912 24550 36964 24556
rect 36372 24398 36492 24426
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36280 24041 36308 24142
rect 36266 24032 36322 24041
rect 36266 23967 36322 23976
rect 36268 23724 36320 23730
rect 36372 23712 36400 24142
rect 36464 24070 36492 24398
rect 36544 24404 36596 24410
rect 36544 24346 36596 24352
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36320 23684 36400 23712
rect 36268 23666 36320 23672
rect 36266 23624 36322 23633
rect 36266 23559 36322 23568
rect 36280 22982 36308 23559
rect 36268 22976 36320 22982
rect 36268 22918 36320 22924
rect 36372 22030 36400 23684
rect 36464 23594 36492 24006
rect 36556 23730 36584 24346
rect 36544 23724 36596 23730
rect 36544 23666 36596 23672
rect 36556 23633 36584 23666
rect 36542 23624 36598 23633
rect 36452 23588 36504 23594
rect 36542 23559 36598 23568
rect 36452 23530 36504 23536
rect 36728 23316 36780 23322
rect 36728 23258 36780 23264
rect 36634 22672 36690 22681
rect 36634 22607 36636 22616
rect 36688 22607 36690 22616
rect 36636 22578 36688 22584
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36452 22160 36504 22166
rect 36452 22102 36504 22108
rect 36360 22024 36412 22030
rect 36360 21966 36412 21972
rect 36372 21078 36400 21966
rect 36360 21072 36412 21078
rect 36360 21014 36412 21020
rect 36176 20392 36228 20398
rect 36176 20334 36228 20340
rect 36464 19938 36492 22102
rect 36556 22098 36584 22374
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 36636 22024 36688 22030
rect 36636 21966 36688 21972
rect 36464 19910 36584 19938
rect 36556 19854 36584 19910
rect 36452 19848 36504 19854
rect 36452 19790 36504 19796
rect 36544 19848 36596 19854
rect 36544 19790 36596 19796
rect 35820 19638 35940 19666
rect 35808 19508 35860 19514
rect 35808 19450 35860 19456
rect 35716 18148 35768 18154
rect 35716 18090 35768 18096
rect 35624 16448 35676 16454
rect 35624 16390 35676 16396
rect 35532 15496 35584 15502
rect 35532 15438 35584 15444
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35544 15042 35572 15438
rect 35624 15428 35676 15434
rect 35624 15370 35676 15376
rect 35452 15014 35572 15042
rect 35348 14340 35400 14346
rect 35348 14282 35400 14288
rect 35164 14272 35216 14278
rect 35216 14232 35296 14260
rect 35164 14214 35216 14220
rect 34888 13932 34940 13938
rect 34888 13874 34940 13880
rect 34900 13802 34928 13874
rect 34888 13796 34940 13802
rect 34888 13738 34940 13744
rect 35268 13682 35296 14232
rect 35452 13734 35480 15014
rect 35532 14884 35584 14890
rect 35532 14826 35584 14832
rect 35544 13938 35572 14826
rect 35636 14521 35664 15370
rect 35622 14512 35678 14521
rect 35622 14447 35678 14456
rect 35624 14000 35676 14006
rect 35624 13942 35676 13948
rect 35532 13932 35584 13938
rect 35532 13874 35584 13880
rect 35440 13728 35492 13734
rect 35268 13654 35388 13682
rect 35440 13670 35492 13676
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 34808 12968 34836 13466
rect 35360 13462 35388 13654
rect 35348 13456 35400 13462
rect 35348 13398 35400 13404
rect 34808 12940 34928 12968
rect 34900 12850 34928 12940
rect 35360 12850 35388 13398
rect 35544 13394 35572 13874
rect 35636 13802 35664 13942
rect 35624 13796 35676 13802
rect 35624 13738 35676 13744
rect 35532 13388 35584 13394
rect 35532 13330 35584 13336
rect 34888 12844 34940 12850
rect 34716 12804 34836 12832
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34624 12102 34652 12718
rect 34704 12708 34756 12714
rect 34704 12650 34756 12656
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34060 11756 34112 11762
rect 34716 11744 34744 12650
rect 34808 12646 34836 12804
rect 34888 12786 34940 12792
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35544 12238 35572 13330
rect 35636 13326 35664 13738
rect 35728 13530 35756 18090
rect 35820 17882 35848 19450
rect 35912 19310 35940 19638
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35900 19304 35952 19310
rect 35900 19246 35952 19252
rect 35808 17876 35860 17882
rect 35808 17818 35860 17824
rect 35912 17610 35940 19246
rect 36004 18698 36032 19314
rect 36464 18970 36492 19790
rect 36452 18964 36504 18970
rect 36452 18906 36504 18912
rect 35992 18692 36044 18698
rect 35992 18634 36044 18640
rect 36360 18624 36412 18630
rect 36360 18566 36412 18572
rect 36372 18154 36400 18566
rect 36464 18426 36492 18906
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36360 18148 36412 18154
rect 36360 18090 36412 18096
rect 36176 18080 36228 18086
rect 36176 18022 36228 18028
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 35912 16046 35940 17546
rect 36188 17338 36216 18022
rect 36268 17876 36320 17882
rect 36268 17818 36320 17824
rect 36280 17746 36308 17818
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 36648 17678 36676 21966
rect 36740 21146 36768 23258
rect 36820 23044 36872 23050
rect 36820 22986 36872 22992
rect 36832 22778 36860 22986
rect 36820 22772 36872 22778
rect 36820 22714 36872 22720
rect 36818 22672 36874 22681
rect 36818 22607 36820 22616
rect 36872 22607 36874 22616
rect 36820 22578 36872 22584
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36740 20058 36768 20878
rect 36728 20052 36780 20058
rect 36728 19994 36780 20000
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36176 17332 36228 17338
rect 36176 17274 36228 17280
rect 35992 17264 36044 17270
rect 35992 17206 36044 17212
rect 36004 16454 36032 17206
rect 36268 16788 36320 16794
rect 36268 16730 36320 16736
rect 35992 16448 36044 16454
rect 35992 16390 36044 16396
rect 36004 16114 36032 16390
rect 36176 16176 36228 16182
rect 36174 16144 36176 16153
rect 36228 16144 36230 16153
rect 35992 16108 36044 16114
rect 36174 16079 36230 16088
rect 35992 16050 36044 16056
rect 35900 16040 35952 16046
rect 35900 15982 35952 15988
rect 35912 15706 35940 15982
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 35900 15088 35952 15094
rect 35898 15056 35900 15065
rect 35952 15056 35954 15065
rect 35898 14991 35954 15000
rect 35806 14920 35862 14929
rect 35806 14855 35862 14864
rect 35820 14414 35848 14855
rect 35900 14544 35952 14550
rect 35900 14486 35952 14492
rect 35808 14408 35860 14414
rect 35808 14350 35860 14356
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 35716 13524 35768 13530
rect 35716 13466 35768 13472
rect 35820 13326 35848 14214
rect 35624 13320 35676 13326
rect 35624 13262 35676 13268
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35636 12918 35664 13262
rect 35624 12912 35676 12918
rect 35624 12854 35676 12860
rect 35532 12232 35584 12238
rect 35532 12174 35584 12180
rect 35912 11898 35940 14486
rect 36004 12782 36032 16050
rect 36280 15570 36308 16730
rect 36452 16516 36504 16522
rect 36452 16458 36504 16464
rect 36268 15564 36320 15570
rect 36268 15506 36320 15512
rect 36084 15428 36136 15434
rect 36084 15370 36136 15376
rect 36096 14074 36124 15370
rect 36280 14822 36308 15506
rect 36464 15026 36492 16458
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36268 14816 36320 14822
rect 36268 14758 36320 14764
rect 36372 14482 36400 14962
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36360 14476 36412 14482
rect 36360 14418 36412 14424
rect 36176 14272 36228 14278
rect 36176 14214 36228 14220
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 34980 11892 35032 11898
rect 34980 11834 35032 11840
rect 35900 11892 35952 11898
rect 35900 11834 35952 11840
rect 34992 11762 35020 11834
rect 36188 11762 36216 14214
rect 36372 13938 36400 14418
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36464 13462 36492 14758
rect 36556 14618 36584 17478
rect 36648 15706 36676 17614
rect 36728 17196 36780 17202
rect 36728 17138 36780 17144
rect 36740 16250 36768 17138
rect 36832 16454 36860 22578
rect 36924 21622 36952 24550
rect 37096 24336 37148 24342
rect 37094 24304 37096 24313
rect 37148 24304 37150 24313
rect 37094 24239 37150 24248
rect 37004 24200 37056 24206
rect 37200 24188 37228 29446
rect 37292 28966 37320 29582
rect 37384 29306 37412 30534
rect 37372 29300 37424 29306
rect 37372 29242 37424 29248
rect 37280 28960 37332 28966
rect 37280 28902 37332 28908
rect 37556 28756 37608 28762
rect 37556 28698 37608 28704
rect 37462 27976 37518 27985
rect 37462 27911 37464 27920
rect 37516 27911 37518 27920
rect 37464 27882 37516 27888
rect 37280 26784 37332 26790
rect 37280 26726 37332 26732
rect 37056 24160 37228 24188
rect 37004 24142 37056 24148
rect 37016 22642 37044 24142
rect 37094 23760 37150 23769
rect 37094 23695 37150 23704
rect 37108 23662 37136 23695
rect 37096 23656 37148 23662
rect 37096 23598 37148 23604
rect 37186 23352 37242 23361
rect 37186 23287 37242 23296
rect 37096 23248 37148 23254
rect 37096 23190 37148 23196
rect 37004 22636 37056 22642
rect 37004 22578 37056 22584
rect 36912 21616 36964 21622
rect 36912 21558 36964 21564
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 36924 19786 36952 20402
rect 36912 19780 36964 19786
rect 36912 19722 36964 19728
rect 36924 19514 36952 19722
rect 36912 19508 36964 19514
rect 36912 19450 36964 19456
rect 36912 18964 36964 18970
rect 36912 18906 36964 18912
rect 36924 17134 36952 18906
rect 36912 17128 36964 17134
rect 36912 17070 36964 17076
rect 36820 16448 36872 16454
rect 36820 16390 36872 16396
rect 36728 16244 36780 16250
rect 36728 16186 36780 16192
rect 36728 15972 36780 15978
rect 36728 15914 36780 15920
rect 36636 15700 36688 15706
rect 36636 15642 36688 15648
rect 36636 15496 36688 15502
rect 36740 15484 36768 15914
rect 36688 15456 36768 15484
rect 36820 15496 36872 15502
rect 36636 15438 36688 15444
rect 36820 15438 36872 15444
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 36452 13456 36504 13462
rect 36452 13398 36504 13404
rect 36648 12306 36676 15438
rect 36726 15328 36782 15337
rect 36726 15263 36782 15272
rect 36740 15026 36768 15263
rect 36832 15162 36860 15438
rect 36820 15156 36872 15162
rect 36820 15098 36872 15104
rect 36728 15020 36780 15026
rect 36728 14962 36780 14968
rect 36728 14884 36780 14890
rect 36728 14826 36780 14832
rect 36740 13870 36768 14826
rect 36820 14340 36872 14346
rect 36820 14282 36872 14288
rect 36728 13864 36780 13870
rect 36728 13806 36780 13812
rect 36832 12986 36860 14282
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 37016 12434 37044 21286
rect 37108 19446 37136 23190
rect 37200 23118 37228 23287
rect 37188 23112 37240 23118
rect 37188 23054 37240 23060
rect 37188 22024 37240 22030
rect 37186 21992 37188 22001
rect 37240 21992 37242 22001
rect 37186 21927 37242 21936
rect 37292 19854 37320 26726
rect 37464 26308 37516 26314
rect 37464 26250 37516 26256
rect 37476 26217 37504 26250
rect 37462 26208 37518 26217
rect 37462 26143 37518 26152
rect 37372 25900 37424 25906
rect 37476 25888 37504 26143
rect 37424 25860 37504 25888
rect 37372 25842 37424 25848
rect 37568 25838 37596 28698
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37370 25528 37426 25537
rect 37370 25463 37372 25472
rect 37424 25463 37426 25472
rect 37372 25434 37424 25440
rect 37372 25220 37424 25226
rect 37372 25162 37424 25168
rect 37384 24410 37412 25162
rect 37464 25152 37516 25158
rect 37464 25094 37516 25100
rect 37476 24410 37504 25094
rect 37554 24712 37610 24721
rect 37554 24647 37610 24656
rect 37372 24404 37424 24410
rect 37372 24346 37424 24352
rect 37464 24404 37516 24410
rect 37464 24346 37516 24352
rect 37476 23662 37504 24346
rect 37464 23656 37516 23662
rect 37464 23598 37516 23604
rect 37464 23520 37516 23526
rect 37464 23462 37516 23468
rect 37476 22030 37504 23462
rect 37568 23118 37596 24647
rect 37660 24206 37688 31078
rect 37752 30938 37780 31826
rect 37740 30932 37792 30938
rect 37740 30874 37792 30880
rect 37936 30326 37964 33272
rect 38120 32042 38148 33646
rect 38304 33522 38332 34478
rect 38396 33998 38424 36343
rect 38476 36032 38528 36038
rect 38476 35974 38528 35980
rect 38488 35766 38516 35974
rect 38476 35760 38528 35766
rect 38476 35702 38528 35708
rect 38476 35080 38528 35086
rect 38476 35022 38528 35028
rect 38488 34626 38516 35022
rect 38580 34746 38608 39238
rect 38660 37256 38712 37262
rect 38764 37244 38792 40326
rect 38856 39982 38884 41006
rect 39040 40390 39068 41126
rect 38936 40384 38988 40390
rect 38936 40326 38988 40332
rect 39028 40384 39080 40390
rect 39028 40326 39080 40332
rect 38844 39976 38896 39982
rect 38844 39918 38896 39924
rect 38856 39370 38884 39918
rect 38844 39364 38896 39370
rect 38844 39306 38896 39312
rect 38856 38894 38884 39306
rect 38948 38978 38976 40326
rect 39120 39432 39172 39438
rect 39120 39374 39172 39380
rect 39132 39030 39160 39374
rect 39120 39024 39172 39030
rect 38948 38950 39068 38978
rect 39120 38966 39172 38972
rect 38844 38888 38896 38894
rect 38844 38830 38896 38836
rect 38712 37216 38792 37244
rect 38660 37198 38712 37204
rect 38672 36650 38700 37198
rect 38660 36644 38712 36650
rect 38660 36586 38712 36592
rect 38752 36372 38804 36378
rect 38752 36314 38804 36320
rect 38764 36174 38792 36314
rect 38752 36168 38804 36174
rect 38752 36110 38804 36116
rect 38568 34740 38620 34746
rect 38568 34682 38620 34688
rect 38488 34598 38608 34626
rect 38476 34400 38528 34406
rect 38476 34342 38528 34348
rect 38384 33992 38436 33998
rect 38384 33934 38436 33940
rect 38488 33862 38516 34342
rect 38384 33856 38436 33862
rect 38384 33798 38436 33804
rect 38476 33856 38528 33862
rect 38476 33798 38528 33804
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38200 32768 38252 32774
rect 38200 32710 38252 32716
rect 38212 32201 38240 32710
rect 38292 32496 38344 32502
rect 38292 32438 38344 32444
rect 38198 32192 38254 32201
rect 38198 32127 38254 32136
rect 38120 32014 38240 32042
rect 38016 31816 38068 31822
rect 38016 31758 38068 31764
rect 37924 30320 37976 30326
rect 37924 30262 37976 30268
rect 37740 30252 37792 30258
rect 37740 30194 37792 30200
rect 37832 30252 37884 30258
rect 37832 30194 37884 30200
rect 37752 29102 37780 30194
rect 37844 29782 37872 30194
rect 37832 29776 37884 29782
rect 37832 29718 37884 29724
rect 37924 29640 37976 29646
rect 37924 29582 37976 29588
rect 37936 29306 37964 29582
rect 37924 29300 37976 29306
rect 37924 29242 37976 29248
rect 37740 29096 37792 29102
rect 37740 29038 37792 29044
rect 37752 27606 37780 29038
rect 37832 28688 37884 28694
rect 37832 28630 37884 28636
rect 37844 27878 37872 28630
rect 37832 27872 37884 27878
rect 37832 27814 37884 27820
rect 37740 27600 37792 27606
rect 37740 27542 37792 27548
rect 37752 26994 37780 27542
rect 37936 27452 37964 29242
rect 38028 28626 38056 31758
rect 38108 31204 38160 31210
rect 38108 31146 38160 31152
rect 38120 31113 38148 31146
rect 38106 31104 38162 31113
rect 38106 31039 38162 31048
rect 38108 30728 38160 30734
rect 38108 30670 38160 30676
rect 38120 30326 38148 30670
rect 38212 30394 38240 32014
rect 38304 31822 38332 32438
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 38292 31340 38344 31346
rect 38292 31282 38344 31288
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 38108 30320 38160 30326
rect 38108 30262 38160 30268
rect 38120 29714 38148 30262
rect 38200 30252 38252 30258
rect 38200 30194 38252 30200
rect 38108 29708 38160 29714
rect 38108 29650 38160 29656
rect 38212 29238 38240 30194
rect 38304 30025 38332 31282
rect 38396 31278 38424 33798
rect 38580 33590 38608 34598
rect 38856 34474 38884 38830
rect 39040 38010 39068 38950
rect 39224 38554 39252 41386
rect 39316 41206 39344 41414
rect 39408 41206 39436 41686
rect 40132 41676 40184 41682
rect 40132 41618 40184 41624
rect 39672 41472 39724 41478
rect 39672 41414 39724 41420
rect 39304 41200 39356 41206
rect 39304 41142 39356 41148
rect 39396 41200 39448 41206
rect 39396 41142 39448 41148
rect 39488 40384 39540 40390
rect 39488 40326 39540 40332
rect 39304 39840 39356 39846
rect 39304 39782 39356 39788
rect 39396 39840 39448 39846
rect 39396 39782 39448 39788
rect 39316 39302 39344 39782
rect 39304 39296 39356 39302
rect 39304 39238 39356 39244
rect 39316 39098 39344 39238
rect 39304 39092 39356 39098
rect 39304 39034 39356 39040
rect 39212 38548 39264 38554
rect 39212 38490 39264 38496
rect 39028 38004 39080 38010
rect 39028 37946 39080 37952
rect 39028 37868 39080 37874
rect 39028 37810 39080 37816
rect 39040 37777 39068 37810
rect 39026 37768 39082 37777
rect 39026 37703 39082 37712
rect 39224 37670 39252 38490
rect 39408 38418 39436 39782
rect 39396 38412 39448 38418
rect 39396 38354 39448 38360
rect 39302 38176 39358 38185
rect 39302 38111 39358 38120
rect 39212 37664 39264 37670
rect 39212 37606 39264 37612
rect 39316 37330 39344 38111
rect 39408 37874 39436 38354
rect 39500 38010 39528 40326
rect 39488 38004 39540 38010
rect 39488 37946 39540 37952
rect 39396 37868 39448 37874
rect 39396 37810 39448 37816
rect 39408 37398 39436 37810
rect 39396 37392 39448 37398
rect 39396 37334 39448 37340
rect 39580 37392 39632 37398
rect 39580 37334 39632 37340
rect 39304 37324 39356 37330
rect 39304 37266 39356 37272
rect 39026 36952 39082 36961
rect 39120 36916 39172 36922
rect 39082 36896 39120 36904
rect 39026 36887 39120 36896
rect 39040 36876 39120 36887
rect 38936 36644 38988 36650
rect 38936 36586 38988 36592
rect 38948 36378 38976 36586
rect 38936 36372 38988 36378
rect 38936 36314 38988 36320
rect 39040 35766 39068 36876
rect 39120 36858 39172 36864
rect 39408 36786 39436 37334
rect 39396 36780 39448 36786
rect 39396 36722 39448 36728
rect 39488 36712 39540 36718
rect 39488 36654 39540 36660
rect 39396 36168 39448 36174
rect 39396 36110 39448 36116
rect 39212 36100 39264 36106
rect 39212 36042 39264 36048
rect 39304 36100 39356 36106
rect 39304 36042 39356 36048
rect 39028 35760 39080 35766
rect 39224 35737 39252 36042
rect 39028 35702 39080 35708
rect 39210 35728 39266 35737
rect 39210 35663 39266 35672
rect 39224 34921 39252 35663
rect 39316 35018 39344 36042
rect 39408 35034 39436 36110
rect 39500 35698 39528 36654
rect 39488 35692 39540 35698
rect 39488 35634 39540 35640
rect 39500 35601 39528 35634
rect 39486 35592 39542 35601
rect 39486 35527 39542 35536
rect 39500 35222 39528 35527
rect 39488 35216 39540 35222
rect 39488 35158 39540 35164
rect 39304 35012 39356 35018
rect 39408 35006 39528 35034
rect 39304 34954 39356 34960
rect 39210 34912 39266 34921
rect 39210 34847 39266 34856
rect 39028 34604 39080 34610
rect 39028 34546 39080 34552
rect 38844 34468 38896 34474
rect 38844 34410 38896 34416
rect 39040 34202 39068 34546
rect 39028 34196 39080 34202
rect 39028 34138 39080 34144
rect 39118 34096 39174 34105
rect 39118 34031 39174 34040
rect 39132 33998 39160 34031
rect 39120 33992 39172 33998
rect 39120 33934 39172 33940
rect 38936 33924 38988 33930
rect 38936 33866 38988 33872
rect 38948 33658 38976 33866
rect 39132 33844 39160 33934
rect 39396 33856 39448 33862
rect 39132 33816 39396 33844
rect 39396 33798 39448 33804
rect 38936 33652 38988 33658
rect 38936 33594 38988 33600
rect 39028 33652 39080 33658
rect 39028 33594 39080 33600
rect 38568 33584 38620 33590
rect 38568 33526 38620 33532
rect 39040 33318 39068 33594
rect 39394 33552 39450 33561
rect 39394 33487 39396 33496
rect 39448 33487 39450 33496
rect 39396 33458 39448 33464
rect 39500 33454 39528 35006
rect 39488 33448 39540 33454
rect 39488 33390 39540 33396
rect 38476 33312 38528 33318
rect 38476 33254 38528 33260
rect 38752 33312 38804 33318
rect 38752 33254 38804 33260
rect 39028 33312 39080 33318
rect 39028 33254 39080 33260
rect 38384 31272 38436 31278
rect 38384 31214 38436 31220
rect 38384 31136 38436 31142
rect 38384 31078 38436 31084
rect 38396 30054 38424 31078
rect 38488 30938 38516 33254
rect 38764 32609 38792 33254
rect 39396 32904 39448 32910
rect 39396 32846 39448 32852
rect 39304 32768 39356 32774
rect 39304 32710 39356 32716
rect 38750 32600 38806 32609
rect 38750 32535 38806 32544
rect 39316 32502 39344 32710
rect 39408 32502 39436 32846
rect 39304 32496 39356 32502
rect 39304 32438 39356 32444
rect 39396 32496 39448 32502
rect 39396 32438 39448 32444
rect 39120 32428 39172 32434
rect 39120 32370 39172 32376
rect 39028 32292 39080 32298
rect 39028 32234 39080 32240
rect 38750 31920 38806 31929
rect 38750 31855 38806 31864
rect 38764 31414 38792 31855
rect 38752 31408 38804 31414
rect 38752 31350 38804 31356
rect 39040 31226 39068 32234
rect 39132 31346 39160 32370
rect 39500 32298 39528 33390
rect 39396 32292 39448 32298
rect 39396 32234 39448 32240
rect 39488 32292 39540 32298
rect 39488 32234 39540 32240
rect 39408 32178 39436 32234
rect 39592 32178 39620 37334
rect 39684 36854 39712 41414
rect 39948 41268 40000 41274
rect 39948 41210 40000 41216
rect 39960 40458 39988 41210
rect 40144 40594 40172 41618
rect 40420 41562 40448 44200
rect 40500 42016 40552 42022
rect 40500 41958 40552 41964
rect 40592 42016 40644 42022
rect 40592 41958 40644 41964
rect 40328 41534 40448 41562
rect 40328 41478 40356 41534
rect 40316 41472 40368 41478
rect 40316 41414 40368 41420
rect 40408 41472 40460 41478
rect 40408 41414 40460 41420
rect 40420 40730 40448 41414
rect 40408 40724 40460 40730
rect 40408 40666 40460 40672
rect 40132 40588 40184 40594
rect 40132 40530 40184 40536
rect 39948 40452 40000 40458
rect 39948 40394 40000 40400
rect 40040 39568 40092 39574
rect 40040 39510 40092 39516
rect 40052 38758 40080 39510
rect 40408 39364 40460 39370
rect 40408 39306 40460 39312
rect 40316 39296 40368 39302
rect 40316 39238 40368 39244
rect 40132 39024 40184 39030
rect 40132 38966 40184 38972
rect 40222 38992 40278 39001
rect 40040 38752 40092 38758
rect 40040 38694 40092 38700
rect 40052 38350 40080 38694
rect 40144 38350 40172 38966
rect 40222 38927 40278 38936
rect 40040 38344 40092 38350
rect 40040 38286 40092 38292
rect 40132 38344 40184 38350
rect 40132 38286 40184 38292
rect 39856 38208 39908 38214
rect 39856 38150 39908 38156
rect 39868 37466 39896 38150
rect 40052 38010 40080 38286
rect 40040 38004 40092 38010
rect 40040 37946 40092 37952
rect 40040 37868 40092 37874
rect 40040 37810 40092 37816
rect 39856 37460 39908 37466
rect 39856 37402 39908 37408
rect 39672 36848 39724 36854
rect 39672 36790 39724 36796
rect 39868 36106 39896 37402
rect 40052 37369 40080 37810
rect 40038 37360 40094 37369
rect 40038 37295 40094 37304
rect 40236 37262 40264 38927
rect 40328 38826 40356 39238
rect 40420 39001 40448 39306
rect 40406 38992 40462 39001
rect 40406 38927 40462 38936
rect 40316 38820 40368 38826
rect 40316 38762 40368 38768
rect 40328 38026 40356 38762
rect 40512 38486 40540 41958
rect 40604 41546 40632 41958
rect 41984 41818 42012 44200
rect 42800 42152 42852 42158
rect 42800 42094 42852 42100
rect 41972 41812 42024 41818
rect 41972 41754 42024 41760
rect 42156 41608 42208 41614
rect 42156 41550 42208 41556
rect 40592 41540 40644 41546
rect 40592 41482 40644 41488
rect 41144 41472 41196 41478
rect 41144 41414 41196 41420
rect 41236 41472 41288 41478
rect 41236 41414 41288 41420
rect 41156 41138 41184 41414
rect 41144 41132 41196 41138
rect 41144 41074 41196 41080
rect 41248 39982 41276 41414
rect 41420 40996 41472 41002
rect 41420 40938 41472 40944
rect 41328 40928 41380 40934
rect 41328 40870 41380 40876
rect 41340 40526 41368 40870
rect 41432 40526 41460 40938
rect 41788 40928 41840 40934
rect 41788 40870 41840 40876
rect 41328 40520 41380 40526
rect 41328 40462 41380 40468
rect 41420 40520 41472 40526
rect 41420 40462 41472 40468
rect 41604 40384 41656 40390
rect 41604 40326 41656 40332
rect 41328 40180 41380 40186
rect 41328 40122 41380 40128
rect 41236 39976 41288 39982
rect 41236 39918 41288 39924
rect 41340 39642 41368 40122
rect 41328 39636 41380 39642
rect 41328 39578 41380 39584
rect 41144 39364 41196 39370
rect 41144 39306 41196 39312
rect 41156 39098 41184 39306
rect 41144 39092 41196 39098
rect 41144 39034 41196 39040
rect 40684 39024 40736 39030
rect 40684 38966 40736 38972
rect 40500 38480 40552 38486
rect 40500 38422 40552 38428
rect 40696 38282 40724 38966
rect 40868 38956 40920 38962
rect 40868 38898 40920 38904
rect 41052 38956 41104 38962
rect 41052 38898 41104 38904
rect 40880 38826 40908 38898
rect 40868 38820 40920 38826
rect 40868 38762 40920 38768
rect 40684 38276 40736 38282
rect 40684 38218 40736 38224
rect 40328 37998 40448 38026
rect 40316 37868 40368 37874
rect 40316 37810 40368 37816
rect 40224 37256 40276 37262
rect 40224 37198 40276 37204
rect 40328 37194 40356 37810
rect 40420 37806 40448 37998
rect 40592 37868 40644 37874
rect 40592 37810 40644 37816
rect 40408 37800 40460 37806
rect 40408 37742 40460 37748
rect 40604 37262 40632 37810
rect 40696 37466 40724 38218
rect 40776 37800 40828 37806
rect 40776 37742 40828 37748
rect 40684 37460 40736 37466
rect 40684 37402 40736 37408
rect 40788 37398 40816 37742
rect 40776 37392 40828 37398
rect 40682 37360 40738 37369
rect 40776 37334 40828 37340
rect 40682 37295 40738 37304
rect 40592 37256 40644 37262
rect 40592 37198 40644 37204
rect 40316 37188 40368 37194
rect 40316 37130 40368 37136
rect 40224 37120 40276 37126
rect 40224 37062 40276 37068
rect 39948 36848 40000 36854
rect 39948 36790 40000 36796
rect 39856 36100 39908 36106
rect 39856 36042 39908 36048
rect 39762 35728 39818 35737
rect 39762 35663 39764 35672
rect 39816 35663 39818 35672
rect 39764 35634 39816 35640
rect 39670 35048 39726 35057
rect 39670 34983 39672 34992
rect 39724 34983 39726 34992
rect 39672 34954 39724 34960
rect 39764 33992 39816 33998
rect 39764 33934 39816 33940
rect 39408 32150 39620 32178
rect 39212 32020 39264 32026
rect 39212 31962 39264 31968
rect 39120 31340 39172 31346
rect 39120 31282 39172 31288
rect 39040 31198 39160 31226
rect 38476 30932 38528 30938
rect 38476 30874 38528 30880
rect 38568 30592 38620 30598
rect 38568 30534 38620 30540
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 38474 30152 38530 30161
rect 38474 30087 38530 30096
rect 38384 30048 38436 30054
rect 38290 30016 38346 30025
rect 38384 29990 38436 29996
rect 38290 29951 38346 29960
rect 38200 29232 38252 29238
rect 38200 29174 38252 29180
rect 38108 29164 38160 29170
rect 38108 29106 38160 29112
rect 38016 28620 38068 28626
rect 38016 28562 38068 28568
rect 38016 28484 38068 28490
rect 38016 28426 38068 28432
rect 38028 28082 38056 28426
rect 38120 28150 38148 29106
rect 38212 28490 38240 29174
rect 38304 28694 38332 29951
rect 38292 28688 38344 28694
rect 38292 28630 38344 28636
rect 38200 28484 38252 28490
rect 38252 28444 38332 28472
rect 38200 28426 38252 28432
rect 38108 28144 38160 28150
rect 38108 28086 38160 28092
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 38120 27674 38148 28086
rect 38200 27872 38252 27878
rect 38200 27814 38252 27820
rect 38108 27668 38160 27674
rect 38108 27610 38160 27616
rect 38212 27577 38240 27814
rect 38198 27568 38254 27577
rect 38198 27503 38254 27512
rect 38016 27464 38068 27470
rect 37936 27424 38016 27452
rect 38016 27406 38068 27412
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 37830 27024 37886 27033
rect 37740 26988 37792 26994
rect 37830 26959 37886 26968
rect 37924 26988 37976 26994
rect 37740 26930 37792 26936
rect 37752 26858 37780 26930
rect 37740 26852 37792 26858
rect 37740 26794 37792 26800
rect 37844 25906 37872 26959
rect 37924 26930 37976 26936
rect 37936 26353 37964 26930
rect 37922 26344 37978 26353
rect 37922 26279 37978 26288
rect 37924 26240 37976 26246
rect 37924 26182 37976 26188
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37832 25764 37884 25770
rect 37832 25706 37884 25712
rect 37740 25696 37792 25702
rect 37740 25638 37792 25644
rect 37752 24818 37780 25638
rect 37844 25294 37872 25706
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37844 24954 37872 25230
rect 37832 24948 37884 24954
rect 37832 24890 37884 24896
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37752 24682 37780 24754
rect 37830 24712 37886 24721
rect 37740 24676 37792 24682
rect 37830 24647 37832 24656
rect 37740 24618 37792 24624
rect 37884 24647 37886 24656
rect 37832 24618 37884 24624
rect 37648 24200 37700 24206
rect 37648 24142 37700 24148
rect 37660 23526 37688 24142
rect 37752 23780 37780 24618
rect 37832 24132 37884 24138
rect 37832 24074 37884 24080
rect 37844 24041 37872 24074
rect 37830 24032 37886 24041
rect 37830 23967 37886 23976
rect 37832 23792 37884 23798
rect 37752 23752 37832 23780
rect 37832 23734 37884 23740
rect 37832 23656 37884 23662
rect 37830 23624 37832 23633
rect 37884 23624 37886 23633
rect 37830 23559 37886 23568
rect 37648 23520 37700 23526
rect 37648 23462 37700 23468
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37556 23112 37608 23118
rect 37556 23054 37608 23060
rect 37556 22976 37608 22982
rect 37556 22918 37608 22924
rect 37648 22976 37700 22982
rect 37648 22918 37700 22924
rect 37568 22642 37596 22918
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 37372 21480 37424 21486
rect 37372 21422 37424 21428
rect 37384 20330 37412 21422
rect 37464 21344 37516 21350
rect 37464 21286 37516 21292
rect 37476 21146 37504 21286
rect 37464 21140 37516 21146
rect 37464 21082 37516 21088
rect 37476 20602 37504 21082
rect 37556 20868 37608 20874
rect 37556 20810 37608 20816
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37372 20324 37424 20330
rect 37372 20266 37424 20272
rect 37464 20256 37516 20262
rect 37464 20198 37516 20204
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37096 19440 37148 19446
rect 37096 19382 37148 19388
rect 37200 19310 37228 19790
rect 37372 19780 37424 19786
rect 37372 19722 37424 19728
rect 37188 19304 37240 19310
rect 37188 19246 37240 19252
rect 37096 18760 37148 18766
rect 37096 18702 37148 18708
rect 37108 17270 37136 18702
rect 37200 18086 37228 19246
rect 37384 18902 37412 19722
rect 37372 18896 37424 18902
rect 37372 18838 37424 18844
rect 37384 18766 37412 18838
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 37476 18426 37504 20198
rect 37568 18970 37596 20810
rect 37660 20466 37688 22918
rect 37740 21956 37792 21962
rect 37740 21898 37792 21904
rect 37752 20874 37780 21898
rect 37844 21078 37872 23122
rect 37936 22778 37964 26182
rect 38028 24682 38056 27406
rect 38120 26897 38148 27406
rect 38106 26888 38162 26897
rect 38106 26823 38162 26832
rect 38108 26784 38160 26790
rect 38108 26726 38160 26732
rect 38120 26042 38148 26726
rect 38108 26036 38160 26042
rect 38108 25978 38160 25984
rect 38016 24676 38068 24682
rect 38016 24618 38068 24624
rect 38014 24304 38070 24313
rect 38014 24239 38070 24248
rect 38028 24206 38056 24239
rect 38016 24200 38068 24206
rect 38016 24142 38068 24148
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38028 23361 38056 24006
rect 38014 23352 38070 23361
rect 38014 23287 38070 23296
rect 37924 22772 37976 22778
rect 37924 22714 37976 22720
rect 37924 22636 37976 22642
rect 37924 22578 37976 22584
rect 37832 21072 37884 21078
rect 37832 21014 37884 21020
rect 37936 20942 37964 22578
rect 38120 22522 38148 25978
rect 38212 22642 38240 27503
rect 38304 27033 38332 28444
rect 38396 27538 38424 29990
rect 38488 29238 38516 30087
rect 38580 29782 38608 30534
rect 38752 30184 38804 30190
rect 38752 30126 38804 30132
rect 38568 29776 38620 29782
rect 38568 29718 38620 29724
rect 38568 29640 38620 29646
rect 38568 29582 38620 29588
rect 38476 29232 38528 29238
rect 38476 29174 38528 29180
rect 38488 29034 38516 29174
rect 38580 29170 38608 29582
rect 38568 29164 38620 29170
rect 38568 29106 38620 29112
rect 38476 29028 38528 29034
rect 38476 28970 38528 28976
rect 38476 28552 38528 28558
rect 38476 28494 38528 28500
rect 38384 27532 38436 27538
rect 38384 27474 38436 27480
rect 38396 27062 38424 27474
rect 38488 27334 38516 28494
rect 38580 28490 38608 29106
rect 38764 28762 38792 30126
rect 38752 28756 38804 28762
rect 38752 28698 38804 28704
rect 38568 28484 38620 28490
rect 38568 28426 38620 28432
rect 38580 27946 38608 28426
rect 38568 27940 38620 27946
rect 38568 27882 38620 27888
rect 38660 27872 38712 27878
rect 38856 27826 38884 30534
rect 39028 30048 39080 30054
rect 39028 29990 39080 29996
rect 39040 29578 39068 29990
rect 39028 29572 39080 29578
rect 39028 29514 39080 29520
rect 39040 29186 39068 29514
rect 38948 29158 39068 29186
rect 38948 29102 38976 29158
rect 38936 29096 38988 29102
rect 39028 29096 39080 29102
rect 38936 29038 38988 29044
rect 39026 29064 39028 29073
rect 39080 29064 39082 29073
rect 38660 27814 38712 27820
rect 38672 27554 38700 27814
rect 38580 27526 38700 27554
rect 38764 27798 38884 27826
rect 38580 27470 38608 27526
rect 38568 27464 38620 27470
rect 38568 27406 38620 27412
rect 38476 27328 38528 27334
rect 38474 27296 38476 27305
rect 38528 27296 38530 27305
rect 38474 27231 38530 27240
rect 38384 27056 38436 27062
rect 38290 27024 38346 27033
rect 38384 26998 38436 27004
rect 38290 26959 38292 26968
rect 38344 26959 38346 26968
rect 38292 26930 38344 26936
rect 38476 26920 38528 26926
rect 38382 26888 38438 26897
rect 38476 26862 38528 26868
rect 38382 26823 38438 26832
rect 38396 26518 38424 26823
rect 38384 26512 38436 26518
rect 38384 26454 38436 26460
rect 38384 26376 38436 26382
rect 38384 26318 38436 26324
rect 38292 25900 38344 25906
rect 38292 25842 38344 25848
rect 38304 25226 38332 25842
rect 38396 25294 38424 26318
rect 38488 26217 38516 26862
rect 38580 26382 38608 27406
rect 38764 26926 38792 27798
rect 38844 27668 38896 27674
rect 38844 27610 38896 27616
rect 38752 26920 38804 26926
rect 38752 26862 38804 26868
rect 38856 26790 38884 27610
rect 38948 27554 38976 29038
rect 39026 28999 39082 29008
rect 39132 28490 39160 31198
rect 39224 31142 39252 31962
rect 39396 31680 39448 31686
rect 39396 31622 39448 31628
rect 39408 31346 39436 31622
rect 39396 31340 39448 31346
rect 39448 31300 39528 31328
rect 39396 31282 39448 31288
rect 39212 31136 39264 31142
rect 39212 31078 39264 31084
rect 39396 30728 39448 30734
rect 39394 30696 39396 30705
rect 39448 30696 39450 30705
rect 39394 30631 39450 30640
rect 39212 29844 39264 29850
rect 39212 29786 39264 29792
rect 39224 29073 39252 29786
rect 39304 29504 39356 29510
rect 39304 29446 39356 29452
rect 39210 29064 39266 29073
rect 39210 28999 39266 29008
rect 39120 28484 39172 28490
rect 39120 28426 39172 28432
rect 39212 27872 39264 27878
rect 39212 27814 39264 27820
rect 38948 27526 39160 27554
rect 39026 27432 39082 27441
rect 39026 27367 39028 27376
rect 39080 27367 39082 27376
rect 39028 27338 39080 27344
rect 39132 26858 39160 27526
rect 39224 26926 39252 27814
rect 39212 26920 39264 26926
rect 39212 26862 39264 26868
rect 39120 26852 39172 26858
rect 39120 26794 39172 26800
rect 38844 26784 38896 26790
rect 38844 26726 38896 26732
rect 39132 26450 39160 26794
rect 39120 26444 39172 26450
rect 39120 26386 39172 26392
rect 38568 26376 38620 26382
rect 38568 26318 38620 26324
rect 38752 26240 38804 26246
rect 38474 26208 38530 26217
rect 38752 26182 38804 26188
rect 38474 26143 38530 26152
rect 38384 25288 38436 25294
rect 38384 25230 38436 25236
rect 38292 25220 38344 25226
rect 38292 25162 38344 25168
rect 38384 24200 38436 24206
rect 38384 24142 38436 24148
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38304 23050 38332 23666
rect 38396 23526 38424 24142
rect 38476 24064 38528 24070
rect 38476 24006 38528 24012
rect 38568 24064 38620 24070
rect 38568 24006 38620 24012
rect 38384 23520 38436 23526
rect 38384 23462 38436 23468
rect 38488 23322 38516 24006
rect 38476 23316 38528 23322
rect 38476 23258 38528 23264
rect 38580 23118 38608 24006
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38568 23112 38620 23118
rect 38568 23054 38620 23060
rect 38292 23044 38344 23050
rect 38292 22986 38344 22992
rect 38200 22636 38252 22642
rect 38200 22578 38252 22584
rect 38120 22494 38240 22522
rect 38212 22098 38240 22494
rect 38200 22092 38252 22098
rect 38200 22034 38252 22040
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37740 20868 37792 20874
rect 37740 20810 37792 20816
rect 37648 20460 37700 20466
rect 37648 20402 37700 20408
rect 37648 20256 37700 20262
rect 37648 20198 37700 20204
rect 37660 19990 37688 20198
rect 37648 19984 37700 19990
rect 37648 19926 37700 19932
rect 37832 19984 37884 19990
rect 37832 19926 37884 19932
rect 37740 19848 37792 19854
rect 37740 19790 37792 19796
rect 37752 19496 37780 19790
rect 37660 19468 37780 19496
rect 37660 19174 37688 19468
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 37648 19168 37700 19174
rect 37648 19110 37700 19116
rect 37556 18964 37608 18970
rect 37556 18906 37608 18912
rect 37556 18760 37608 18766
rect 37556 18702 37608 18708
rect 37464 18420 37516 18426
rect 37464 18362 37516 18368
rect 37568 18306 37596 18702
rect 37476 18278 37596 18306
rect 37188 18080 37240 18086
rect 37188 18022 37240 18028
rect 37096 17264 37148 17270
rect 37096 17206 37148 17212
rect 37108 16153 37136 17206
rect 37200 16726 37228 18022
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37188 16720 37240 16726
rect 37188 16662 37240 16668
rect 37200 16590 37228 16662
rect 37384 16658 37412 17138
rect 37476 17066 37504 18278
rect 37556 18216 37608 18222
rect 37556 18158 37608 18164
rect 37568 18086 37596 18158
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 37464 17060 37516 17066
rect 37464 17002 37516 17008
rect 37568 16998 37596 18022
rect 37660 17882 37688 19110
rect 37752 18698 37780 19314
rect 37740 18692 37792 18698
rect 37740 18634 37792 18640
rect 37752 18290 37780 18634
rect 37740 18284 37792 18290
rect 37740 18226 37792 18232
rect 37648 17876 37700 17882
rect 37648 17818 37700 17824
rect 37752 17678 37780 18226
rect 37844 17746 37872 19926
rect 37936 18970 37964 20878
rect 38028 20806 38056 21966
rect 38108 21888 38160 21894
rect 38108 21830 38160 21836
rect 38120 21554 38148 21830
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 38028 20466 38056 20742
rect 38016 20460 38068 20466
rect 38016 20402 38068 20408
rect 38016 20256 38068 20262
rect 38016 20198 38068 20204
rect 38028 19922 38056 20198
rect 38016 19916 38068 19922
rect 38016 19858 38068 19864
rect 38304 19514 38332 22986
rect 38384 22772 38436 22778
rect 38384 22714 38436 22720
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38396 19428 38424 22714
rect 38568 22024 38620 22030
rect 38568 21966 38620 21972
rect 38476 21480 38528 21486
rect 38476 21422 38528 21428
rect 38488 21010 38516 21422
rect 38476 21004 38528 21010
rect 38476 20946 38528 20952
rect 38580 20058 38608 21966
rect 38568 20052 38620 20058
rect 38568 19994 38620 20000
rect 38580 19786 38608 19994
rect 38672 19854 38700 23258
rect 38764 23186 38792 26182
rect 39224 26042 39252 26862
rect 39212 26036 39264 26042
rect 39212 25978 39264 25984
rect 39210 25936 39266 25945
rect 39120 25900 39172 25906
rect 39210 25871 39212 25880
rect 39120 25842 39172 25848
rect 39264 25871 39266 25880
rect 39212 25842 39264 25848
rect 39132 25498 39160 25842
rect 39120 25492 39172 25498
rect 39120 25434 39172 25440
rect 39132 25276 39160 25434
rect 39224 25430 39252 25842
rect 39212 25424 39264 25430
rect 39212 25366 39264 25372
rect 39316 25294 39344 29446
rect 39408 29050 39436 30631
rect 39500 29170 39528 31300
rect 39580 31272 39632 31278
rect 39580 31214 39632 31220
rect 39592 30258 39620 31214
rect 39580 30252 39632 30258
rect 39580 30194 39632 30200
rect 39592 30122 39620 30194
rect 39580 30116 39632 30122
rect 39580 30058 39632 30064
rect 39592 29850 39620 30058
rect 39672 30048 39724 30054
rect 39672 29990 39724 29996
rect 39580 29844 39632 29850
rect 39580 29786 39632 29792
rect 39580 29504 39632 29510
rect 39580 29446 39632 29452
rect 39592 29238 39620 29446
rect 39580 29232 39632 29238
rect 39580 29174 39632 29180
rect 39684 29170 39712 29990
rect 39488 29164 39540 29170
rect 39488 29106 39540 29112
rect 39672 29164 39724 29170
rect 39672 29106 39724 29112
rect 39580 29096 39632 29102
rect 39408 29044 39580 29050
rect 39408 29038 39632 29044
rect 39408 29022 39620 29038
rect 39672 28484 39724 28490
rect 39672 28426 39724 28432
rect 39396 27872 39448 27878
rect 39396 27814 39448 27820
rect 39408 27062 39436 27814
rect 39488 27464 39540 27470
rect 39488 27406 39540 27412
rect 39396 27056 39448 27062
rect 39396 26998 39448 27004
rect 39408 26450 39436 26998
rect 39396 26444 39448 26450
rect 39396 26386 39448 26392
rect 39396 26036 39448 26042
rect 39396 25978 39448 25984
rect 39212 25288 39264 25294
rect 39132 25248 39212 25276
rect 39212 25230 39264 25236
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 39120 25152 39172 25158
rect 39120 25094 39172 25100
rect 39028 24608 39080 24614
rect 39028 24550 39080 24556
rect 39040 23798 39068 24550
rect 39028 23792 39080 23798
rect 38934 23760 38990 23769
rect 39028 23734 39080 23740
rect 38934 23695 38990 23704
rect 38752 23180 38804 23186
rect 38752 23122 38804 23128
rect 38844 23180 38896 23186
rect 38844 23122 38896 23128
rect 38856 22506 38884 23122
rect 38948 22930 38976 23695
rect 38948 22902 39068 22930
rect 38936 22772 38988 22778
rect 38936 22714 38988 22720
rect 38844 22500 38896 22506
rect 38844 22442 38896 22448
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 38856 21690 38884 21966
rect 38844 21684 38896 21690
rect 38844 21626 38896 21632
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38764 20942 38792 21490
rect 38752 20936 38804 20942
rect 38752 20878 38804 20884
rect 38660 19848 38712 19854
rect 38660 19790 38712 19796
rect 38568 19780 38620 19786
rect 38568 19722 38620 19728
rect 38568 19440 38620 19446
rect 38396 19400 38568 19428
rect 38568 19382 38620 19388
rect 37924 18964 37976 18970
rect 37924 18906 37976 18912
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 37936 18358 37964 18702
rect 38660 18692 38712 18698
rect 38660 18634 38712 18640
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 37924 18352 37976 18358
rect 37924 18294 37976 18300
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 37832 17740 37884 17746
rect 37832 17682 37884 17688
rect 37648 17672 37700 17678
rect 37648 17614 37700 17620
rect 37740 17672 37792 17678
rect 37740 17614 37792 17620
rect 37660 17338 37688 17614
rect 37752 17542 37780 17614
rect 37740 17536 37792 17542
rect 37740 17478 37792 17484
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 37556 16992 37608 16998
rect 37556 16934 37608 16940
rect 37844 16794 37872 17682
rect 37936 17678 37964 17818
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37924 17536 37976 17542
rect 37924 17478 37976 17484
rect 37740 16788 37792 16794
rect 37740 16730 37792 16736
rect 37832 16788 37884 16794
rect 37832 16730 37884 16736
rect 37372 16652 37424 16658
rect 37372 16594 37424 16600
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37200 16250 37228 16526
rect 37188 16244 37240 16250
rect 37188 16186 37240 16192
rect 37094 16144 37150 16153
rect 37094 16079 37150 16088
rect 37108 15162 37136 16079
rect 37200 15910 37228 16186
rect 37292 15978 37320 16526
rect 37280 15972 37332 15978
rect 37280 15914 37332 15920
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37096 15156 37148 15162
rect 37096 15098 37148 15104
rect 37200 14414 37228 15506
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 37096 14068 37148 14074
rect 37096 14010 37148 14016
rect 37108 12442 37136 14010
rect 37292 13258 37320 14894
rect 37384 14074 37412 16594
rect 37648 16516 37700 16522
rect 37648 16458 37700 16464
rect 37660 15026 37688 16458
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37384 13410 37412 14010
rect 37476 13938 37504 14962
rect 37752 14414 37780 16730
rect 37936 16674 37964 17478
rect 37844 16646 37964 16674
rect 37844 14822 37872 16646
rect 38028 16522 38056 18362
rect 38476 17604 38528 17610
rect 38476 17546 38528 17552
rect 38384 17196 38436 17202
rect 38384 17138 38436 17144
rect 38292 16992 38344 16998
rect 38292 16934 38344 16940
rect 38108 16584 38160 16590
rect 38108 16526 38160 16532
rect 38016 16516 38068 16522
rect 38016 16458 38068 16464
rect 37924 16448 37976 16454
rect 37924 16390 37976 16396
rect 37936 15978 37964 16390
rect 37924 15972 37976 15978
rect 37924 15914 37976 15920
rect 37936 15502 37964 15914
rect 37924 15496 37976 15502
rect 37924 15438 37976 15444
rect 38120 15094 38148 16526
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38212 15706 38240 16050
rect 38200 15700 38252 15706
rect 38200 15642 38252 15648
rect 37924 15088 37976 15094
rect 37924 15030 37976 15036
rect 38108 15088 38160 15094
rect 38108 15030 38160 15036
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37740 14408 37792 14414
rect 37740 14350 37792 14356
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37476 13530 37504 13874
rect 37464 13524 37516 13530
rect 37464 13466 37516 13472
rect 37384 13382 37504 13410
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 36924 12406 37044 12434
rect 37096 12436 37148 12442
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 34796 11756 34848 11762
rect 34716 11716 34796 11744
rect 34060 11698 34112 11704
rect 34796 11698 34848 11704
rect 34980 11756 35032 11762
rect 34980 11698 35032 11704
rect 36176 11756 36228 11762
rect 36176 11698 36228 11704
rect 34992 11626 35020 11698
rect 34980 11620 35032 11626
rect 34980 11562 35032 11568
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 34152 11144 34204 11150
rect 34152 11086 34204 11092
rect 33140 11076 33192 11082
rect 33140 11018 33192 11024
rect 33692 11076 33744 11082
rect 33692 11018 33744 11024
rect 33152 10810 33180 11018
rect 34164 10810 34192 11086
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 34152 10804 34204 10810
rect 34152 10746 34204 10752
rect 32864 10600 32916 10606
rect 32864 10542 32916 10548
rect 34440 10538 34468 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35452 10810 35480 11494
rect 36924 11286 36952 12406
rect 37096 12378 37148 12384
rect 37292 12170 37320 13194
rect 37280 12164 37332 12170
rect 37280 12106 37332 12112
rect 37292 11830 37320 12106
rect 37384 11898 37412 13262
rect 37476 12850 37504 13382
rect 37568 13326 37596 14350
rect 37752 13870 37780 14350
rect 37936 14278 37964 15030
rect 38120 14618 38148 15030
rect 38108 14612 38160 14618
rect 38108 14554 38160 14560
rect 38120 14482 38148 14554
rect 38198 14512 38254 14521
rect 38108 14476 38160 14482
rect 38198 14447 38200 14456
rect 38108 14418 38160 14424
rect 38252 14447 38254 14456
rect 38200 14418 38252 14424
rect 38304 14346 38332 16934
rect 38396 16794 38424 17138
rect 38488 16998 38516 17546
rect 38476 16992 38528 16998
rect 38528 16952 38608 16980
rect 38476 16934 38528 16940
rect 38384 16788 38436 16794
rect 38384 16730 38436 16736
rect 38396 16114 38424 16730
rect 38476 16652 38528 16658
rect 38476 16594 38528 16600
rect 38488 16114 38516 16594
rect 38384 16108 38436 16114
rect 38384 16050 38436 16056
rect 38476 16108 38528 16114
rect 38476 16050 38528 16056
rect 38396 15570 38424 16050
rect 38384 15564 38436 15570
rect 38384 15506 38436 15512
rect 38396 15162 38424 15506
rect 38384 15156 38436 15162
rect 38384 15098 38436 15104
rect 38292 14340 38344 14346
rect 38292 14282 38344 14288
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 38304 14074 38332 14282
rect 38580 14278 38608 16952
rect 38672 16250 38700 18634
rect 38764 18086 38792 20878
rect 38948 20398 38976 22714
rect 39040 22438 39068 22902
rect 39028 22432 39080 22438
rect 39028 22374 39080 22380
rect 39028 22228 39080 22234
rect 39028 22170 39080 22176
rect 39040 21010 39068 22170
rect 39132 22098 39160 25094
rect 39408 24206 39436 25978
rect 39500 25974 39528 27406
rect 39580 26852 39632 26858
rect 39684 26840 39712 28426
rect 39776 26908 39804 33934
rect 39960 33522 39988 36790
rect 40236 36786 40264 37062
rect 40328 36786 40356 37130
rect 40604 36786 40632 37198
rect 40132 36780 40184 36786
rect 40132 36722 40184 36728
rect 40224 36780 40276 36786
rect 40224 36722 40276 36728
rect 40316 36780 40368 36786
rect 40316 36722 40368 36728
rect 40592 36780 40644 36786
rect 40592 36722 40644 36728
rect 40144 36310 40172 36722
rect 40132 36304 40184 36310
rect 40132 36246 40184 36252
rect 40222 36272 40278 36281
rect 40222 36207 40278 36216
rect 40236 36174 40264 36207
rect 40224 36168 40276 36174
rect 40224 36110 40276 36116
rect 40328 36106 40356 36722
rect 40500 36168 40552 36174
rect 40420 36128 40500 36156
rect 40316 36100 40368 36106
rect 40316 36042 40368 36048
rect 40328 35834 40356 36042
rect 40316 35828 40368 35834
rect 40316 35770 40368 35776
rect 40328 35630 40356 35770
rect 40420 35698 40448 36128
rect 40604 36156 40632 36722
rect 40552 36128 40632 36156
rect 40500 36110 40552 36116
rect 40408 35692 40460 35698
rect 40408 35634 40460 35640
rect 40500 35692 40552 35698
rect 40500 35634 40552 35640
rect 40592 35692 40644 35698
rect 40696 35680 40724 37295
rect 40776 37188 40828 37194
rect 40776 37130 40828 37136
rect 40788 36922 40816 37130
rect 40776 36916 40828 36922
rect 40776 36858 40828 36864
rect 40880 35986 40908 38762
rect 41064 38554 41092 38898
rect 41144 38888 41196 38894
rect 41144 38830 41196 38836
rect 41052 38548 41104 38554
rect 41052 38490 41104 38496
rect 41052 38412 41104 38418
rect 41052 38354 41104 38360
rect 40960 37936 41012 37942
rect 40960 37878 41012 37884
rect 40644 35652 40724 35680
rect 40788 35958 40908 35986
rect 40592 35634 40644 35640
rect 40316 35624 40368 35630
rect 40316 35566 40368 35572
rect 40420 35562 40448 35634
rect 40408 35556 40460 35562
rect 40408 35498 40460 35504
rect 40420 35154 40448 35498
rect 40512 35290 40540 35634
rect 40592 35488 40644 35494
rect 40592 35430 40644 35436
rect 40500 35284 40552 35290
rect 40500 35226 40552 35232
rect 40604 35154 40632 35430
rect 40408 35148 40460 35154
rect 40408 35090 40460 35096
rect 40592 35148 40644 35154
rect 40592 35090 40644 35096
rect 40132 35080 40184 35086
rect 40132 35022 40184 35028
rect 40144 34542 40172 35022
rect 40316 34672 40368 34678
rect 40314 34640 40316 34649
rect 40368 34640 40370 34649
rect 40224 34604 40276 34610
rect 40314 34575 40370 34584
rect 40224 34546 40276 34552
rect 40132 34536 40184 34542
rect 40132 34478 40184 34484
rect 40040 33992 40092 33998
rect 40038 33960 40040 33969
rect 40092 33960 40094 33969
rect 40038 33895 40094 33904
rect 39948 33516 40000 33522
rect 39948 33458 40000 33464
rect 40236 33153 40264 34546
rect 40222 33144 40278 33153
rect 40222 33079 40278 33088
rect 40040 32904 40092 32910
rect 40040 32846 40092 32852
rect 39948 32836 40000 32842
rect 39948 32778 40000 32784
rect 39856 32564 39908 32570
rect 39856 32506 39908 32512
rect 39868 32026 39896 32506
rect 39856 32020 39908 32026
rect 39856 31962 39908 31968
rect 39868 30734 39896 31962
rect 39960 31754 39988 32778
rect 40052 32366 40080 32846
rect 40040 32360 40092 32366
rect 40040 32302 40092 32308
rect 39948 31748 40000 31754
rect 39948 31690 40000 31696
rect 39856 30728 39908 30734
rect 39856 30670 39908 30676
rect 39868 28014 39896 30670
rect 39960 29646 39988 31690
rect 40052 31414 40080 32302
rect 40316 31952 40368 31958
rect 40316 31894 40368 31900
rect 40132 31884 40184 31890
rect 40132 31826 40184 31832
rect 40040 31408 40092 31414
rect 40040 31350 40092 31356
rect 40144 31210 40172 31826
rect 40224 31816 40276 31822
rect 40328 31793 40356 31894
rect 40224 31758 40276 31764
rect 40314 31784 40370 31793
rect 40040 31204 40092 31210
rect 40040 31146 40092 31152
rect 40132 31204 40184 31210
rect 40132 31146 40184 31152
rect 40052 30394 40080 31146
rect 40236 31142 40264 31758
rect 40314 31719 40370 31728
rect 40420 31686 40448 35090
rect 40500 34944 40552 34950
rect 40500 34886 40552 34892
rect 40512 34678 40540 34886
rect 40500 34672 40552 34678
rect 40500 34614 40552 34620
rect 40788 33522 40816 35958
rect 40866 35864 40922 35873
rect 40866 35799 40922 35808
rect 40880 35698 40908 35799
rect 40868 35692 40920 35698
rect 40868 35634 40920 35640
rect 40880 35601 40908 35634
rect 40866 35592 40922 35601
rect 40866 35527 40922 35536
rect 40972 35018 41000 37878
rect 41064 37652 41092 38354
rect 41156 38350 41184 38830
rect 41144 38344 41196 38350
rect 41144 38286 41196 38292
rect 41156 37942 41184 38286
rect 41144 37936 41196 37942
rect 41328 37936 41380 37942
rect 41196 37896 41276 37924
rect 41144 37878 41196 37884
rect 41144 37664 41196 37670
rect 41064 37624 41144 37652
rect 41144 37606 41196 37612
rect 41156 37262 41184 37606
rect 41248 37262 41276 37896
rect 41328 37878 41380 37884
rect 41144 37256 41196 37262
rect 41144 37198 41196 37204
rect 41236 37256 41288 37262
rect 41236 37198 41288 37204
rect 41052 36712 41104 36718
rect 41052 36654 41104 36660
rect 41064 36038 41092 36654
rect 41156 36378 41184 37198
rect 41340 37194 41368 37878
rect 41512 37664 41564 37670
rect 41512 37606 41564 37612
rect 41420 37392 41472 37398
rect 41420 37334 41472 37340
rect 41328 37188 41380 37194
rect 41328 37130 41380 37136
rect 41432 36922 41460 37334
rect 41420 36916 41472 36922
rect 41420 36858 41472 36864
rect 41524 36786 41552 37606
rect 41236 36780 41288 36786
rect 41512 36780 41564 36786
rect 41236 36722 41288 36728
rect 41432 36740 41512 36768
rect 41144 36372 41196 36378
rect 41144 36314 41196 36320
rect 41248 36174 41276 36722
rect 41328 36576 41380 36582
rect 41328 36518 41380 36524
rect 41236 36168 41288 36174
rect 41236 36110 41288 36116
rect 41052 36032 41104 36038
rect 41052 35974 41104 35980
rect 41248 35834 41276 36110
rect 41236 35828 41288 35834
rect 41236 35770 41288 35776
rect 41340 35630 41368 36518
rect 41432 36174 41460 36740
rect 41512 36722 41564 36728
rect 41420 36168 41472 36174
rect 41420 36110 41472 36116
rect 41512 36168 41564 36174
rect 41512 36110 41564 36116
rect 41328 35624 41380 35630
rect 41328 35566 41380 35572
rect 41340 35086 41368 35566
rect 41524 35154 41552 36110
rect 41512 35148 41564 35154
rect 41512 35090 41564 35096
rect 41328 35080 41380 35086
rect 41328 35022 41380 35028
rect 40960 35012 41012 35018
rect 40960 34954 41012 34960
rect 40960 34400 41012 34406
rect 40960 34342 41012 34348
rect 40972 34202 41000 34342
rect 40960 34196 41012 34202
rect 40960 34138 41012 34144
rect 41052 34196 41104 34202
rect 41052 34138 41104 34144
rect 41064 33590 41092 34138
rect 41420 34128 41472 34134
rect 41420 34070 41472 34076
rect 41328 33992 41380 33998
rect 41328 33934 41380 33940
rect 41052 33584 41104 33590
rect 41052 33526 41104 33532
rect 40776 33516 40828 33522
rect 40776 33458 40828 33464
rect 40868 33516 40920 33522
rect 40868 33458 40920 33464
rect 40880 33289 40908 33458
rect 40866 33280 40922 33289
rect 40866 33215 40922 33224
rect 40960 33040 41012 33046
rect 40960 32982 41012 32988
rect 40776 32904 40828 32910
rect 40776 32846 40828 32852
rect 40868 32904 40920 32910
rect 40868 32846 40920 32852
rect 40500 32768 40552 32774
rect 40500 32710 40552 32716
rect 40684 32768 40736 32774
rect 40684 32710 40736 32716
rect 40512 32366 40540 32710
rect 40592 32428 40644 32434
rect 40592 32370 40644 32376
rect 40500 32360 40552 32366
rect 40500 32302 40552 32308
rect 40604 32026 40632 32370
rect 40592 32020 40644 32026
rect 40592 31962 40644 31968
rect 40498 31920 40554 31929
rect 40498 31855 40554 31864
rect 40408 31680 40460 31686
rect 40408 31622 40460 31628
rect 40512 31464 40540 31855
rect 40696 31822 40724 32710
rect 40788 32434 40816 32846
rect 40776 32428 40828 32434
rect 40776 32370 40828 32376
rect 40684 31816 40736 31822
rect 40590 31784 40646 31793
rect 40684 31758 40736 31764
rect 40590 31719 40646 31728
rect 40420 31436 40540 31464
rect 40316 31408 40368 31414
rect 40316 31350 40368 31356
rect 40224 31136 40276 31142
rect 40224 31078 40276 31084
rect 40328 30954 40356 31350
rect 40132 30932 40184 30938
rect 40132 30874 40184 30880
rect 40236 30926 40356 30954
rect 40040 30388 40092 30394
rect 40040 30330 40092 30336
rect 40144 30258 40172 30874
rect 40236 30734 40264 30926
rect 40224 30728 40276 30734
rect 40224 30670 40276 30676
rect 40132 30252 40184 30258
rect 40132 30194 40184 30200
rect 39948 29640 40000 29646
rect 39948 29582 40000 29588
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 40052 28082 40080 28494
rect 40040 28076 40092 28082
rect 40040 28018 40092 28024
rect 39856 28008 39908 28014
rect 39856 27950 39908 27956
rect 39868 27062 39896 27950
rect 39948 27940 40000 27946
rect 39948 27882 40000 27888
rect 39960 27606 39988 27882
rect 39948 27600 40000 27606
rect 39948 27542 40000 27548
rect 39856 27056 39908 27062
rect 39856 26998 39908 27004
rect 39776 26880 39896 26908
rect 39684 26812 39804 26840
rect 39580 26794 39632 26800
rect 39488 25968 39540 25974
rect 39488 25910 39540 25916
rect 39488 25696 39540 25702
rect 39592 25684 39620 26794
rect 39672 26376 39724 26382
rect 39672 26318 39724 26324
rect 39540 25656 39620 25684
rect 39488 25638 39540 25644
rect 39500 24750 39528 25638
rect 39580 25220 39632 25226
rect 39580 25162 39632 25168
rect 39488 24744 39540 24750
rect 39488 24686 39540 24692
rect 39488 24608 39540 24614
rect 39488 24550 39540 24556
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39212 23792 39264 23798
rect 39408 23769 39436 24142
rect 39212 23734 39264 23740
rect 39394 23760 39450 23769
rect 39224 23322 39252 23734
rect 39500 23730 39528 24550
rect 39394 23695 39450 23704
rect 39488 23724 39540 23730
rect 39488 23666 39540 23672
rect 39212 23316 39264 23322
rect 39212 23258 39264 23264
rect 39500 23202 39528 23666
rect 39316 23186 39528 23202
rect 39304 23180 39528 23186
rect 39356 23174 39528 23180
rect 39304 23122 39356 23128
rect 39212 23112 39264 23118
rect 39212 23054 39264 23060
rect 39488 23112 39540 23118
rect 39488 23054 39540 23060
rect 39224 22642 39252 23054
rect 39304 22976 39356 22982
rect 39304 22918 39356 22924
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 39316 22506 39344 22918
rect 39500 22778 39528 23054
rect 39488 22772 39540 22778
rect 39488 22714 39540 22720
rect 39396 22636 39448 22642
rect 39396 22578 39448 22584
rect 39304 22500 39356 22506
rect 39304 22442 39356 22448
rect 39304 22228 39356 22234
rect 39304 22170 39356 22176
rect 39120 22092 39172 22098
rect 39172 22052 39252 22080
rect 39120 22034 39172 22040
rect 39120 21956 39172 21962
rect 39120 21898 39172 21904
rect 39028 21004 39080 21010
rect 39028 20946 39080 20952
rect 39028 20800 39080 20806
rect 39028 20742 39080 20748
rect 38936 20392 38988 20398
rect 38936 20334 38988 20340
rect 39040 19854 39068 20742
rect 39132 20330 39160 21898
rect 39224 21350 39252 22052
rect 39316 21894 39344 22170
rect 39304 21888 39356 21894
rect 39304 21830 39356 21836
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 39212 20936 39264 20942
rect 39212 20878 39264 20884
rect 39224 20466 39252 20878
rect 39212 20460 39264 20466
rect 39212 20402 39264 20408
rect 39120 20324 39172 20330
rect 39120 20266 39172 20272
rect 39028 19848 39080 19854
rect 39028 19790 39080 19796
rect 39304 19712 39356 19718
rect 39304 19654 39356 19660
rect 39120 19508 39172 19514
rect 39316 19496 39344 19654
rect 39172 19468 39344 19496
rect 39120 19450 39172 19456
rect 39316 19378 39344 19468
rect 39028 19372 39080 19378
rect 39028 19314 39080 19320
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 39304 19372 39356 19378
rect 39304 19314 39356 19320
rect 38936 19304 38988 19310
rect 38936 19246 38988 19252
rect 38844 18896 38896 18902
rect 38844 18838 38896 18844
rect 38856 18290 38884 18838
rect 38948 18630 38976 19246
rect 39040 18630 39068 19314
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 39028 18624 39080 18630
rect 39028 18566 39080 18572
rect 39120 18624 39172 18630
rect 39120 18566 39172 18572
rect 39040 18426 39068 18566
rect 39028 18420 39080 18426
rect 39028 18362 39080 18368
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38856 17762 38884 18226
rect 39028 17876 39080 17882
rect 39028 17818 39080 17824
rect 38856 17734 38976 17762
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38752 17536 38804 17542
rect 38752 17478 38804 17484
rect 38764 17270 38792 17478
rect 38752 17264 38804 17270
rect 38752 17206 38804 17212
rect 38764 16590 38792 17206
rect 38856 17134 38884 17614
rect 38948 17202 38976 17734
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38844 17128 38896 17134
rect 39040 17082 39068 17818
rect 39132 17814 39160 18566
rect 39224 18426 39252 19314
rect 39302 19000 39358 19009
rect 39302 18935 39304 18944
rect 39356 18935 39358 18944
rect 39304 18906 39356 18912
rect 39212 18420 39264 18426
rect 39212 18362 39264 18368
rect 39212 18284 39264 18290
rect 39212 18226 39264 18232
rect 39120 17808 39172 17814
rect 39120 17750 39172 17756
rect 38844 17070 38896 17076
rect 38948 17054 39068 17082
rect 39120 17128 39172 17134
rect 39120 17070 39172 17076
rect 38752 16584 38804 16590
rect 38752 16526 38804 16532
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38764 15094 38792 16526
rect 38948 15638 38976 17054
rect 39028 15904 39080 15910
rect 39028 15846 39080 15852
rect 38936 15632 38988 15638
rect 38936 15574 38988 15580
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 38568 14272 38620 14278
rect 38568 14214 38620 14220
rect 38292 14068 38344 14074
rect 38292 14010 38344 14016
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 37740 13864 37792 13870
rect 37740 13806 37792 13812
rect 38568 13864 38620 13870
rect 38568 13806 38620 13812
rect 38580 13326 38608 13806
rect 38672 13530 38700 13942
rect 38764 13802 38792 15030
rect 39040 14890 39068 15846
rect 39028 14884 39080 14890
rect 39028 14826 39080 14832
rect 39040 13938 39068 14826
rect 39132 14414 39160 17070
rect 39224 16590 39252 18226
rect 39304 18216 39356 18222
rect 39304 18158 39356 18164
rect 39212 16584 39264 16590
rect 39212 16526 39264 16532
rect 39224 16182 39252 16526
rect 39212 16176 39264 16182
rect 39212 16118 39264 16124
rect 39316 16114 39344 18158
rect 39408 17338 39436 22578
rect 39488 22500 39540 22506
rect 39488 22442 39540 22448
rect 39500 17542 39528 22442
rect 39592 21554 39620 25162
rect 39684 24750 39712 26318
rect 39672 24744 39724 24750
rect 39672 24686 39724 24692
rect 39672 24200 39724 24206
rect 39672 24142 39724 24148
rect 39684 23866 39712 24142
rect 39672 23860 39724 23866
rect 39672 23802 39724 23808
rect 39776 23746 39804 26812
rect 39684 23718 39804 23746
rect 39684 22982 39712 23718
rect 39764 23044 39816 23050
rect 39764 22986 39816 22992
rect 39672 22976 39724 22982
rect 39672 22918 39724 22924
rect 39670 22808 39726 22817
rect 39670 22743 39726 22752
rect 39684 22710 39712 22743
rect 39672 22704 39724 22710
rect 39672 22646 39724 22652
rect 39684 22137 39712 22646
rect 39670 22128 39726 22137
rect 39670 22063 39726 22072
rect 39672 21888 39724 21894
rect 39672 21830 39724 21836
rect 39580 21548 39632 21554
rect 39580 21490 39632 21496
rect 39684 21350 39712 21830
rect 39672 21344 39724 21350
rect 39672 21286 39724 21292
rect 39672 19440 39724 19446
rect 39670 19408 39672 19417
rect 39724 19408 39726 19417
rect 39670 19343 39726 19352
rect 39672 19304 39724 19310
rect 39672 19246 39724 19252
rect 39684 18902 39712 19246
rect 39776 19242 39804 22986
rect 39868 21146 39896 26880
rect 39960 26382 39988 27542
rect 40040 26988 40092 26994
rect 40040 26930 40092 26936
rect 40052 26450 40080 26930
rect 40040 26444 40092 26450
rect 40040 26386 40092 26392
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 40040 26036 40092 26042
rect 40040 25978 40092 25984
rect 40052 25430 40080 25978
rect 40040 25424 40092 25430
rect 40040 25366 40092 25372
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40052 24818 40080 25230
rect 40144 24818 40172 30194
rect 40236 28558 40264 30670
rect 40420 29714 40448 31436
rect 40500 31340 40552 31346
rect 40500 31282 40552 31288
rect 40512 30122 40540 31282
rect 40604 30326 40632 31719
rect 40788 31328 40816 32370
rect 40880 31793 40908 32846
rect 40972 32570 41000 32982
rect 41340 32978 41368 33934
rect 41432 33522 41460 34070
rect 41616 33658 41644 40326
rect 41800 36650 41828 40870
rect 41880 40520 41932 40526
rect 41880 40462 41932 40468
rect 41892 39438 41920 40462
rect 41880 39432 41932 39438
rect 41880 39374 41932 39380
rect 41892 38350 41920 39374
rect 41880 38344 41932 38350
rect 41880 38286 41932 38292
rect 41892 37262 41920 38286
rect 42064 37664 42116 37670
rect 42064 37606 42116 37612
rect 41880 37256 41932 37262
rect 41880 37198 41932 37204
rect 41788 36644 41840 36650
rect 41788 36586 41840 36592
rect 41696 36236 41748 36242
rect 41696 36178 41748 36184
rect 41604 33652 41656 33658
rect 41604 33594 41656 33600
rect 41420 33516 41472 33522
rect 41420 33458 41472 33464
rect 41604 33380 41656 33386
rect 41604 33322 41656 33328
rect 41616 32978 41644 33322
rect 41052 32972 41104 32978
rect 41052 32914 41104 32920
rect 41328 32972 41380 32978
rect 41328 32914 41380 32920
rect 41604 32972 41656 32978
rect 41604 32914 41656 32920
rect 40960 32564 41012 32570
rect 40960 32506 41012 32512
rect 40866 31784 40922 31793
rect 40866 31719 40922 31728
rect 40960 31340 41012 31346
rect 40788 31300 40908 31328
rect 40880 31142 40908 31300
rect 40960 31282 41012 31288
rect 40868 31136 40920 31142
rect 40868 31078 40920 31084
rect 40880 30734 40908 31078
rect 40972 30870 41000 31282
rect 40960 30864 41012 30870
rect 40960 30806 41012 30812
rect 40684 30728 40736 30734
rect 40684 30670 40736 30676
rect 40868 30728 40920 30734
rect 40868 30670 40920 30676
rect 40592 30320 40644 30326
rect 40592 30262 40644 30268
rect 40500 30116 40552 30122
rect 40500 30058 40552 30064
rect 40316 29708 40368 29714
rect 40316 29650 40368 29656
rect 40408 29708 40460 29714
rect 40408 29650 40460 29656
rect 40328 29238 40356 29650
rect 40316 29232 40368 29238
rect 40316 29174 40368 29180
rect 40420 29170 40448 29650
rect 40408 29164 40460 29170
rect 40408 29106 40460 29112
rect 40512 29050 40540 30058
rect 40592 29776 40644 29782
rect 40592 29718 40644 29724
rect 40328 29022 40540 29050
rect 40604 29034 40632 29718
rect 40592 29028 40644 29034
rect 40224 28552 40276 28558
rect 40224 28494 40276 28500
rect 40328 27441 40356 29022
rect 40592 28970 40644 28976
rect 40500 28960 40552 28966
rect 40500 28902 40552 28908
rect 40408 28008 40460 28014
rect 40408 27950 40460 27956
rect 40420 27674 40448 27950
rect 40512 27674 40540 28902
rect 40696 28422 40724 30670
rect 40868 30388 40920 30394
rect 40868 30330 40920 30336
rect 40776 29232 40828 29238
rect 40776 29174 40828 29180
rect 40684 28416 40736 28422
rect 40684 28358 40736 28364
rect 40592 28076 40644 28082
rect 40592 28018 40644 28024
rect 40408 27668 40460 27674
rect 40408 27610 40460 27616
rect 40500 27668 40552 27674
rect 40500 27610 40552 27616
rect 40314 27432 40370 27441
rect 40224 27396 40276 27402
rect 40314 27367 40370 27376
rect 40224 27338 40276 27344
rect 40236 26994 40264 27338
rect 40224 26988 40276 26994
rect 40224 26930 40276 26936
rect 40316 26920 40368 26926
rect 40316 26862 40368 26868
rect 40224 26784 40276 26790
rect 40224 26726 40276 26732
rect 40040 24812 40092 24818
rect 40040 24754 40092 24760
rect 40132 24812 40184 24818
rect 40132 24754 40184 24760
rect 40038 24440 40094 24449
rect 40038 24375 40040 24384
rect 40092 24375 40094 24384
rect 40040 24346 40092 24352
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39960 22166 39988 22918
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 39948 22160 40000 22166
rect 39948 22102 40000 22108
rect 40052 21622 40080 22374
rect 40040 21616 40092 21622
rect 40040 21558 40092 21564
rect 39856 21140 39908 21146
rect 39856 21082 39908 21088
rect 40040 21140 40092 21146
rect 40040 21082 40092 21088
rect 39764 19236 39816 19242
rect 39764 19178 39816 19184
rect 39672 18896 39724 18902
rect 39672 18838 39724 18844
rect 39488 17536 39540 17542
rect 39488 17478 39540 17484
rect 39396 17332 39448 17338
rect 39396 17274 39448 17280
rect 39868 16794 39896 21082
rect 39948 19712 40000 19718
rect 39948 19654 40000 19660
rect 39960 19446 39988 19654
rect 39948 19440 40000 19446
rect 39948 19382 40000 19388
rect 40052 19242 40080 21082
rect 40144 21026 40172 24142
rect 40236 23322 40264 26726
rect 40328 26042 40356 26862
rect 40420 26382 40448 27610
rect 40500 27328 40552 27334
rect 40500 27270 40552 27276
rect 40512 26382 40540 27270
rect 40408 26376 40460 26382
rect 40408 26318 40460 26324
rect 40500 26376 40552 26382
rect 40500 26318 40552 26324
rect 40316 26036 40368 26042
rect 40316 25978 40368 25984
rect 40500 25900 40552 25906
rect 40500 25842 40552 25848
rect 40512 25430 40540 25842
rect 40500 25424 40552 25430
rect 40500 25366 40552 25372
rect 40512 24818 40540 25366
rect 40316 24812 40368 24818
rect 40316 24754 40368 24760
rect 40500 24812 40552 24818
rect 40500 24754 40552 24760
rect 40328 24698 40356 24754
rect 40604 24698 40632 28018
rect 40696 27130 40724 28358
rect 40684 27124 40736 27130
rect 40684 27066 40736 27072
rect 40696 26382 40724 27066
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 40788 24732 40816 29174
rect 40880 28218 40908 30330
rect 40972 29102 41000 30806
rect 41064 29306 41092 32914
rect 41144 32836 41196 32842
rect 41144 32778 41196 32784
rect 41156 30394 41184 32778
rect 41236 32496 41288 32502
rect 41236 32438 41288 32444
rect 41248 31890 41276 32438
rect 41604 32428 41656 32434
rect 41604 32370 41656 32376
rect 41616 31929 41644 32370
rect 41602 31920 41658 31929
rect 41236 31884 41288 31890
rect 41602 31855 41658 31864
rect 41236 31826 41288 31832
rect 41708 31804 41736 36178
rect 41892 36174 41920 37198
rect 41972 37188 42024 37194
rect 41972 37130 42024 37136
rect 41984 36922 42012 37130
rect 41972 36916 42024 36922
rect 41972 36858 42024 36864
rect 41880 36168 41932 36174
rect 41880 36110 41932 36116
rect 41788 36032 41840 36038
rect 41788 35974 41840 35980
rect 41800 35698 41828 35974
rect 41788 35692 41840 35698
rect 41788 35634 41840 35640
rect 41880 33856 41932 33862
rect 41880 33798 41932 33804
rect 41892 33318 41920 33798
rect 41880 33312 41932 33318
rect 41880 33254 41932 33260
rect 42076 32570 42104 37606
rect 42168 34406 42196 41550
rect 42616 41472 42668 41478
rect 42616 41414 42668 41420
rect 42536 41386 42656 41414
rect 42340 40384 42392 40390
rect 42340 40326 42392 40332
rect 42248 36576 42300 36582
rect 42248 36518 42300 36524
rect 42156 34400 42208 34406
rect 42156 34342 42208 34348
rect 42156 33924 42208 33930
rect 42156 33866 42208 33872
rect 42064 32564 42116 32570
rect 42064 32506 42116 32512
rect 41880 32020 41932 32026
rect 41880 31962 41932 31968
rect 41616 31776 41736 31804
rect 41420 31680 41472 31686
rect 41420 31622 41472 31628
rect 41432 31346 41460 31622
rect 41328 31340 41380 31346
rect 41248 31300 41328 31328
rect 41248 30802 41276 31300
rect 41328 31282 41380 31288
rect 41420 31340 41472 31346
rect 41420 31282 41472 31288
rect 41236 30796 41288 30802
rect 41236 30738 41288 30744
rect 41144 30388 41196 30394
rect 41144 30330 41196 30336
rect 41144 29708 41196 29714
rect 41144 29650 41196 29656
rect 41156 29306 41184 29650
rect 41052 29300 41104 29306
rect 41052 29242 41104 29248
rect 41144 29300 41196 29306
rect 41144 29242 41196 29248
rect 41052 29164 41104 29170
rect 41104 29124 41184 29152
rect 41052 29106 41104 29112
rect 40960 29096 41012 29102
rect 40960 29038 41012 29044
rect 41052 28960 41104 28966
rect 41052 28902 41104 28908
rect 41064 28694 41092 28902
rect 41052 28688 41104 28694
rect 41052 28630 41104 28636
rect 40868 28212 40920 28218
rect 40868 28154 40920 28160
rect 41064 28014 41092 28630
rect 41052 28008 41104 28014
rect 41052 27950 41104 27956
rect 41156 27962 41184 29124
rect 41248 28082 41276 30738
rect 41328 30592 41380 30598
rect 41328 30534 41380 30540
rect 41340 30394 41368 30534
rect 41328 30388 41380 30394
rect 41328 30330 41380 30336
rect 41420 30320 41472 30326
rect 41420 30262 41472 30268
rect 41328 29844 41380 29850
rect 41328 29786 41380 29792
rect 41340 29578 41368 29786
rect 41432 29714 41460 30262
rect 41420 29708 41472 29714
rect 41420 29650 41472 29656
rect 41512 29640 41564 29646
rect 41512 29582 41564 29588
rect 41328 29572 41380 29578
rect 41328 29514 41380 29520
rect 41340 28694 41368 29514
rect 41420 29164 41472 29170
rect 41420 29106 41472 29112
rect 41328 28688 41380 28694
rect 41328 28630 41380 28636
rect 41432 28626 41460 29106
rect 41524 29102 41552 29582
rect 41512 29096 41564 29102
rect 41512 29038 41564 29044
rect 41420 28620 41472 28626
rect 41420 28562 41472 28568
rect 41236 28076 41288 28082
rect 41236 28018 41288 28024
rect 41064 27470 41092 27950
rect 41156 27934 41368 27962
rect 41144 27600 41196 27606
rect 41144 27542 41196 27548
rect 40868 27464 40920 27470
rect 40868 27406 40920 27412
rect 41052 27464 41104 27470
rect 41052 27406 41104 27412
rect 40880 26926 40908 27406
rect 40960 26988 41012 26994
rect 40960 26930 41012 26936
rect 40868 26920 40920 26926
rect 40868 26862 40920 26868
rect 40972 26382 41000 26930
rect 41052 26444 41104 26450
rect 41052 26386 41104 26392
rect 40960 26376 41012 26382
rect 40960 26318 41012 26324
rect 41064 25974 41092 26386
rect 41052 25968 41104 25974
rect 41052 25910 41104 25916
rect 41156 24818 41184 27542
rect 41236 27532 41288 27538
rect 41236 27474 41288 27480
rect 41248 26790 41276 27474
rect 41340 27334 41368 27934
rect 41432 27674 41460 28562
rect 41420 27668 41472 27674
rect 41420 27610 41472 27616
rect 41328 27328 41380 27334
rect 41328 27270 41380 27276
rect 41236 26784 41288 26790
rect 41236 26726 41288 26732
rect 41248 26246 41276 26726
rect 41236 26240 41288 26246
rect 41236 26182 41288 26188
rect 41248 26042 41276 26182
rect 41236 26036 41288 26042
rect 41236 25978 41288 25984
rect 41248 25362 41276 25978
rect 41236 25356 41288 25362
rect 41236 25298 41288 25304
rect 41144 24812 41196 24818
rect 41144 24754 41196 24760
rect 40328 24676 40632 24698
rect 40328 24670 40500 24676
rect 40552 24670 40632 24676
rect 40696 24704 40816 24732
rect 40500 24618 40552 24624
rect 40406 24440 40462 24449
rect 40406 24375 40408 24384
rect 40460 24375 40462 24384
rect 40408 24346 40460 24352
rect 40696 23866 40724 24704
rect 40958 24168 41014 24177
rect 40958 24103 41014 24112
rect 40972 24070 41000 24103
rect 40960 24064 41012 24070
rect 40960 24006 41012 24012
rect 40684 23860 40736 23866
rect 40684 23802 40736 23808
rect 40696 23662 40724 23802
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 41156 23594 41184 24754
rect 41248 24750 41276 25298
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 41248 24410 41276 24686
rect 41236 24404 41288 24410
rect 41236 24346 41288 24352
rect 41340 24274 41368 27270
rect 41432 26926 41460 27610
rect 41512 27464 41564 27470
rect 41512 27406 41564 27412
rect 41524 26994 41552 27406
rect 41512 26988 41564 26994
rect 41512 26930 41564 26936
rect 41420 26920 41472 26926
rect 41420 26862 41472 26868
rect 41432 25820 41460 26862
rect 41512 25832 41564 25838
rect 41432 25792 41512 25820
rect 41512 25774 41564 25780
rect 41524 25294 41552 25774
rect 41512 25288 41564 25294
rect 41512 25230 41564 25236
rect 41328 24268 41380 24274
rect 41328 24210 41380 24216
rect 41512 23724 41564 23730
rect 41512 23666 41564 23672
rect 41144 23588 41196 23594
rect 41144 23530 41196 23536
rect 41524 23322 41552 23666
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 41512 23316 41564 23322
rect 41512 23258 41564 23264
rect 40868 22636 40920 22642
rect 40868 22578 40920 22584
rect 40408 22500 40460 22506
rect 40408 22442 40460 22448
rect 40316 22092 40368 22098
rect 40316 22034 40368 22040
rect 40224 22024 40276 22030
rect 40224 21966 40276 21972
rect 40236 21146 40264 21966
rect 40328 21554 40356 22034
rect 40316 21548 40368 21554
rect 40316 21490 40368 21496
rect 40224 21140 40276 21146
rect 40224 21082 40276 21088
rect 40144 20998 40264 21026
rect 40132 20936 40184 20942
rect 40132 20878 40184 20884
rect 40144 20602 40172 20878
rect 40132 20596 40184 20602
rect 40132 20538 40184 20544
rect 40236 20482 40264 20998
rect 40328 20602 40356 21490
rect 40420 20874 40448 22442
rect 40684 21888 40736 21894
rect 40684 21830 40736 21836
rect 40696 21622 40724 21830
rect 40880 21690 40908 22578
rect 41326 22128 41382 22137
rect 41616 22094 41644 31776
rect 41892 31482 41920 31962
rect 41880 31476 41932 31482
rect 41880 31418 41932 31424
rect 41696 31272 41748 31278
rect 41696 31214 41748 31220
rect 41708 30598 41736 31214
rect 41972 31136 42024 31142
rect 41972 31078 42024 31084
rect 41984 30734 42012 31078
rect 41972 30728 42024 30734
rect 41786 30696 41842 30705
rect 41972 30670 42024 30676
rect 41786 30631 41842 30640
rect 41696 30592 41748 30598
rect 41696 30534 41748 30540
rect 41708 30394 41736 30534
rect 41696 30388 41748 30394
rect 41696 30330 41748 30336
rect 41696 28484 41748 28490
rect 41696 28426 41748 28432
rect 41708 25974 41736 28426
rect 41800 28218 41828 30631
rect 42064 30116 42116 30122
rect 42064 30058 42116 30064
rect 41880 28960 41932 28966
rect 41880 28902 41932 28908
rect 41972 28960 42024 28966
rect 41972 28902 42024 28908
rect 41892 28558 41920 28902
rect 41984 28558 42012 28902
rect 41880 28552 41932 28558
rect 41880 28494 41932 28500
rect 41972 28552 42024 28558
rect 41972 28494 42024 28500
rect 41788 28212 41840 28218
rect 41788 28154 41840 28160
rect 41788 27396 41840 27402
rect 41788 27338 41840 27344
rect 41800 26382 41828 27338
rect 41892 26874 41920 28494
rect 41984 28014 42012 28494
rect 41972 28008 42024 28014
rect 41972 27950 42024 27956
rect 42076 27606 42104 30058
rect 42064 27600 42116 27606
rect 42064 27542 42116 27548
rect 41892 26846 42012 26874
rect 41880 26444 41932 26450
rect 41880 26386 41932 26392
rect 41788 26376 41840 26382
rect 41788 26318 41840 26324
rect 41696 25968 41748 25974
rect 41696 25910 41748 25916
rect 41708 25786 41736 25910
rect 41708 25758 41828 25786
rect 41696 25696 41748 25702
rect 41696 25638 41748 25644
rect 41708 24274 41736 25638
rect 41800 24886 41828 25758
rect 41892 25430 41920 26386
rect 41984 26314 42012 26846
rect 41972 26308 42024 26314
rect 41972 26250 42024 26256
rect 41880 25424 41932 25430
rect 41880 25366 41932 25372
rect 41788 24880 41840 24886
rect 41788 24822 41840 24828
rect 41892 24614 41920 25366
rect 41984 25276 42012 26250
rect 42168 25514 42196 33866
rect 42260 29782 42288 36518
rect 42352 36378 42380 40326
rect 42536 36718 42564 41386
rect 42616 40928 42668 40934
rect 42616 40870 42668 40876
rect 42628 40458 42656 40870
rect 42616 40452 42668 40458
rect 42616 40394 42668 40400
rect 42708 39908 42760 39914
rect 42708 39850 42760 39856
rect 42616 39840 42668 39846
rect 42616 39782 42668 39788
rect 42628 39098 42656 39782
rect 42616 39092 42668 39098
rect 42616 39034 42668 39040
rect 42614 37768 42670 37777
rect 42614 37703 42670 37712
rect 42524 36712 42576 36718
rect 42524 36654 42576 36660
rect 42628 36378 42656 37703
rect 42340 36372 42392 36378
rect 42340 36314 42392 36320
rect 42616 36372 42668 36378
rect 42616 36314 42668 36320
rect 42616 36100 42668 36106
rect 42616 36042 42668 36048
rect 42628 35834 42656 36042
rect 42720 35834 42748 39850
rect 42616 35828 42668 35834
rect 42616 35770 42668 35776
rect 42708 35828 42760 35834
rect 42708 35770 42760 35776
rect 42720 34746 42748 35770
rect 42708 34740 42760 34746
rect 42708 34682 42760 34688
rect 42720 34626 42748 34682
rect 42628 34598 42748 34626
rect 42812 34610 42840 42094
rect 43548 41614 43576 44200
rect 43994 42664 44050 42673
rect 43994 42599 44050 42608
rect 44008 42226 44036 42599
rect 43996 42220 44048 42226
rect 43996 42162 44048 42168
rect 43536 41608 43588 41614
rect 43536 41550 43588 41556
rect 43076 41540 43128 41546
rect 43076 41482 43128 41488
rect 42892 41472 42944 41478
rect 42892 41414 42944 41420
rect 42904 41274 42932 41414
rect 43088 41274 43116 41482
rect 42892 41268 42944 41274
rect 42892 41210 42944 41216
rect 43076 41268 43128 41274
rect 43076 41210 43128 41216
rect 42892 40384 42944 40390
rect 42892 40326 42944 40332
rect 42904 35737 42932 40326
rect 43444 39840 43496 39846
rect 43444 39782 43496 39788
rect 43352 36780 43404 36786
rect 43352 36722 43404 36728
rect 43364 36689 43392 36722
rect 43350 36680 43406 36689
rect 43350 36615 43406 36624
rect 42984 36576 43036 36582
rect 42984 36518 43036 36524
rect 42890 35728 42946 35737
rect 42890 35663 42946 35672
rect 42800 34604 42852 34610
rect 42432 33312 42484 33318
rect 42432 33254 42484 33260
rect 42444 31754 42472 33254
rect 42432 31748 42484 31754
rect 42432 31690 42484 31696
rect 42628 30705 42656 34598
rect 42800 34546 42852 34552
rect 42708 34536 42760 34542
rect 42708 34478 42760 34484
rect 42720 32910 42748 34478
rect 42812 33930 42840 34546
rect 42800 33924 42852 33930
rect 42800 33866 42852 33872
rect 42812 33522 42840 33866
rect 42800 33516 42852 33522
rect 42800 33458 42852 33464
rect 42904 33436 42932 35663
rect 42996 33930 43024 36518
rect 43076 34468 43128 34474
rect 43076 34410 43128 34416
rect 42984 33924 43036 33930
rect 42984 33866 43036 33872
rect 42996 33590 43024 33866
rect 43088 33658 43116 34410
rect 43168 33992 43220 33998
rect 43168 33934 43220 33940
rect 43076 33652 43128 33658
rect 43076 33594 43128 33600
rect 42984 33584 43036 33590
rect 42984 33526 43036 33532
rect 42904 33408 43024 33436
rect 42800 32972 42852 32978
rect 42800 32914 42852 32920
rect 42708 32904 42760 32910
rect 42708 32846 42760 32852
rect 42708 31272 42760 31278
rect 42706 31240 42708 31249
rect 42760 31240 42762 31249
rect 42706 31175 42762 31184
rect 42720 30802 42748 31175
rect 42812 31142 42840 32914
rect 42892 32224 42944 32230
rect 42892 32166 42944 32172
rect 42904 31890 42932 32166
rect 42892 31884 42944 31890
rect 42892 31826 42944 31832
rect 42892 31340 42944 31346
rect 42892 31282 42944 31288
rect 42800 31136 42852 31142
rect 42800 31078 42852 31084
rect 42798 30832 42854 30841
rect 42708 30796 42760 30802
rect 42798 30767 42800 30776
rect 42708 30738 42760 30744
rect 42852 30767 42854 30776
rect 42800 30738 42852 30744
rect 42614 30696 42670 30705
rect 42904 30682 42932 31282
rect 42614 30631 42670 30640
rect 42812 30654 42932 30682
rect 42812 30054 42840 30654
rect 42890 30288 42946 30297
rect 42890 30223 42946 30232
rect 42800 30048 42852 30054
rect 42800 29990 42852 29996
rect 42248 29776 42300 29782
rect 42300 29724 42380 29730
rect 42248 29718 42380 29724
rect 42260 29702 42380 29718
rect 42248 29572 42300 29578
rect 42248 29514 42300 29520
rect 42260 29170 42288 29514
rect 42248 29164 42300 29170
rect 42248 29106 42300 29112
rect 42168 25486 42288 25514
rect 42064 25288 42116 25294
rect 41984 25248 42064 25276
rect 42064 25230 42116 25236
rect 41972 25152 42024 25158
rect 41972 25094 42024 25100
rect 41984 24818 42012 25094
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 41880 24608 41932 24614
rect 41880 24550 41932 24556
rect 41696 24268 41748 24274
rect 41696 24210 41748 24216
rect 41708 24138 41736 24210
rect 41788 24200 41840 24206
rect 41788 24142 41840 24148
rect 41696 24132 41748 24138
rect 41696 24074 41748 24080
rect 41800 23322 41828 24142
rect 41788 23316 41840 23322
rect 41788 23258 41840 23264
rect 41800 22710 41828 23258
rect 41892 23118 41920 24550
rect 41984 23186 42012 24754
rect 42076 24410 42104 25230
rect 42064 24404 42116 24410
rect 42064 24346 42116 24352
rect 41972 23180 42024 23186
rect 41972 23122 42024 23128
rect 41880 23112 41932 23118
rect 41880 23054 41932 23060
rect 41788 22704 41840 22710
rect 41788 22646 41840 22652
rect 42064 22704 42116 22710
rect 42064 22646 42116 22652
rect 41788 22432 41840 22438
rect 41788 22374 41840 22380
rect 41800 22098 41828 22374
rect 41326 22063 41382 22072
rect 41524 22066 41644 22094
rect 41788 22092 41840 22098
rect 40868 21684 40920 21690
rect 40868 21626 40920 21632
rect 40500 21616 40552 21622
rect 40500 21558 40552 21564
rect 40684 21616 40736 21622
rect 40684 21558 40736 21564
rect 40512 21078 40540 21558
rect 40500 21072 40552 21078
rect 40500 21014 40552 21020
rect 40500 20936 40552 20942
rect 40500 20878 40552 20884
rect 40408 20868 40460 20874
rect 40408 20810 40460 20816
rect 40316 20596 40368 20602
rect 40316 20538 40368 20544
rect 40144 20454 40264 20482
rect 40144 19514 40172 20454
rect 40328 19922 40356 20538
rect 40420 19990 40448 20810
rect 40512 20398 40540 20878
rect 41340 20874 41368 22063
rect 41328 20868 41380 20874
rect 41328 20810 41380 20816
rect 41340 20777 41368 20810
rect 41326 20768 41382 20777
rect 41326 20703 41382 20712
rect 40500 20392 40552 20398
rect 40500 20334 40552 20340
rect 40512 20058 40540 20334
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 40408 19984 40460 19990
rect 40408 19926 40460 19932
rect 40316 19916 40368 19922
rect 40316 19858 40368 19864
rect 40132 19508 40184 19514
rect 40132 19450 40184 19456
rect 40774 19408 40830 19417
rect 40132 19372 40184 19378
rect 40132 19314 40184 19320
rect 40684 19372 40736 19378
rect 40774 19343 40776 19352
rect 40684 19314 40736 19320
rect 40828 19343 40830 19352
rect 41052 19372 41104 19378
rect 40776 19314 40828 19320
rect 41052 19314 41104 19320
rect 40040 19236 40092 19242
rect 40040 19178 40092 19184
rect 40144 19122 40172 19314
rect 40316 19304 40368 19310
rect 40316 19246 40368 19252
rect 39960 19094 40172 19122
rect 39960 18698 39988 19094
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 39948 18692 40000 18698
rect 39948 18634 40000 18640
rect 40144 17882 40172 18702
rect 40132 17876 40184 17882
rect 40052 17836 40132 17864
rect 39946 17776 40002 17785
rect 39946 17711 40002 17720
rect 39960 17066 39988 17711
rect 40052 17202 40080 17836
rect 40132 17818 40184 17824
rect 40236 17678 40264 18770
rect 40328 17678 40356 19246
rect 40696 18970 40724 19314
rect 40788 18970 40816 19314
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40684 18964 40736 18970
rect 40684 18906 40736 18912
rect 40776 18964 40828 18970
rect 40776 18906 40828 18912
rect 40788 18698 40816 18906
rect 40776 18692 40828 18698
rect 40776 18634 40828 18640
rect 40972 18358 41000 19110
rect 41064 18698 41092 19314
rect 41052 18692 41104 18698
rect 41052 18634 41104 18640
rect 40960 18352 41012 18358
rect 40960 18294 41012 18300
rect 40224 17672 40276 17678
rect 40224 17614 40276 17620
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 40132 17196 40184 17202
rect 40132 17138 40184 17144
rect 39948 17060 40000 17066
rect 39948 17002 40000 17008
rect 39856 16788 39908 16794
rect 39856 16730 39908 16736
rect 39304 16108 39356 16114
rect 39304 16050 39356 16056
rect 39856 16040 39908 16046
rect 39856 15982 39908 15988
rect 39210 15600 39266 15609
rect 39210 15535 39266 15544
rect 39224 15502 39252 15535
rect 39212 15496 39264 15502
rect 39212 15438 39264 15444
rect 39120 14408 39172 14414
rect 39120 14350 39172 14356
rect 39132 14006 39160 14350
rect 39120 14000 39172 14006
rect 39120 13942 39172 13948
rect 39028 13932 39080 13938
rect 39028 13874 39080 13880
rect 38752 13796 38804 13802
rect 38752 13738 38804 13744
rect 38660 13524 38712 13530
rect 38660 13466 38712 13472
rect 38764 13410 38792 13738
rect 38672 13382 38792 13410
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38580 12850 38608 13262
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 38568 12844 38620 12850
rect 38568 12786 38620 12792
rect 38580 12434 38608 12786
rect 38672 12782 38700 13382
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 38764 12986 38792 13262
rect 38752 12980 38804 12986
rect 38752 12922 38804 12928
rect 38660 12776 38712 12782
rect 38660 12718 38712 12724
rect 38660 12436 38712 12442
rect 38580 12406 38660 12434
rect 38660 12378 38712 12384
rect 38672 12238 38700 12378
rect 39224 12374 39252 15438
rect 39764 15020 39816 15026
rect 39764 14962 39816 14968
rect 39776 14482 39804 14962
rect 39868 14958 39896 15982
rect 40144 15094 40172 17138
rect 40236 16590 40264 17614
rect 40328 16590 40356 17614
rect 41064 17338 41092 18634
rect 41144 18624 41196 18630
rect 41144 18566 41196 18572
rect 41156 17678 41184 18566
rect 41328 18080 41380 18086
rect 41328 18022 41380 18028
rect 41340 17762 41368 18022
rect 41340 17746 41460 17762
rect 41340 17740 41472 17746
rect 41340 17734 41420 17740
rect 41420 17682 41472 17688
rect 41144 17672 41196 17678
rect 41144 17614 41196 17620
rect 41052 17332 41104 17338
rect 41052 17274 41104 17280
rect 41524 17270 41552 22066
rect 41788 22034 41840 22040
rect 42076 21690 42104 22646
rect 42260 22642 42288 25486
rect 42352 24070 42380 29702
rect 42616 29572 42668 29578
rect 42812 29560 42840 29990
rect 42904 29782 42932 30223
rect 42892 29776 42944 29782
rect 42892 29718 42944 29724
rect 42892 29572 42944 29578
rect 42812 29532 42892 29560
rect 42616 29514 42668 29520
rect 42892 29514 42944 29520
rect 42628 27470 42656 29514
rect 42800 28620 42852 28626
rect 42800 28562 42852 28568
rect 42812 28150 42840 28562
rect 42904 28558 42932 29514
rect 42996 28994 43024 33408
rect 43088 32570 43116 33594
rect 43076 32564 43128 32570
rect 43076 32506 43128 32512
rect 43180 31890 43208 33934
rect 43352 32564 43404 32570
rect 43352 32506 43404 32512
rect 43260 32428 43312 32434
rect 43260 32370 43312 32376
rect 43168 31884 43220 31890
rect 43168 31826 43220 31832
rect 43272 31754 43300 32370
rect 43180 31726 43300 31754
rect 42996 28966 43116 28994
rect 42984 28688 43036 28694
rect 42984 28630 43036 28636
rect 42892 28552 42944 28558
rect 42892 28494 42944 28500
rect 42800 28144 42852 28150
rect 42800 28086 42852 28092
rect 42616 27464 42668 27470
rect 42616 27406 42668 27412
rect 42628 27130 42656 27406
rect 42616 27124 42668 27130
rect 42616 27066 42668 27072
rect 42432 26784 42484 26790
rect 42432 26726 42484 26732
rect 42444 25226 42472 26726
rect 42996 26194 43024 28630
rect 43088 27878 43116 28966
rect 43076 27872 43128 27878
rect 43076 27814 43128 27820
rect 43076 26988 43128 26994
rect 43076 26930 43128 26936
rect 43088 26450 43116 26930
rect 43076 26444 43128 26450
rect 43076 26386 43128 26392
rect 42996 26166 43116 26194
rect 43088 25945 43116 26166
rect 43074 25936 43130 25945
rect 42524 25900 42576 25906
rect 43074 25871 43130 25880
rect 42524 25842 42576 25848
rect 42432 25220 42484 25226
rect 42432 25162 42484 25168
rect 42444 24750 42472 25162
rect 42536 25158 42564 25842
rect 42800 25764 42852 25770
rect 42800 25706 42852 25712
rect 42616 25492 42668 25498
rect 42616 25434 42668 25440
rect 42524 25152 42576 25158
rect 42524 25094 42576 25100
rect 42628 24818 42656 25434
rect 42616 24812 42668 24818
rect 42616 24754 42668 24760
rect 42432 24744 42484 24750
rect 42432 24686 42484 24692
rect 42444 24206 42472 24686
rect 42432 24200 42484 24206
rect 42432 24142 42484 24148
rect 42340 24064 42392 24070
rect 42340 24006 42392 24012
rect 42340 23792 42392 23798
rect 42340 23734 42392 23740
rect 42352 22778 42380 23734
rect 42444 23050 42472 24142
rect 42524 24064 42576 24070
rect 42524 24006 42576 24012
rect 42432 23044 42484 23050
rect 42432 22986 42484 22992
rect 42340 22772 42392 22778
rect 42340 22714 42392 22720
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 42156 22432 42208 22438
rect 42156 22374 42208 22380
rect 42168 21962 42196 22374
rect 42156 21956 42208 21962
rect 42156 21898 42208 21904
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 42260 21554 42288 22578
rect 42536 22234 42564 24006
rect 42812 23730 42840 25706
rect 42984 25696 43036 25702
rect 42984 25638 43036 25644
rect 42996 24886 43024 25638
rect 42984 24880 43036 24886
rect 42984 24822 43036 24828
rect 43088 24818 43116 25871
rect 42892 24812 42944 24818
rect 42892 24754 42944 24760
rect 43076 24812 43128 24818
rect 43076 24754 43128 24760
rect 42904 24274 42932 24754
rect 42892 24268 42944 24274
rect 42892 24210 42944 24216
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42904 23322 42932 24210
rect 43180 24154 43208 31726
rect 43260 31136 43312 31142
rect 43260 31078 43312 31084
rect 43272 30258 43300 31078
rect 43260 30252 43312 30258
rect 43260 30194 43312 30200
rect 43272 29578 43300 30194
rect 43260 29572 43312 29578
rect 43260 29514 43312 29520
rect 43272 28626 43300 29514
rect 43260 28620 43312 28626
rect 43260 28562 43312 28568
rect 43364 27062 43392 32506
rect 43456 28082 43484 39782
rect 43996 36780 44048 36786
rect 43996 36722 44048 36728
rect 44008 35329 44036 36722
rect 43994 35320 44050 35329
rect 43994 35255 44050 35264
rect 43994 31648 44050 31657
rect 43994 31583 44050 31592
rect 44008 31278 44036 31583
rect 43996 31272 44048 31278
rect 43996 31214 44048 31220
rect 43444 28076 43496 28082
rect 43444 28018 43496 28024
rect 43996 28076 44048 28082
rect 43996 28018 44048 28024
rect 44008 27985 44036 28018
rect 43994 27976 44050 27985
rect 43994 27911 44050 27920
rect 43536 27872 43588 27878
rect 43536 27814 43588 27820
rect 43352 27056 43404 27062
rect 43352 26998 43404 27004
rect 43088 24126 43208 24154
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 42984 24064 43036 24070
rect 42984 24006 43036 24012
rect 42996 23866 43024 24006
rect 42984 23860 43036 23866
rect 42984 23802 43036 23808
rect 42892 23316 42944 23322
rect 42892 23258 42944 23264
rect 43088 23254 43116 24126
rect 43168 24064 43220 24070
rect 43168 24006 43220 24012
rect 43076 23248 43128 23254
rect 43076 23190 43128 23196
rect 42892 23180 42944 23186
rect 42892 23122 42944 23128
rect 42708 23112 42760 23118
rect 42708 23054 42760 23060
rect 42904 23066 42932 23122
rect 42720 22438 42748 23054
rect 42904 23038 43024 23066
rect 42996 22574 43024 23038
rect 43076 23044 43128 23050
rect 43076 22986 43128 22992
rect 43088 22642 43116 22986
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 42984 22568 43036 22574
rect 42984 22510 43036 22516
rect 42708 22432 42760 22438
rect 42708 22374 42760 22380
rect 42524 22228 42576 22234
rect 42524 22170 42576 22176
rect 42248 21548 42300 21554
rect 42248 21490 42300 21496
rect 42260 20806 42288 21490
rect 42248 20800 42300 20806
rect 42248 20742 42300 20748
rect 41880 20528 41932 20534
rect 41880 20470 41932 20476
rect 41892 19514 41920 20470
rect 42260 20466 42288 20742
rect 42720 20602 42748 22374
rect 42996 22234 43024 22510
rect 42984 22228 43036 22234
rect 42984 22170 43036 22176
rect 42708 20596 42760 20602
rect 42708 20538 42760 20544
rect 42248 20460 42300 20466
rect 42248 20402 42300 20408
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 42260 19378 42288 20402
rect 42892 20256 42944 20262
rect 42892 20198 42944 20204
rect 42904 19854 42932 20198
rect 42892 19848 42944 19854
rect 42892 19790 42944 19796
rect 42248 19372 42300 19378
rect 42248 19314 42300 19320
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 41696 18760 41748 18766
rect 41696 18702 41748 18708
rect 41708 18086 41736 18702
rect 41696 18080 41748 18086
rect 41696 18022 41748 18028
rect 41708 17270 41736 18022
rect 41512 17264 41564 17270
rect 41512 17206 41564 17212
rect 41696 17264 41748 17270
rect 41696 17206 41748 17212
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 40236 15910 40264 16526
rect 40224 15904 40276 15910
rect 40224 15846 40276 15852
rect 40132 15088 40184 15094
rect 40132 15030 40184 15036
rect 39856 14952 39908 14958
rect 39856 14894 39908 14900
rect 39868 14482 39896 14894
rect 40144 14618 40172 15030
rect 40236 14618 40264 15846
rect 40132 14612 40184 14618
rect 40132 14554 40184 14560
rect 40224 14612 40276 14618
rect 40224 14554 40276 14560
rect 39764 14476 39816 14482
rect 39764 14418 39816 14424
rect 39856 14476 39908 14482
rect 39856 14418 39908 14424
rect 39580 14408 39632 14414
rect 39580 14350 39632 14356
rect 39592 13938 39620 14350
rect 39776 13938 39804 14418
rect 40144 14414 40172 14554
rect 40132 14408 40184 14414
rect 40132 14350 40184 14356
rect 40328 14346 40356 16526
rect 41524 16522 41552 17206
rect 41708 16658 41736 17206
rect 41696 16652 41748 16658
rect 41696 16594 41748 16600
rect 41512 16516 41564 16522
rect 41512 16458 41564 16464
rect 41052 16448 41104 16454
rect 41052 16390 41104 16396
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 40972 15570 41000 16186
rect 40960 15564 41012 15570
rect 40960 15506 41012 15512
rect 41064 15366 41092 16390
rect 41236 16108 41288 16114
rect 41236 16050 41288 16056
rect 41144 15564 41196 15570
rect 41144 15506 41196 15512
rect 40500 15360 40552 15366
rect 40500 15302 40552 15308
rect 41052 15360 41104 15366
rect 41052 15302 41104 15308
rect 40316 14340 40368 14346
rect 40316 14282 40368 14288
rect 40512 14278 40540 15302
rect 41064 15026 41092 15302
rect 41052 15020 41104 15026
rect 41052 14962 41104 14968
rect 40592 14340 40644 14346
rect 40592 14282 40644 14288
rect 40500 14272 40552 14278
rect 40500 14214 40552 14220
rect 40512 13938 40540 14214
rect 39580 13932 39632 13938
rect 39580 13874 39632 13880
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 40040 13796 40092 13802
rect 40040 13738 40092 13744
rect 40052 13462 40080 13738
rect 40040 13456 40092 13462
rect 40040 13398 40092 13404
rect 40408 13252 40460 13258
rect 40408 13194 40460 13200
rect 39212 12368 39264 12374
rect 39212 12310 39264 12316
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 38660 12232 38712 12238
rect 38660 12174 38712 12180
rect 39396 12232 39448 12238
rect 39396 12174 39448 12180
rect 37648 12096 37700 12102
rect 37648 12038 37700 12044
rect 37372 11892 37424 11898
rect 37372 11834 37424 11840
rect 37280 11824 37332 11830
rect 37280 11766 37332 11772
rect 36912 11280 36964 11286
rect 36912 11222 36964 11228
rect 36924 10810 36952 11222
rect 37292 11150 37320 11766
rect 37660 11762 37688 12038
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37660 11218 37688 11698
rect 37648 11212 37700 11218
rect 37648 11154 37700 11160
rect 38304 11150 38332 12174
rect 38672 11762 38700 12174
rect 39118 12064 39174 12073
rect 39118 11999 39174 12008
rect 38660 11756 38712 11762
rect 38660 11698 38712 11704
rect 38384 11552 38436 11558
rect 38384 11494 38436 11500
rect 38396 11218 38424 11494
rect 38384 11212 38436 11218
rect 38384 11154 38436 11160
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 35440 10804 35492 10810
rect 35440 10746 35492 10752
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 37292 10742 37320 11086
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37936 10742 37964 10950
rect 37280 10736 37332 10742
rect 37280 10678 37332 10684
rect 37924 10736 37976 10742
rect 37924 10678 37976 10684
rect 31852 10532 31904 10538
rect 31852 10474 31904 10480
rect 34428 10532 34480 10538
rect 34428 10474 34480 10480
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 38304 10266 38332 11086
rect 39132 11014 39160 11999
rect 39408 11898 39436 12174
rect 39670 12064 39726 12073
rect 39670 11999 39726 12008
rect 39396 11892 39448 11898
rect 39396 11834 39448 11840
rect 39684 11830 39712 11999
rect 39672 11824 39724 11830
rect 39672 11766 39724 11772
rect 40040 11824 40092 11830
rect 40040 11766 40092 11772
rect 39120 11008 39172 11014
rect 39120 10950 39172 10956
rect 39396 11008 39448 11014
rect 39396 10950 39448 10956
rect 39028 10668 39080 10674
rect 39028 10610 39080 10616
rect 39040 10266 39068 10610
rect 38292 10260 38344 10266
rect 38292 10202 38344 10208
rect 39028 10260 39080 10266
rect 39028 10202 39080 10208
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 39408 10062 39436 10950
rect 40052 10266 40080 11766
rect 40132 11756 40184 11762
rect 40132 11698 40184 11704
rect 40144 11082 40172 11698
rect 40420 11150 40448 13194
rect 40604 12442 40632 14282
rect 41052 13864 41104 13870
rect 41052 13806 41104 13812
rect 41064 13190 41092 13806
rect 41156 13802 41184 15506
rect 41248 15162 41276 16050
rect 41328 15904 41380 15910
rect 41328 15846 41380 15852
rect 41340 15502 41368 15846
rect 41328 15496 41380 15502
rect 41328 15438 41380 15444
rect 41236 15156 41288 15162
rect 41236 15098 41288 15104
rect 41234 14104 41290 14113
rect 41234 14039 41236 14048
rect 41288 14039 41290 14048
rect 41236 14010 41288 14016
rect 41144 13796 41196 13802
rect 41144 13738 41196 13744
rect 41052 13184 41104 13190
rect 41052 13126 41104 13132
rect 41064 12986 41092 13126
rect 41052 12980 41104 12986
rect 41052 12922 41104 12928
rect 41156 12866 41184 13738
rect 41064 12838 41184 12866
rect 41248 12850 41276 14010
rect 41340 13326 41368 15438
rect 41524 14906 41552 16458
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 41616 15026 41644 15846
rect 41708 15570 41736 16594
rect 41696 15564 41748 15570
rect 41696 15506 41748 15512
rect 41604 15020 41656 15026
rect 41604 14962 41656 14968
rect 41524 14878 41736 14906
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 41420 12980 41472 12986
rect 41420 12922 41472 12928
rect 41236 12844 41288 12850
rect 41064 12782 41092 12838
rect 41236 12786 41288 12792
rect 41052 12776 41104 12782
rect 41052 12718 41104 12724
rect 40592 12436 40644 12442
rect 40592 12378 40644 12384
rect 40866 11928 40922 11937
rect 40866 11863 40868 11872
rect 40920 11863 40922 11872
rect 40868 11834 40920 11840
rect 40408 11144 40460 11150
rect 40408 11086 40460 11092
rect 40132 11076 40184 11082
rect 40132 11018 40184 11024
rect 40144 10810 40172 11018
rect 40132 10804 40184 10810
rect 40132 10746 40184 10752
rect 40420 10742 40448 11086
rect 40684 11076 40736 11082
rect 40684 11018 40736 11024
rect 40408 10736 40460 10742
rect 40408 10678 40460 10684
rect 40696 10266 40724 11018
rect 40880 10810 40908 11834
rect 41064 11694 41092 12718
rect 41248 12434 41276 12786
rect 41432 12434 41460 12922
rect 41512 12436 41564 12442
rect 41248 12406 41368 12434
rect 41432 12406 41512 12434
rect 41144 11756 41196 11762
rect 41144 11698 41196 11704
rect 41052 11688 41104 11694
rect 41052 11630 41104 11636
rect 41156 11354 41184 11698
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 41144 11348 41196 11354
rect 41144 11290 41196 11296
rect 41064 11082 41092 11290
rect 41052 11076 41104 11082
rect 41052 11018 41104 11024
rect 40868 10804 40920 10810
rect 40868 10746 40920 10752
rect 41064 10606 41092 11018
rect 41156 10810 41184 11290
rect 41144 10804 41196 10810
rect 41144 10746 41196 10752
rect 41052 10600 41104 10606
rect 41052 10542 41104 10548
rect 40868 10464 40920 10470
rect 40868 10406 40920 10412
rect 40040 10260 40092 10266
rect 40040 10202 40092 10208
rect 40684 10260 40736 10266
rect 40684 10202 40736 10208
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 39396 10056 39448 10062
rect 39396 9998 39448 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 40052 9722 40080 10202
rect 40880 10062 40908 10406
rect 40868 10056 40920 10062
rect 40868 9998 40920 10004
rect 40040 9716 40092 9722
rect 40040 9658 40092 9664
rect 40052 9382 40080 9658
rect 41340 9654 41368 12406
rect 41512 12378 41564 12384
rect 41420 10736 41472 10742
rect 41420 10678 41472 10684
rect 41328 9648 41380 9654
rect 41328 9590 41380 9596
rect 40040 9376 40092 9382
rect 40040 9318 40092 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 41432 9178 41460 10678
rect 41708 10470 41736 14878
rect 41800 14618 41828 18906
rect 42616 18760 42668 18766
rect 42616 18702 42668 18708
rect 42248 18624 42300 18630
rect 42248 18566 42300 18572
rect 41972 17740 42024 17746
rect 41972 17682 42024 17688
rect 41880 17332 41932 17338
rect 41880 17274 41932 17280
rect 41892 15162 41920 17274
rect 41984 15570 42012 17682
rect 42260 17678 42288 18566
rect 42628 18426 42656 18702
rect 42616 18420 42668 18426
rect 42616 18362 42668 18368
rect 43076 18216 43128 18222
rect 43076 18158 43128 18164
rect 42984 18148 43036 18154
rect 42984 18090 43036 18096
rect 42996 17882 43024 18090
rect 43088 17882 43116 18158
rect 42984 17876 43036 17882
rect 42984 17818 43036 17824
rect 43076 17876 43128 17882
rect 43076 17818 43128 17824
rect 42248 17672 42300 17678
rect 42248 17614 42300 17620
rect 42248 17196 42300 17202
rect 42248 17138 42300 17144
rect 41972 15564 42024 15570
rect 41972 15506 42024 15512
rect 41880 15156 41932 15162
rect 41880 15098 41932 15104
rect 41788 14612 41840 14618
rect 41788 14554 41840 14560
rect 41892 14006 41920 15098
rect 41880 14000 41932 14006
rect 41880 13942 41932 13948
rect 41892 12986 41920 13942
rect 41972 13320 42024 13326
rect 41972 13262 42024 13268
rect 41880 12980 41932 12986
rect 41880 12922 41932 12928
rect 41984 12306 42012 13262
rect 42156 13252 42208 13258
rect 42156 13194 42208 13200
rect 42168 12986 42196 13194
rect 42156 12980 42208 12986
rect 42156 12922 42208 12928
rect 41972 12300 42024 12306
rect 41972 12242 42024 12248
rect 42064 12164 42116 12170
rect 42064 12106 42116 12112
rect 42076 11898 42104 12106
rect 42064 11892 42116 11898
rect 42064 11834 42116 11840
rect 42260 10810 42288 17138
rect 42892 16652 42944 16658
rect 42892 16594 42944 16600
rect 42800 16448 42852 16454
rect 42800 16390 42852 16396
rect 42616 15428 42668 15434
rect 42616 15370 42668 15376
rect 42628 15162 42656 15370
rect 42616 15156 42668 15162
rect 42616 15098 42668 15104
rect 42812 15026 42840 16390
rect 42904 15706 42932 16594
rect 42996 16590 43024 17818
rect 43088 17338 43116 17818
rect 43076 17332 43128 17338
rect 43076 17274 43128 17280
rect 42984 16584 43036 16590
rect 42984 16526 43036 16532
rect 42996 15978 43024 16526
rect 43180 16182 43208 24006
rect 43260 22636 43312 22642
rect 43260 22578 43312 22584
rect 43272 20058 43300 22578
rect 43364 21690 43392 24142
rect 43352 21684 43404 21690
rect 43352 21626 43404 21632
rect 43352 20868 43404 20874
rect 43352 20810 43404 20816
rect 43260 20052 43312 20058
rect 43260 19994 43312 20000
rect 43168 16176 43220 16182
rect 43168 16118 43220 16124
rect 42984 15972 43036 15978
rect 42984 15914 43036 15920
rect 42892 15700 42944 15706
rect 42892 15642 42944 15648
rect 42996 15586 43024 15914
rect 42904 15558 43024 15586
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42904 13870 42932 15558
rect 43180 15502 43208 16118
rect 43168 15496 43220 15502
rect 43220 15456 43300 15484
rect 43168 15438 43220 15444
rect 43074 14376 43130 14385
rect 43074 14311 43076 14320
rect 43128 14311 43130 14320
rect 43076 14282 43128 14288
rect 43088 14074 43116 14282
rect 43076 14068 43128 14074
rect 42996 14028 43076 14056
rect 42892 13864 42944 13870
rect 42892 13806 42944 13812
rect 42798 13288 42854 13297
rect 42798 13223 42854 13232
rect 42524 12912 42576 12918
rect 42524 12854 42576 12860
rect 42536 12434 42564 12854
rect 42536 12406 42656 12434
rect 42628 11898 42656 12406
rect 42616 11892 42668 11898
rect 42616 11834 42668 11840
rect 42340 11756 42392 11762
rect 42340 11698 42392 11704
rect 42352 11354 42380 11698
rect 42340 11348 42392 11354
rect 42340 11290 42392 11296
rect 42248 10804 42300 10810
rect 42248 10746 42300 10752
rect 41696 10464 41748 10470
rect 41696 10406 41748 10412
rect 42064 10464 42116 10470
rect 42064 10406 42116 10412
rect 42076 10266 42104 10406
rect 42064 10260 42116 10266
rect 42064 10202 42116 10208
rect 42812 9654 42840 13223
rect 42904 12782 42932 13806
rect 42996 12986 43024 14028
rect 43076 14010 43128 14016
rect 43076 13864 43128 13870
rect 43076 13806 43128 13812
rect 43088 13530 43116 13806
rect 43168 13796 43220 13802
rect 43168 13738 43220 13744
rect 43076 13524 43128 13530
rect 43076 13466 43128 13472
rect 43088 12986 43116 13466
rect 42984 12980 43036 12986
rect 42984 12922 43036 12928
rect 43076 12980 43128 12986
rect 43076 12922 43128 12928
rect 42892 12776 42944 12782
rect 42892 12718 42944 12724
rect 42904 11218 42932 12718
rect 43076 12096 43128 12102
rect 43076 12038 43128 12044
rect 43088 11898 43116 12038
rect 43076 11892 43128 11898
rect 43076 11834 43128 11840
rect 42984 11756 43036 11762
rect 42984 11698 43036 11704
rect 42996 11354 43024 11698
rect 42984 11348 43036 11354
rect 42984 11290 43036 11296
rect 42892 11212 42944 11218
rect 42892 11154 42944 11160
rect 42996 10130 43024 11290
rect 43088 11286 43116 11834
rect 43180 11694 43208 13738
rect 43168 11688 43220 11694
rect 43168 11630 43220 11636
rect 43076 11280 43128 11286
rect 43076 11222 43128 11228
rect 42984 10124 43036 10130
rect 42984 10066 43036 10072
rect 42800 9648 42852 9654
rect 42800 9590 42852 9596
rect 42996 9466 43024 10066
rect 43272 9926 43300 15456
rect 43364 15162 43392 20810
rect 43548 18290 43576 27814
rect 43994 24304 44050 24313
rect 43994 24239 44050 24248
rect 44008 24206 44036 24239
rect 43996 24200 44048 24206
rect 43996 24142 44048 24148
rect 43996 20868 44048 20874
rect 43996 20810 44048 20816
rect 44008 20641 44036 20810
rect 43994 20632 44050 20641
rect 43994 20567 44050 20576
rect 43536 18284 43588 18290
rect 43536 18226 43588 18232
rect 43548 17610 43576 18226
rect 43536 17604 43588 17610
rect 43536 17546 43588 17552
rect 43548 17134 43576 17546
rect 43996 17196 44048 17202
rect 43996 17138 44048 17144
rect 43536 17128 43588 17134
rect 43536 17070 43588 17076
rect 43352 15156 43404 15162
rect 43352 15098 43404 15104
rect 43352 14408 43404 14414
rect 43352 14350 43404 14356
rect 43364 13297 43392 14350
rect 43350 13288 43406 13297
rect 43350 13223 43406 13232
rect 43352 12912 43404 12918
rect 43352 12854 43404 12860
rect 43260 9920 43312 9926
rect 43260 9862 43312 9868
rect 43272 9722 43300 9862
rect 43260 9716 43312 9722
rect 43260 9658 43312 9664
rect 42904 9438 43024 9466
rect 41420 9172 41472 9178
rect 41420 9114 41472 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 42904 8634 42932 9438
rect 42984 9376 43036 9382
rect 42984 9318 43036 9324
rect 42892 8628 42944 8634
rect 42892 8570 42944 8576
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 42996 2514 43024 9318
rect 43364 9178 43392 12854
rect 43548 10810 43576 17070
rect 44008 16969 44036 17138
rect 43994 16960 44050 16969
rect 43994 16895 44050 16904
rect 43536 10804 43588 10810
rect 43536 10746 43588 10752
rect 43996 10056 44048 10062
rect 43996 9998 44048 10004
rect 44008 9625 44036 9998
rect 43994 9616 44050 9625
rect 43994 9551 44050 9560
rect 43076 9172 43128 9178
rect 43076 9114 43128 9120
rect 43352 9172 43404 9178
rect 43352 9114 43404 9120
rect 43088 6390 43116 9114
rect 44008 8090 44036 9551
rect 43996 8084 44048 8090
rect 43996 8026 44048 8032
rect 43076 6384 43128 6390
rect 43076 6326 43128 6332
rect 43352 6316 43404 6322
rect 43352 6258 43404 6264
rect 43364 5953 43392 6258
rect 43350 5944 43406 5953
rect 43350 5879 43352 5888
rect 43404 5879 43406 5888
rect 43352 5850 43404 5856
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 42984 2508 43036 2514
rect 42984 2450 43036 2456
rect 43364 2446 43392 2790
rect 43352 2440 43404 2446
rect 43352 2382 43404 2388
rect 43996 2440 44048 2446
rect 43996 2382 44048 2388
rect 44008 2281 44036 2382
rect 43994 2272 44050 2281
rect 19574 2204 19882 2213
rect 43994 2207 44050 2216
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
<< via2 >>
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 10414 34584 10470 34640
rect 7562 34448 7618 34504
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 15198 37884 15200 37904
rect 15200 37884 15252 37904
rect 15252 37884 15254 37904
rect 15198 37848 15254 37884
rect 15566 37576 15622 37632
rect 14094 36644 14150 36680
rect 14094 36624 14096 36644
rect 14096 36624 14148 36644
rect 14148 36624 14150 36644
rect 12254 34992 12310 35048
rect 10690 33904 10746 33960
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 16946 38820 17002 38856
rect 16946 38800 16948 38820
rect 16948 38800 17000 38820
rect 17000 38800 17002 38820
rect 16670 37460 16726 37496
rect 16670 37440 16672 37460
rect 16672 37440 16724 37460
rect 16724 37440 16726 37460
rect 17222 38392 17278 38448
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 16486 31728 16542 31784
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19982 34856 20038 34912
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 17590 31728 17646 31784
rect 18142 31184 18198 31240
rect 18234 31048 18290 31104
rect 18142 29044 18144 29064
rect 18144 29044 18196 29064
rect 18196 29044 18198 29064
rect 18142 29008 18198 29044
rect 18418 29144 18474 29200
rect 18786 31048 18842 31104
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19430 33496 19486 33552
rect 18878 29588 18880 29608
rect 18880 29588 18932 29608
rect 18932 29588 18934 29608
rect 18878 29552 18934 29588
rect 18970 29008 19026 29064
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 20534 34468 20590 34504
rect 20534 34448 20536 34468
rect 20536 34448 20588 34468
rect 20588 34448 20590 34468
rect 20258 33496 20314 33552
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19982 31048 20038 31104
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 20810 34040 20866 34096
rect 21546 38256 21602 38312
rect 21454 37984 21510 38040
rect 22006 35808 22062 35864
rect 22098 35264 22154 35320
rect 22282 36896 22338 36952
rect 22558 37848 22614 37904
rect 22926 37984 22982 38040
rect 22282 36352 22338 36408
rect 23018 37848 23074 37904
rect 21454 34040 21510 34096
rect 20626 32816 20682 32872
rect 20534 32544 20590 32600
rect 19154 29552 19210 29608
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19982 29280 20038 29336
rect 20074 29144 20130 29200
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 21914 31728 21970 31784
rect 22098 30368 22154 30424
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 23202 36524 23204 36544
rect 23204 36524 23256 36544
rect 23256 36524 23258 36544
rect 23202 36488 23258 36524
rect 23570 38256 23626 38312
rect 23294 36216 23350 36272
rect 23570 37032 23626 37088
rect 24306 38120 24362 38176
rect 23754 36352 23810 36408
rect 24122 36352 24178 36408
rect 23938 35980 23940 36000
rect 23940 35980 23992 36000
rect 23992 35980 23994 36000
rect 23938 35944 23994 35980
rect 24030 35672 24086 35728
rect 23570 33088 23626 33144
rect 23846 32952 23902 33008
rect 24766 38292 24768 38312
rect 24768 38292 24820 38312
rect 24820 38292 24822 38312
rect 24766 38256 24822 38292
rect 24766 37304 24822 37360
rect 24766 36896 24822 36952
rect 25226 37712 25282 37768
rect 25502 38392 25558 38448
rect 25318 37304 25374 37360
rect 20534 26036 20590 26072
rect 20534 26016 20536 26036
rect 20536 26016 20588 26036
rect 20588 26016 20590 26036
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 17866 19216 17922 19272
rect 17222 17620 17224 17640
rect 17224 17620 17276 17640
rect 17276 17620 17278 17640
rect 17222 17584 17278 17620
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 22742 19508 22798 19544
rect 22742 19488 22744 19508
rect 22744 19488 22796 19508
rect 22796 19488 22798 19508
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 24306 32428 24362 32464
rect 24582 36116 24584 36136
rect 24584 36116 24636 36136
rect 24636 36116 24638 36136
rect 24582 36080 24638 36116
rect 24582 35808 24638 35864
rect 24674 35128 24730 35184
rect 24306 32408 24308 32428
rect 24308 32408 24360 32428
rect 24360 32408 24362 32428
rect 24674 32272 24730 32328
rect 25042 35264 25098 35320
rect 25502 36760 25558 36816
rect 25318 36100 25374 36136
rect 25318 36080 25320 36100
rect 25320 36080 25372 36100
rect 25372 36080 25374 36100
rect 25686 38156 25688 38176
rect 25688 38156 25740 38176
rect 25740 38156 25742 38176
rect 25686 38120 25742 38156
rect 25870 37984 25926 38040
rect 25870 37032 25926 37088
rect 25870 36780 25926 36816
rect 25870 36760 25872 36780
rect 25872 36760 25924 36780
rect 25924 36760 25926 36780
rect 25502 35944 25558 36000
rect 25778 35808 25834 35864
rect 25226 34312 25282 34368
rect 25594 34720 25650 34776
rect 25226 33768 25282 33824
rect 24950 32564 25006 32600
rect 24950 32544 24952 32564
rect 24952 32544 25004 32564
rect 25004 32544 25006 32564
rect 24398 29008 24454 29064
rect 24306 26288 24362 26344
rect 25226 32544 25282 32600
rect 25226 32272 25282 32328
rect 25410 32272 25466 32328
rect 25134 31764 25136 31784
rect 25136 31764 25188 31784
rect 25188 31764 25190 31784
rect 25134 31728 25190 31764
rect 25410 31864 25466 31920
rect 25042 31048 25098 31104
rect 24950 30776 25006 30832
rect 24582 29280 24638 29336
rect 26146 38392 26202 38448
rect 26238 38292 26240 38312
rect 26240 38292 26292 38312
rect 26292 38292 26294 38312
rect 26238 38256 26294 38292
rect 26054 33632 26110 33688
rect 26514 36488 26570 36544
rect 26974 37984 27030 38040
rect 26974 36760 27030 36816
rect 26422 36352 26478 36408
rect 26422 33904 26478 33960
rect 26330 33768 26386 33824
rect 25870 30252 25926 30288
rect 25870 30232 25872 30252
rect 25872 30232 25924 30252
rect 25924 30232 25926 30252
rect 26146 19932 26148 19952
rect 26148 19932 26200 19952
rect 26200 19932 26202 19952
rect 26146 19896 26202 19932
rect 24582 16788 24638 16824
rect 24582 16768 24584 16788
rect 24584 16768 24636 16788
rect 24636 16768 24638 16788
rect 26054 15308 26056 15328
rect 26056 15308 26108 15328
rect 26108 15308 26110 15328
rect 26054 15272 26110 15308
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 26882 32408 26938 32464
rect 27526 38972 27528 38992
rect 27528 38972 27580 38992
rect 27580 38972 27582 38992
rect 27526 38936 27582 38972
rect 27158 35400 27214 35456
rect 26790 31764 26792 31784
rect 26792 31764 26844 31784
rect 26844 31764 26846 31784
rect 26790 31728 26846 31764
rect 26698 27648 26754 27704
rect 26606 16244 26662 16280
rect 26606 16224 26608 16244
rect 26608 16224 26660 16244
rect 26660 16224 26662 16244
rect 27434 37576 27490 37632
rect 27342 35672 27398 35728
rect 27342 34992 27398 35048
rect 27894 39888 27950 39944
rect 28354 38428 28356 38448
rect 28356 38428 28408 38448
rect 28408 38428 28410 38448
rect 28354 38392 28410 38428
rect 28262 37848 28318 37904
rect 27710 36080 27766 36136
rect 27618 35944 27674 36000
rect 27526 35572 27528 35592
rect 27528 35572 27580 35592
rect 27580 35572 27582 35592
rect 27526 35536 27582 35572
rect 27342 34448 27398 34504
rect 27526 33360 27582 33416
rect 27342 31728 27398 31784
rect 27986 34176 28042 34232
rect 27894 30504 27950 30560
rect 27434 20596 27490 20632
rect 28354 35028 28356 35048
rect 28356 35028 28408 35048
rect 28408 35028 28410 35048
rect 28354 34992 28410 35028
rect 28170 32544 28226 32600
rect 28998 38800 29054 38856
rect 28906 38700 28908 38720
rect 28908 38700 28960 38720
rect 28960 38700 28962 38720
rect 28906 38664 28962 38700
rect 28630 38292 28632 38312
rect 28632 38292 28684 38312
rect 28684 38292 28686 38312
rect 28630 38256 28686 38292
rect 28906 38256 28962 38312
rect 28722 37984 28778 38040
rect 28630 35808 28686 35864
rect 28630 34856 28686 34912
rect 28998 37984 29054 38040
rect 29366 37848 29422 37904
rect 29274 37304 29330 37360
rect 28814 34176 28870 34232
rect 28998 34992 29054 35048
rect 28998 34584 29054 34640
rect 28998 33496 29054 33552
rect 29366 35808 29422 35864
rect 29734 37576 29790 37632
rect 29918 37204 29920 37224
rect 29920 37204 29972 37224
rect 29972 37204 29974 37224
rect 29918 37168 29974 37204
rect 30010 37032 30066 37088
rect 30378 38936 30434 38992
rect 31482 39888 31538 39944
rect 30286 37304 30342 37360
rect 30286 36080 30342 36136
rect 30010 35536 30066 35592
rect 29458 33940 29460 33960
rect 29460 33940 29512 33960
rect 29512 33940 29514 33960
rect 29458 33904 29514 33940
rect 28906 31764 28908 31784
rect 28908 31764 28960 31784
rect 28960 31764 28962 31784
rect 28906 31728 28962 31764
rect 28814 30252 28870 30288
rect 28814 30232 28816 30252
rect 28816 30232 28868 30252
rect 28868 30232 28870 30252
rect 29918 34584 29974 34640
rect 30194 35692 30250 35728
rect 30194 35672 30196 35692
rect 30196 35672 30248 35692
rect 30248 35672 30250 35692
rect 30654 35808 30710 35864
rect 30286 35536 30342 35592
rect 30562 34312 30618 34368
rect 30470 33632 30526 33688
rect 30378 33108 30434 33144
rect 30378 33088 30380 33108
rect 30380 33088 30432 33108
rect 30432 33088 30434 33108
rect 29734 31084 29736 31104
rect 29736 31084 29788 31104
rect 29788 31084 29790 31104
rect 29734 31048 29790 31084
rect 29734 30932 29790 30968
rect 29734 30912 29736 30932
rect 29736 30912 29788 30932
rect 29788 30912 29790 30932
rect 30010 31084 30012 31104
rect 30012 31084 30064 31104
rect 30064 31084 30066 31104
rect 30010 31048 30066 31084
rect 28354 24112 28410 24168
rect 27434 20576 27436 20596
rect 27436 20576 27488 20596
rect 27488 20576 27490 20596
rect 26974 14320 27030 14376
rect 27986 17720 28042 17776
rect 27894 16496 27950 16552
rect 29734 29008 29790 29064
rect 28998 22108 29000 22128
rect 29000 22108 29052 22128
rect 29052 22108 29054 22128
rect 28998 22072 29054 22108
rect 28814 21936 28870 21992
rect 28906 19916 28962 19952
rect 28906 19896 28908 19916
rect 28908 19896 28960 19916
rect 28960 19896 28962 19916
rect 28814 15136 28870 15192
rect 29182 15136 29238 15192
rect 29918 27512 29974 27568
rect 30746 33360 30802 33416
rect 31574 38276 31630 38312
rect 31574 38256 31576 38276
rect 31576 38256 31628 38276
rect 31628 38256 31630 38276
rect 31666 37168 31722 37224
rect 31114 32952 31170 33008
rect 31206 32544 31262 32600
rect 31206 30132 31208 30152
rect 31208 30132 31260 30152
rect 31260 30132 31262 30152
rect 31206 30096 31262 30132
rect 30286 28328 30342 28384
rect 29734 20576 29790 20632
rect 30654 26308 30710 26344
rect 30654 26288 30656 26308
rect 30656 26288 30708 26308
rect 30708 26288 30710 26308
rect 32402 38392 32458 38448
rect 32034 37304 32090 37360
rect 31942 36896 31998 36952
rect 31758 35808 31814 35864
rect 32034 35944 32090 36000
rect 32494 37848 32550 37904
rect 32218 34992 32274 35048
rect 33690 39344 33746 39400
rect 33230 39244 33232 39264
rect 33232 39244 33284 39264
rect 33284 39244 33286 39264
rect 33230 39208 33286 39244
rect 32954 38800 33010 38856
rect 32770 36780 32826 36816
rect 32770 36760 32772 36780
rect 32772 36760 32824 36780
rect 32824 36760 32826 36780
rect 32770 36216 32826 36272
rect 33046 37168 33102 37224
rect 32494 34720 32550 34776
rect 32494 34584 32550 34640
rect 33598 38800 33654 38856
rect 32402 32952 32458 33008
rect 32126 32272 32182 32328
rect 32034 32000 32090 32056
rect 31850 31340 31906 31376
rect 31850 31320 31852 31340
rect 31852 31320 31904 31340
rect 31904 31320 31906 31340
rect 31942 30540 31944 30560
rect 31944 30540 31996 30560
rect 31996 30540 31998 30560
rect 31942 30504 31998 30540
rect 31482 28056 31538 28112
rect 31390 21936 31446 21992
rect 32862 32952 32918 33008
rect 31850 23740 31852 23760
rect 31852 23740 31904 23760
rect 31904 23740 31906 23760
rect 31850 23704 31906 23740
rect 32034 24656 32090 24712
rect 32034 22108 32036 22128
rect 32036 22108 32088 22128
rect 32088 22108 32090 22128
rect 32034 22072 32090 22108
rect 29826 14864 29882 14920
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 31666 14184 31722 14240
rect 32310 24792 32366 24848
rect 32402 22616 32458 22672
rect 32310 22208 32366 22264
rect 32678 23724 32734 23760
rect 32678 23704 32680 23724
rect 32680 23704 32732 23724
rect 32732 23704 32734 23724
rect 33966 37868 34022 37904
rect 33966 37848 33968 37868
rect 33968 37848 34020 37868
rect 34020 37848 34022 37868
rect 33230 31884 33286 31920
rect 33230 31864 33232 31884
rect 33232 31864 33284 31884
rect 33284 31864 33286 31884
rect 33046 29008 33102 29064
rect 33322 30912 33378 30968
rect 33598 33924 33654 33960
rect 33598 33904 33600 33924
rect 33600 33904 33652 33924
rect 33652 33904 33654 33924
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34242 37168 34298 37224
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35254 38256 35310 38312
rect 35162 38120 35218 38176
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34610 37168 34666 37224
rect 34150 34312 34206 34368
rect 33782 32836 33838 32872
rect 33782 32816 33784 32836
rect 33784 32816 33836 32836
rect 33836 32816 33838 32836
rect 33690 32272 33746 32328
rect 33230 28212 33286 28248
rect 33230 28192 33232 28212
rect 33232 28192 33284 28212
rect 33284 28192 33286 28212
rect 33966 32000 34022 32056
rect 34058 31592 34114 31648
rect 33046 26016 33102 26072
rect 33322 26288 33378 26344
rect 33138 23160 33194 23216
rect 32310 16360 32366 16416
rect 32586 16088 32642 16144
rect 32494 15272 32550 15328
rect 32218 11348 32274 11384
rect 32218 11328 32220 11348
rect 32220 11328 32272 11348
rect 32272 11328 32274 11348
rect 34426 30368 34482 30424
rect 35162 36896 35218 36952
rect 35530 38956 35586 38992
rect 35530 38936 35532 38956
rect 35532 38936 35584 38956
rect 35584 38936 35586 38956
rect 35530 37868 35586 37904
rect 35530 37848 35532 37868
rect 35532 37848 35584 37868
rect 35584 37848 35586 37868
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35346 35808 35402 35864
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34886 35164 34888 35184
rect 34888 35164 34940 35184
rect 34940 35164 34942 35184
rect 34886 35128 34942 35164
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35162 32428 35218 32464
rect 35162 32408 35164 32428
rect 35164 32408 35216 32428
rect 35216 32408 35218 32428
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34610 31864 34666 31920
rect 34518 30252 34574 30288
rect 34518 30232 34520 30252
rect 34520 30232 34572 30252
rect 34572 30232 34574 30252
rect 34518 29588 34520 29608
rect 34520 29588 34572 29608
rect 34572 29588 34574 29608
rect 34518 29552 34574 29588
rect 33782 26324 33784 26344
rect 33784 26324 33836 26344
rect 33836 26324 33838 26344
rect 33782 26288 33838 26324
rect 34058 26152 34114 26208
rect 34518 27920 34574 27976
rect 34518 27512 34574 27568
rect 34334 26868 34336 26888
rect 34336 26868 34388 26888
rect 34388 26868 34390 26888
rect 34334 26832 34390 26868
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35530 36760 35586 36816
rect 36082 39888 36138 39944
rect 35898 36116 35900 36136
rect 35900 36116 35952 36136
rect 35952 36116 35954 36136
rect 35898 36080 35954 36116
rect 36174 37848 36230 37904
rect 35806 33940 35808 33960
rect 35808 33940 35860 33960
rect 35860 33940 35862 33960
rect 35806 33904 35862 33940
rect 36542 37440 36598 37496
rect 35714 32544 35770 32600
rect 35438 31048 35494 31104
rect 35346 30776 35402 30832
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35714 31320 35770 31376
rect 35622 29144 35678 29200
rect 35438 28464 35494 28520
rect 35162 28076 35218 28112
rect 35162 28056 35164 28076
rect 35164 28056 35216 28076
rect 35216 28056 35218 28076
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34426 26152 34482 26208
rect 34242 24248 34298 24304
rect 34150 23840 34206 23896
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35254 26308 35310 26344
rect 35254 26288 35256 26308
rect 35256 26288 35308 26308
rect 35308 26288 35310 26308
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 36450 34448 36506 34504
rect 36266 33088 36322 33144
rect 36082 32272 36138 32328
rect 37278 38256 37334 38312
rect 36818 36216 36874 36272
rect 36726 36116 36728 36136
rect 36728 36116 36780 36136
rect 36780 36116 36782 36136
rect 36726 36080 36782 36116
rect 36634 35808 36690 35864
rect 36818 35944 36874 36000
rect 36542 33496 36598 33552
rect 36634 32952 36690 33008
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35438 23296 35494 23352
rect 35990 27240 36046 27296
rect 35990 24792 36046 24848
rect 35346 20576 35402 20632
rect 33966 19352 34022 19408
rect 33506 15272 33562 15328
rect 33322 15036 33324 15056
rect 33324 15036 33376 15056
rect 33376 15036 33378 15056
rect 33322 15000 33378 15036
rect 33322 14184 33378 14240
rect 32862 11328 32918 11384
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34150 16496 34206 16552
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34886 16360 34942 16416
rect 35254 16532 35256 16552
rect 35256 16532 35308 16552
rect 35308 16532 35310 16552
rect 35254 16496 35310 16532
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35070 14864 35126 14920
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35070 14456 35126 14512
rect 36818 31864 36874 31920
rect 36450 31048 36506 31104
rect 36358 30096 36414 30152
rect 36450 29960 36506 30016
rect 36358 29008 36414 29064
rect 36358 27532 36414 27568
rect 36358 27512 36360 27532
rect 36360 27512 36412 27532
rect 36412 27512 36414 27532
rect 37186 35808 37242 35864
rect 37462 35980 37464 36000
rect 37464 35980 37516 36000
rect 37516 35980 37518 36000
rect 37462 35944 37518 35980
rect 38014 39380 38016 39400
rect 38016 39380 38068 39400
rect 38068 39380 38070 39400
rect 38014 39344 38070 39380
rect 37922 37168 37978 37224
rect 37830 36352 37886 36408
rect 37738 36116 37740 36136
rect 37740 36116 37792 36136
rect 37792 36116 37794 36136
rect 37738 36080 37794 36116
rect 37002 32000 37058 32056
rect 37002 31764 37004 31784
rect 37004 31764 37056 31784
rect 37056 31764 37058 31784
rect 37002 31728 37058 31764
rect 37002 31356 37004 31376
rect 37004 31356 37056 31376
rect 37056 31356 37058 31376
rect 37002 31320 37058 31356
rect 37738 34856 37794 34912
rect 37462 32680 37518 32736
rect 37370 32272 37426 32328
rect 38382 36352 38438 36408
rect 38106 35672 38162 35728
rect 38014 33632 38070 33688
rect 37922 33360 37978 33416
rect 37094 24792 37150 24848
rect 36266 23976 36322 24032
rect 36266 23568 36322 23624
rect 36542 23568 36598 23624
rect 36634 22636 36690 22672
rect 36634 22616 36636 22636
rect 36636 22616 36688 22636
rect 36688 22616 36690 22636
rect 35622 14456 35678 14512
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 36818 22636 36874 22672
rect 36818 22616 36820 22636
rect 36820 22616 36872 22636
rect 36872 22616 36874 22636
rect 36174 16124 36176 16144
rect 36176 16124 36228 16144
rect 36228 16124 36230 16144
rect 36174 16088 36230 16124
rect 35898 15036 35900 15056
rect 35900 15036 35952 15056
rect 35952 15036 35954 15056
rect 35898 15000 35954 15036
rect 35806 14864 35862 14920
rect 37094 24284 37096 24304
rect 37096 24284 37148 24304
rect 37148 24284 37150 24304
rect 37094 24248 37150 24284
rect 37462 27940 37518 27976
rect 37462 27920 37464 27940
rect 37464 27920 37516 27940
rect 37516 27920 37518 27940
rect 37094 23704 37150 23760
rect 37186 23296 37242 23352
rect 36726 15272 36782 15328
rect 37186 21972 37188 21992
rect 37188 21972 37240 21992
rect 37240 21972 37242 21992
rect 37186 21936 37242 21972
rect 37462 26152 37518 26208
rect 37370 25492 37426 25528
rect 37370 25472 37372 25492
rect 37372 25472 37424 25492
rect 37424 25472 37426 25492
rect 37554 24656 37610 24712
rect 38198 32136 38254 32192
rect 38106 31048 38162 31104
rect 39026 37712 39082 37768
rect 39302 38120 39358 38176
rect 39026 36896 39082 36952
rect 39210 35672 39266 35728
rect 39486 35536 39542 35592
rect 39210 34856 39266 34912
rect 39118 34040 39174 34096
rect 39394 33516 39450 33552
rect 39394 33496 39396 33516
rect 39396 33496 39448 33516
rect 39448 33496 39450 33516
rect 38750 32544 38806 32600
rect 38750 31864 38806 31920
rect 40222 38936 40278 38992
rect 40038 37304 40094 37360
rect 40406 38936 40462 38992
rect 40682 37304 40738 37360
rect 39762 35692 39818 35728
rect 39762 35672 39764 35692
rect 39764 35672 39816 35692
rect 39816 35672 39818 35692
rect 39670 35012 39726 35048
rect 39670 34992 39672 35012
rect 39672 34992 39724 35012
rect 39724 34992 39726 35012
rect 38474 30096 38530 30152
rect 38290 29960 38346 30016
rect 38198 27512 38254 27568
rect 37830 26968 37886 27024
rect 37922 26288 37978 26344
rect 37830 24676 37886 24712
rect 37830 24656 37832 24676
rect 37832 24656 37884 24676
rect 37884 24656 37886 24676
rect 37830 23976 37886 24032
rect 37830 23604 37832 23624
rect 37832 23604 37884 23624
rect 37884 23604 37886 23624
rect 37830 23568 37886 23604
rect 38106 26832 38162 26888
rect 38014 24248 38070 24304
rect 38014 23296 38070 23352
rect 39026 29044 39028 29064
rect 39028 29044 39080 29064
rect 39080 29044 39082 29064
rect 38474 27276 38476 27296
rect 38476 27276 38528 27296
rect 38528 27276 38530 27296
rect 38474 27240 38530 27276
rect 38290 26988 38346 27024
rect 38290 26968 38292 26988
rect 38292 26968 38344 26988
rect 38344 26968 38346 26988
rect 38382 26832 38438 26888
rect 39026 29008 39082 29044
rect 39394 30676 39396 30696
rect 39396 30676 39448 30696
rect 39448 30676 39450 30696
rect 39394 30640 39450 30676
rect 39210 29008 39266 29064
rect 39026 27396 39082 27432
rect 39026 27376 39028 27396
rect 39028 27376 39080 27396
rect 39080 27376 39082 27396
rect 38474 26152 38530 26208
rect 39210 25900 39266 25936
rect 39210 25880 39212 25900
rect 39212 25880 39264 25900
rect 39264 25880 39266 25900
rect 38934 23704 38990 23760
rect 37094 16088 37150 16144
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38198 14476 38254 14512
rect 38198 14456 38200 14476
rect 38200 14456 38252 14476
rect 38252 14456 38254 14476
rect 40222 36216 40278 36272
rect 40314 34620 40316 34640
rect 40316 34620 40368 34640
rect 40368 34620 40370 34640
rect 40314 34584 40370 34620
rect 40038 33940 40040 33960
rect 40040 33940 40092 33960
rect 40092 33940 40094 33960
rect 40038 33904 40094 33940
rect 40222 33088 40278 33144
rect 40314 31728 40370 31784
rect 40866 35808 40922 35864
rect 40866 35536 40922 35592
rect 40866 33224 40922 33280
rect 40498 31864 40554 31920
rect 40590 31728 40646 31784
rect 39394 23704 39450 23760
rect 39302 18964 39358 19000
rect 39302 18944 39304 18964
rect 39304 18944 39356 18964
rect 39356 18944 39358 18964
rect 39670 22752 39726 22808
rect 39670 22072 39726 22128
rect 39670 19388 39672 19408
rect 39672 19388 39724 19408
rect 39724 19388 39726 19408
rect 39670 19352 39726 19388
rect 40866 31728 40922 31784
rect 40314 27376 40370 27432
rect 40038 24404 40094 24440
rect 40038 24384 40040 24404
rect 40040 24384 40092 24404
rect 40092 24384 40094 24404
rect 41602 31864 41658 31920
rect 40406 24404 40462 24440
rect 40406 24384 40408 24404
rect 40408 24384 40460 24404
rect 40460 24384 40462 24404
rect 40958 24112 41014 24168
rect 41326 22072 41382 22128
rect 41786 30640 41842 30696
rect 42614 37712 42670 37768
rect 43994 42608 44050 42664
rect 43350 36624 43406 36680
rect 42890 35672 42946 35728
rect 42706 31220 42708 31240
rect 42708 31220 42760 31240
rect 42760 31220 42762 31240
rect 42706 31184 42762 31220
rect 42798 30796 42854 30832
rect 42798 30776 42800 30796
rect 42800 30776 42852 30796
rect 42852 30776 42854 30796
rect 42614 30640 42670 30696
rect 42890 30232 42946 30288
rect 41326 20712 41382 20768
rect 40774 19372 40830 19408
rect 40774 19352 40776 19372
rect 40776 19352 40828 19372
rect 40828 19352 40830 19372
rect 39946 17720 40002 17776
rect 39210 15544 39266 15600
rect 43074 25880 43130 25936
rect 43994 35264 44050 35320
rect 43994 31592 44050 31648
rect 43994 27920 44050 27976
rect 39118 12008 39174 12064
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 39670 12008 39726 12064
rect 41234 14068 41290 14104
rect 41234 14048 41236 14068
rect 41236 14048 41288 14068
rect 41288 14048 41290 14068
rect 40866 11892 40922 11928
rect 40866 11872 40868 11892
rect 40868 11872 40920 11892
rect 40920 11872 40922 11892
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 43074 14340 43130 14376
rect 43074 14320 43076 14340
rect 43076 14320 43128 14340
rect 43128 14320 43130 14340
rect 42798 13232 42854 13288
rect 43994 24248 44050 24304
rect 43994 20576 44050 20632
rect 43350 13232 43406 13288
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 43994 16904 44050 16960
rect 43994 9560 44050 9616
rect 43350 5908 43406 5944
rect 43350 5888 43352 5908
rect 43352 5888 43404 5908
rect 43404 5888 43406 5908
rect 43994 2216 44050 2272
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 43989 42666 44055 42669
rect 44200 42666 45000 42756
rect 43989 42664 45000 42666
rect 43989 42608 43994 42664
rect 44050 42608 45000 42664
rect 43989 42606 45000 42608
rect 43989 42603 44055 42606
rect 44200 42516 45000 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 27889 39946 27955 39949
rect 28758 39946 28764 39948
rect 27889 39944 28764 39946
rect 27889 39888 27894 39944
rect 27950 39888 28764 39944
rect 27889 39886 28764 39888
rect 27889 39883 27955 39886
rect 28758 39884 28764 39886
rect 28828 39884 28834 39948
rect 31477 39946 31543 39949
rect 36077 39946 36143 39949
rect 31477 39944 36143 39946
rect 31477 39888 31482 39944
rect 31538 39888 36082 39944
rect 36138 39888 36143 39944
rect 31477 39886 36143 39888
rect 31477 39883 31543 39886
rect 36077 39883 36143 39886
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 33685 39402 33751 39405
rect 38009 39402 38075 39405
rect 33685 39400 38075 39402
rect 33685 39344 33690 39400
rect 33746 39344 38014 39400
rect 38070 39344 38075 39400
rect 33685 39342 38075 39344
rect 33685 39339 33751 39342
rect 38009 39339 38075 39342
rect 33225 39268 33291 39269
rect 33174 39204 33180 39268
rect 33244 39266 33291 39268
rect 33244 39264 33336 39266
rect 33286 39208 33336 39264
rect 33244 39206 33336 39208
rect 33244 39204 33291 39206
rect 33225 39203 33291 39204
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 27521 38996 27587 38997
rect 27470 38932 27476 38996
rect 27540 38994 27587 38996
rect 30373 38994 30439 38997
rect 35525 38994 35591 38997
rect 40217 38994 40283 38997
rect 40401 38994 40467 38997
rect 27540 38992 27632 38994
rect 27582 38936 27632 38992
rect 27540 38934 27632 38936
rect 30373 38992 40467 38994
rect 30373 38936 30378 38992
rect 30434 38936 35530 38992
rect 35586 38936 40222 38992
rect 40278 38936 40406 38992
rect 40462 38936 40467 38992
rect 30373 38934 40467 38936
rect 27540 38932 27587 38934
rect 27521 38931 27587 38932
rect 30373 38931 30439 38934
rect 35525 38931 35591 38934
rect 40217 38931 40283 38934
rect 40401 38931 40467 38934
rect 40534 38932 40540 38996
rect 40604 38994 40610 38996
rect 44200 38994 45000 39084
rect 40604 38934 45000 38994
rect 40604 38932 40610 38934
rect 16941 38858 17007 38861
rect 28993 38858 29059 38861
rect 16941 38856 29059 38858
rect 16941 38800 16946 38856
rect 17002 38800 28998 38856
rect 29054 38800 29059 38856
rect 16941 38798 29059 38800
rect 16941 38795 17007 38798
rect 28993 38795 29059 38798
rect 32949 38858 33015 38861
rect 33593 38858 33659 38861
rect 32949 38856 33659 38858
rect 32949 38800 32954 38856
rect 33010 38800 33598 38856
rect 33654 38800 33659 38856
rect 44200 38844 45000 38934
rect 32949 38798 33659 38800
rect 32949 38795 33015 38798
rect 33593 38795 33659 38798
rect 28758 38660 28764 38724
rect 28828 38722 28834 38724
rect 28901 38722 28967 38725
rect 28828 38720 28967 38722
rect 28828 38664 28906 38720
rect 28962 38664 28967 38720
rect 28828 38662 28967 38664
rect 28828 38660 28834 38662
rect 28901 38659 28967 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 17217 38450 17283 38453
rect 25497 38450 25563 38453
rect 26141 38450 26207 38453
rect 17217 38448 26207 38450
rect 17217 38392 17222 38448
rect 17278 38392 25502 38448
rect 25558 38392 26146 38448
rect 26202 38392 26207 38448
rect 17217 38390 26207 38392
rect 17217 38387 17283 38390
rect 25497 38387 25563 38390
rect 26141 38387 26207 38390
rect 28349 38450 28415 38453
rect 28574 38450 28580 38452
rect 28349 38448 28580 38450
rect 28349 38392 28354 38448
rect 28410 38392 28580 38448
rect 28349 38390 28580 38392
rect 28349 38387 28415 38390
rect 28574 38388 28580 38390
rect 28644 38450 28650 38452
rect 32397 38450 32463 38453
rect 28644 38448 32463 38450
rect 28644 38392 32402 38448
rect 32458 38392 32463 38448
rect 28644 38390 32463 38392
rect 28644 38388 28650 38390
rect 32397 38387 32463 38390
rect 21541 38314 21607 38317
rect 23565 38314 23631 38317
rect 21541 38312 23631 38314
rect 21541 38256 21546 38312
rect 21602 38256 23570 38312
rect 23626 38256 23631 38312
rect 21541 38254 23631 38256
rect 21541 38251 21607 38254
rect 23565 38251 23631 38254
rect 24761 38314 24827 38317
rect 26233 38314 26299 38317
rect 28625 38314 28691 38317
rect 24761 38312 28691 38314
rect 24761 38256 24766 38312
rect 24822 38256 26238 38312
rect 26294 38256 28630 38312
rect 28686 38256 28691 38312
rect 24761 38254 28691 38256
rect 24761 38251 24827 38254
rect 26233 38251 26299 38254
rect 28625 38251 28691 38254
rect 28901 38314 28967 38317
rect 31569 38314 31635 38317
rect 35249 38314 35315 38317
rect 37273 38314 37339 38317
rect 28901 38312 37339 38314
rect 28901 38256 28906 38312
rect 28962 38256 31574 38312
rect 31630 38256 35254 38312
rect 35310 38256 37278 38312
rect 37334 38256 37339 38312
rect 28901 38254 37339 38256
rect 28901 38251 28967 38254
rect 31569 38251 31635 38254
rect 35249 38251 35315 38254
rect 37273 38251 37339 38254
rect 24301 38178 24367 38181
rect 24894 38178 24900 38180
rect 24301 38176 24900 38178
rect 24301 38120 24306 38176
rect 24362 38120 24900 38176
rect 24301 38118 24900 38120
rect 24301 38115 24367 38118
rect 24894 38116 24900 38118
rect 24964 38178 24970 38180
rect 25681 38178 25747 38181
rect 24964 38176 25747 38178
rect 24964 38120 25686 38176
rect 25742 38120 25747 38176
rect 24964 38118 25747 38120
rect 24964 38116 24970 38118
rect 25681 38115 25747 38118
rect 35157 38178 35223 38181
rect 35382 38178 35388 38180
rect 35157 38176 35388 38178
rect 35157 38120 35162 38176
rect 35218 38120 35388 38176
rect 35157 38118 35388 38120
rect 35157 38115 35223 38118
rect 35382 38116 35388 38118
rect 35452 38178 35458 38180
rect 39297 38178 39363 38181
rect 35452 38176 39363 38178
rect 35452 38120 39302 38176
rect 39358 38120 39363 38176
rect 35452 38118 39363 38120
rect 35452 38116 35458 38118
rect 39297 38115 39363 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 21449 38042 21515 38045
rect 22921 38042 22987 38045
rect 21449 38040 22987 38042
rect 21449 37984 21454 38040
rect 21510 37984 22926 38040
rect 22982 37984 22987 38040
rect 21449 37982 22987 37984
rect 21449 37979 21515 37982
rect 22921 37979 22987 37982
rect 25865 38042 25931 38045
rect 26969 38042 27035 38045
rect 25865 38040 27035 38042
rect 25865 37984 25870 38040
rect 25926 37984 26974 38040
rect 27030 37984 27035 38040
rect 25865 37982 27035 37984
rect 25865 37979 25931 37982
rect 26969 37979 27035 37982
rect 28717 38042 28783 38045
rect 28993 38042 29059 38045
rect 28717 38040 39084 38042
rect 28717 37984 28722 38040
rect 28778 37984 28998 38040
rect 29054 37984 39084 38040
rect 28717 37982 39084 37984
rect 28717 37979 28783 37982
rect 28993 37979 29059 37982
rect 15193 37906 15259 37909
rect 22553 37906 22619 37909
rect 23013 37906 23079 37909
rect 28257 37906 28323 37909
rect 29361 37906 29427 37909
rect 15193 37904 23079 37906
rect 15193 37848 15198 37904
rect 15254 37848 22558 37904
rect 22614 37848 23018 37904
rect 23074 37848 23079 37904
rect 15193 37846 23079 37848
rect 15193 37843 15259 37846
rect 22553 37843 22619 37846
rect 23013 37843 23079 37846
rect 25086 37904 29427 37906
rect 25086 37848 28262 37904
rect 28318 37848 29366 37904
rect 29422 37848 29427 37904
rect 25086 37846 29427 37848
rect 15561 37634 15627 37637
rect 25086 37634 25146 37846
rect 28257 37843 28323 37846
rect 29361 37843 29427 37846
rect 32489 37906 32555 37909
rect 33961 37906 34027 37909
rect 32489 37904 34027 37906
rect 32489 37848 32494 37904
rect 32550 37848 33966 37904
rect 34022 37848 34027 37904
rect 32489 37846 34027 37848
rect 32489 37843 32555 37846
rect 33961 37843 34027 37846
rect 35525 37906 35591 37909
rect 36169 37906 36235 37909
rect 35525 37904 36235 37906
rect 35525 37848 35530 37904
rect 35586 37848 36174 37904
rect 36230 37848 36235 37904
rect 35525 37846 36235 37848
rect 35525 37843 35591 37846
rect 36169 37843 36235 37846
rect 39024 37773 39084 37982
rect 25221 37770 25287 37773
rect 36302 37770 36308 37772
rect 25221 37768 36308 37770
rect 25221 37712 25226 37768
rect 25282 37712 36308 37768
rect 25221 37710 36308 37712
rect 25221 37707 25287 37710
rect 36302 37708 36308 37710
rect 36372 37708 36378 37772
rect 39021 37770 39087 37773
rect 42609 37770 42675 37773
rect 39021 37768 42675 37770
rect 39021 37712 39026 37768
rect 39082 37712 42614 37768
rect 42670 37712 42675 37768
rect 39021 37710 42675 37712
rect 39021 37707 39087 37710
rect 15561 37632 25146 37634
rect 15561 37576 15566 37632
rect 15622 37576 25146 37632
rect 15561 37574 25146 37576
rect 15561 37571 15627 37574
rect 27286 37572 27292 37636
rect 27356 37634 27362 37636
rect 27429 37634 27495 37637
rect 27356 37632 27495 37634
rect 27356 37576 27434 37632
rect 27490 37576 27495 37632
rect 27356 37574 27495 37576
rect 27356 37572 27362 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 16665 37498 16731 37501
rect 27294 37498 27354 37572
rect 27429 37571 27495 37574
rect 29729 37634 29795 37637
rect 29862 37634 29868 37636
rect 29729 37632 29868 37634
rect 29729 37576 29734 37632
rect 29790 37576 29868 37632
rect 29729 37574 29868 37576
rect 29729 37571 29795 37574
rect 29862 37572 29868 37574
rect 29932 37572 29938 37636
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 16665 37496 27354 37498
rect 16665 37440 16670 37496
rect 16726 37440 27354 37496
rect 16665 37438 27354 37440
rect 36537 37498 36603 37501
rect 37222 37498 37228 37500
rect 36537 37496 37228 37498
rect 36537 37440 36542 37496
rect 36598 37440 37228 37496
rect 36537 37438 37228 37440
rect 16665 37435 16731 37438
rect 36537 37435 36603 37438
rect 37222 37436 37228 37438
rect 37292 37436 37298 37500
rect 40726 37365 40786 37710
rect 42609 37707 42675 37710
rect 24761 37362 24827 37365
rect 25078 37362 25084 37364
rect 24761 37360 25084 37362
rect 24761 37304 24766 37360
rect 24822 37304 25084 37360
rect 24761 37302 25084 37304
rect 24761 37299 24827 37302
rect 25078 37300 25084 37302
rect 25148 37362 25154 37364
rect 25313 37362 25379 37365
rect 25148 37360 25379 37362
rect 25148 37304 25318 37360
rect 25374 37304 25379 37360
rect 25148 37302 25379 37304
rect 25148 37300 25154 37302
rect 25313 37299 25379 37302
rect 29269 37362 29335 37365
rect 30281 37362 30347 37365
rect 32029 37362 32095 37365
rect 40033 37362 40099 37365
rect 29269 37360 29746 37362
rect 29269 37304 29274 37360
rect 29330 37304 29746 37360
rect 29269 37302 29746 37304
rect 29269 37299 29335 37302
rect 23565 37090 23631 37093
rect 25865 37090 25931 37093
rect 23565 37088 25931 37090
rect 23565 37032 23570 37088
rect 23626 37032 25870 37088
rect 25926 37032 25931 37088
rect 23565 37030 25931 37032
rect 29686 37090 29746 37302
rect 30281 37360 32095 37362
rect 30281 37304 30286 37360
rect 30342 37304 32034 37360
rect 32090 37304 32095 37360
rect 30281 37302 32095 37304
rect 30281 37299 30347 37302
rect 32029 37299 32095 37302
rect 34470 37360 40099 37362
rect 34470 37304 40038 37360
rect 40094 37304 40099 37360
rect 34470 37302 40099 37304
rect 29913 37226 29979 37229
rect 31661 37226 31727 37229
rect 33041 37226 33107 37229
rect 29913 37224 33107 37226
rect 29913 37168 29918 37224
rect 29974 37168 31666 37224
rect 31722 37168 33046 37224
rect 33102 37168 33107 37224
rect 29913 37166 33107 37168
rect 29913 37163 29979 37166
rect 31661 37163 31727 37166
rect 33041 37163 33107 37166
rect 34237 37226 34303 37229
rect 34470 37226 34530 37302
rect 40033 37299 40099 37302
rect 40677 37360 40786 37365
rect 40677 37304 40682 37360
rect 40738 37304 40786 37360
rect 40677 37302 40786 37304
rect 40677 37299 40743 37302
rect 34237 37224 34530 37226
rect 34237 37168 34242 37224
rect 34298 37168 34530 37224
rect 34237 37166 34530 37168
rect 34605 37226 34671 37229
rect 37917 37226 37983 37229
rect 34605 37224 37983 37226
rect 34605 37168 34610 37224
rect 34666 37168 37922 37224
rect 37978 37168 37983 37224
rect 34605 37166 37983 37168
rect 34237 37163 34303 37166
rect 34605 37163 34671 37166
rect 37917 37163 37983 37166
rect 30005 37090 30071 37093
rect 29686 37088 30071 37090
rect 29686 37032 30010 37088
rect 30066 37032 30071 37088
rect 29686 37030 30071 37032
rect 23565 37027 23631 37030
rect 25865 37027 25931 37030
rect 30005 37027 30071 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 22277 36954 22343 36957
rect 24761 36954 24827 36957
rect 22277 36952 24827 36954
rect 22277 36896 22282 36952
rect 22338 36896 24766 36952
rect 24822 36896 24827 36952
rect 22277 36894 24827 36896
rect 22277 36891 22343 36894
rect 24761 36891 24827 36894
rect 31937 36954 32003 36957
rect 33174 36954 33180 36956
rect 31937 36952 33180 36954
rect 31937 36896 31942 36952
rect 31998 36896 33180 36952
rect 31937 36894 33180 36896
rect 31937 36891 32003 36894
rect 33174 36892 33180 36894
rect 33244 36954 33250 36956
rect 35157 36954 35223 36957
rect 39021 36954 39087 36957
rect 33244 36952 39087 36954
rect 33244 36896 35162 36952
rect 35218 36896 39026 36952
rect 39082 36896 39087 36952
rect 33244 36894 39087 36896
rect 33244 36892 33250 36894
rect 35157 36891 35223 36894
rect 39021 36891 39087 36894
rect 25497 36818 25563 36821
rect 25865 36818 25931 36821
rect 26969 36818 27035 36821
rect 25497 36816 27035 36818
rect 25497 36760 25502 36816
rect 25558 36760 25870 36816
rect 25926 36760 26974 36816
rect 27030 36760 27035 36816
rect 25497 36758 27035 36760
rect 25497 36755 25563 36758
rect 25865 36755 25931 36758
rect 26969 36755 27035 36758
rect 32765 36818 32831 36821
rect 35525 36818 35591 36821
rect 32765 36816 35591 36818
rect 32765 36760 32770 36816
rect 32826 36760 35530 36816
rect 35586 36760 35591 36816
rect 32765 36758 35591 36760
rect 32765 36755 32831 36758
rect 35525 36755 35591 36758
rect 14089 36682 14155 36685
rect 43345 36682 43411 36685
rect 14089 36680 43411 36682
rect 14089 36624 14094 36680
rect 14150 36624 43350 36680
rect 43406 36624 43411 36680
rect 14089 36622 43411 36624
rect 14089 36619 14155 36622
rect 43345 36619 43411 36622
rect 23197 36546 23263 36549
rect 26509 36546 26575 36549
rect 23197 36544 26575 36546
rect 23197 36488 23202 36544
rect 23258 36488 26514 36544
rect 26570 36488 26575 36544
rect 23197 36486 26575 36488
rect 23197 36483 23263 36486
rect 26509 36483 26575 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 22277 36410 22343 36413
rect 23749 36410 23815 36413
rect 22277 36408 23815 36410
rect 22277 36352 22282 36408
rect 22338 36352 23754 36408
rect 23810 36352 23815 36408
rect 22277 36350 23815 36352
rect 22277 36347 22343 36350
rect 23749 36347 23815 36350
rect 24117 36410 24183 36413
rect 26417 36410 26483 36413
rect 37825 36410 37891 36413
rect 38377 36410 38443 36413
rect 24117 36408 26483 36410
rect 24117 36352 24122 36408
rect 24178 36352 26422 36408
rect 26478 36352 26483 36408
rect 24117 36350 26483 36352
rect 24117 36347 24183 36350
rect 26417 36347 26483 36350
rect 36862 36408 38443 36410
rect 36862 36352 37830 36408
rect 37886 36352 38382 36408
rect 38438 36352 38443 36408
rect 36862 36350 38443 36352
rect 36862 36277 36922 36350
rect 37825 36347 37891 36350
rect 38377 36347 38443 36350
rect 23289 36274 23355 36277
rect 25814 36274 25820 36276
rect 23289 36272 25820 36274
rect 23289 36216 23294 36272
rect 23350 36216 25820 36272
rect 23289 36214 25820 36216
rect 23289 36211 23355 36214
rect 25814 36212 25820 36214
rect 25884 36274 25890 36276
rect 32765 36274 32831 36277
rect 25884 36272 32831 36274
rect 25884 36216 32770 36272
rect 32826 36216 32831 36272
rect 25884 36214 32831 36216
rect 25884 36212 25890 36214
rect 32765 36211 32831 36214
rect 36813 36272 36922 36277
rect 36813 36216 36818 36272
rect 36874 36216 36922 36272
rect 36813 36214 36922 36216
rect 36813 36211 36879 36214
rect 37222 36212 37228 36276
rect 37292 36274 37298 36276
rect 40217 36274 40283 36277
rect 37292 36272 40283 36274
rect 37292 36216 40222 36272
rect 40278 36216 40283 36272
rect 37292 36214 40283 36216
rect 37292 36212 37298 36214
rect 40217 36211 40283 36214
rect 24577 36138 24643 36141
rect 24894 36138 24900 36140
rect 24577 36136 24900 36138
rect 24577 36080 24582 36136
rect 24638 36080 24900 36136
rect 24577 36078 24900 36080
rect 24577 36075 24643 36078
rect 24894 36076 24900 36078
rect 24964 36076 24970 36140
rect 25313 36138 25379 36141
rect 27705 36138 27771 36141
rect 25313 36136 27771 36138
rect 25313 36080 25318 36136
rect 25374 36080 27710 36136
rect 27766 36080 27771 36136
rect 25313 36078 27771 36080
rect 25313 36075 25379 36078
rect 27705 36075 27771 36078
rect 30281 36138 30347 36141
rect 35893 36138 35959 36141
rect 30281 36136 35959 36138
rect 30281 36080 30286 36136
rect 30342 36080 35898 36136
rect 35954 36080 35959 36136
rect 30281 36078 35959 36080
rect 30281 36075 30347 36078
rect 35893 36075 35959 36078
rect 36721 36138 36787 36141
rect 37733 36138 37799 36141
rect 36721 36136 37799 36138
rect 36721 36080 36726 36136
rect 36782 36080 37738 36136
rect 37794 36080 37799 36136
rect 36721 36078 37799 36080
rect 36721 36075 36787 36078
rect 37733 36075 37799 36078
rect 23933 36002 23999 36005
rect 25497 36002 25563 36005
rect 27613 36002 27679 36005
rect 23933 36000 27679 36002
rect 23933 35944 23938 36000
rect 23994 35944 25502 36000
rect 25558 35944 27618 36000
rect 27674 35944 27679 36000
rect 23933 35942 27679 35944
rect 23933 35939 23999 35942
rect 25497 35939 25563 35942
rect 27613 35939 27679 35942
rect 32029 36002 32095 36005
rect 36813 36002 36879 36005
rect 37457 36002 37523 36005
rect 32029 36000 36879 36002
rect 32029 35944 32034 36000
rect 32090 35944 36818 36000
rect 36874 35944 36879 36000
rect 32029 35942 36879 35944
rect 32029 35939 32095 35942
rect 36813 35939 36879 35942
rect 37046 36000 37523 36002
rect 37046 35944 37462 36000
rect 37518 35944 37523 36000
rect 37046 35942 37523 35944
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 22001 35866 22067 35869
rect 24577 35866 24643 35869
rect 25773 35866 25839 35869
rect 22001 35864 25839 35866
rect 22001 35808 22006 35864
rect 22062 35808 24582 35864
rect 24638 35808 25778 35864
rect 25834 35808 25839 35864
rect 22001 35806 25839 35808
rect 22001 35803 22067 35806
rect 24577 35803 24643 35806
rect 25773 35803 25839 35806
rect 28625 35866 28691 35869
rect 29361 35866 29427 35869
rect 28625 35864 29427 35866
rect 28625 35808 28630 35864
rect 28686 35808 29366 35864
rect 29422 35808 29427 35864
rect 28625 35806 29427 35808
rect 28625 35803 28691 35806
rect 29361 35803 29427 35806
rect 30649 35866 30715 35869
rect 31753 35866 31819 35869
rect 35341 35866 35407 35869
rect 30649 35864 35407 35866
rect 30649 35808 30654 35864
rect 30710 35808 31758 35864
rect 31814 35808 35346 35864
rect 35402 35808 35407 35864
rect 30649 35806 35407 35808
rect 30649 35803 30715 35806
rect 31753 35803 31819 35806
rect 35341 35803 35407 35806
rect 36629 35866 36695 35869
rect 37046 35866 37106 35942
rect 37457 35939 37523 35942
rect 36629 35864 37106 35866
rect 36629 35808 36634 35864
rect 36690 35808 37106 35864
rect 36629 35806 37106 35808
rect 37181 35866 37247 35869
rect 40861 35866 40927 35869
rect 37181 35864 40927 35866
rect 37181 35808 37186 35864
rect 37242 35808 40866 35864
rect 40922 35808 40927 35864
rect 37181 35806 40927 35808
rect 36629 35803 36695 35806
rect 37181 35803 37247 35806
rect 40861 35803 40927 35806
rect 24025 35730 24091 35733
rect 27337 35730 27403 35733
rect 24025 35728 27403 35730
rect 24025 35672 24030 35728
rect 24086 35672 27342 35728
rect 27398 35672 27403 35728
rect 24025 35670 27403 35672
rect 24025 35667 24091 35670
rect 27337 35667 27403 35670
rect 30189 35730 30255 35733
rect 38101 35730 38167 35733
rect 30189 35728 38167 35730
rect 30189 35672 30194 35728
rect 30250 35672 38106 35728
rect 38162 35672 38167 35728
rect 30189 35670 38167 35672
rect 30189 35667 30255 35670
rect 38101 35667 38167 35670
rect 39205 35730 39271 35733
rect 39757 35730 39823 35733
rect 42885 35730 42951 35733
rect 39205 35728 42951 35730
rect 39205 35672 39210 35728
rect 39266 35672 39762 35728
rect 39818 35672 42890 35728
rect 42946 35672 42951 35728
rect 39205 35670 42951 35672
rect 39205 35667 39271 35670
rect 39757 35667 39823 35670
rect 42885 35667 42951 35670
rect 27521 35596 27587 35597
rect 27470 35594 27476 35596
rect 27430 35534 27476 35594
rect 27540 35592 27587 35596
rect 27582 35536 27587 35592
rect 27470 35532 27476 35534
rect 27540 35532 27587 35536
rect 27521 35531 27587 35532
rect 30005 35594 30071 35597
rect 30281 35594 30347 35597
rect 39481 35594 39547 35597
rect 40861 35596 40927 35597
rect 40861 35594 40908 35596
rect 30005 35592 30114 35594
rect 30005 35536 30010 35592
rect 30066 35536 30114 35592
rect 30005 35531 30114 35536
rect 30281 35592 39547 35594
rect 30281 35536 30286 35592
rect 30342 35536 39486 35592
rect 39542 35536 39547 35592
rect 30281 35534 39547 35536
rect 40816 35592 40908 35594
rect 40816 35536 40866 35592
rect 40816 35534 40908 35536
rect 30281 35531 30347 35534
rect 39481 35531 39547 35534
rect 40861 35532 40908 35534
rect 40972 35532 40978 35596
rect 40861 35531 40927 35532
rect 27153 35458 27219 35461
rect 30054 35458 30114 35531
rect 32070 35458 32076 35460
rect 27153 35456 32076 35458
rect 27153 35400 27158 35456
rect 27214 35400 32076 35456
rect 27153 35398 32076 35400
rect 27153 35395 27219 35398
rect 32070 35396 32076 35398
rect 32140 35396 32146 35460
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 22093 35322 22159 35325
rect 25037 35322 25103 35325
rect 22093 35320 25103 35322
rect 22093 35264 22098 35320
rect 22154 35264 25042 35320
rect 25098 35264 25103 35320
rect 22093 35262 25103 35264
rect 22093 35259 22159 35262
rect 25037 35259 25103 35262
rect 43989 35322 44055 35325
rect 44200 35322 45000 35412
rect 43989 35320 45000 35322
rect 43989 35264 43994 35320
rect 44050 35264 45000 35320
rect 43989 35262 45000 35264
rect 43989 35259 44055 35262
rect 24669 35186 24735 35189
rect 34881 35186 34947 35189
rect 24669 35184 34947 35186
rect 24669 35128 24674 35184
rect 24730 35128 34886 35184
rect 34942 35128 34947 35184
rect 44200 35172 45000 35262
rect 24669 35126 34947 35128
rect 24669 35123 24735 35126
rect 34881 35123 34947 35126
rect 12249 35050 12315 35053
rect 27337 35050 27403 35053
rect 12249 35048 27403 35050
rect 12249 34992 12254 35048
rect 12310 34992 27342 35048
rect 27398 34992 27403 35048
rect 12249 34990 27403 34992
rect 12249 34987 12315 34990
rect 27337 34987 27403 34990
rect 28349 35050 28415 35053
rect 28758 35050 28764 35052
rect 28349 35048 28764 35050
rect 28349 34992 28354 35048
rect 28410 34992 28764 35048
rect 28349 34990 28764 34992
rect 28349 34987 28415 34990
rect 28758 34988 28764 34990
rect 28828 35050 28834 35052
rect 28993 35050 29059 35053
rect 28828 35048 29059 35050
rect 28828 34992 28998 35048
rect 29054 34992 29059 35048
rect 28828 34990 29059 34992
rect 28828 34988 28834 34990
rect 28993 34987 29059 34990
rect 32213 35050 32279 35053
rect 39665 35050 39731 35053
rect 32213 35048 39731 35050
rect 32213 34992 32218 35048
rect 32274 34992 39670 35048
rect 39726 34992 39731 35048
rect 32213 34990 39731 34992
rect 32213 34987 32279 34990
rect 39665 34987 39731 34990
rect 19977 34914 20043 34917
rect 28625 34914 28691 34917
rect 19977 34912 28691 34914
rect 19977 34856 19982 34912
rect 20038 34856 28630 34912
rect 28686 34856 28691 34912
rect 19977 34854 28691 34856
rect 19977 34851 20043 34854
rect 28625 34851 28691 34854
rect 32070 34852 32076 34916
rect 32140 34914 32146 34916
rect 37733 34914 37799 34917
rect 39205 34914 39271 34917
rect 32140 34912 39271 34914
rect 32140 34856 37738 34912
rect 37794 34856 39210 34912
rect 39266 34856 39271 34912
rect 32140 34854 39271 34856
rect 32140 34852 32146 34854
rect 37733 34851 37799 34854
rect 39205 34851 39271 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 25589 34778 25655 34781
rect 32489 34778 32555 34781
rect 25589 34776 32555 34778
rect 25589 34720 25594 34776
rect 25650 34720 32494 34776
rect 32550 34720 32555 34776
rect 25589 34718 32555 34720
rect 25589 34715 25655 34718
rect 32489 34715 32555 34718
rect 10409 34642 10475 34645
rect 28993 34642 29059 34645
rect 10409 34640 29059 34642
rect 10409 34584 10414 34640
rect 10470 34584 28998 34640
rect 29054 34584 29059 34640
rect 10409 34582 29059 34584
rect 10409 34579 10475 34582
rect 28993 34579 29059 34582
rect 29913 34642 29979 34645
rect 32489 34642 32555 34645
rect 29913 34640 32555 34642
rect 29913 34584 29918 34640
rect 29974 34584 32494 34640
rect 32550 34584 32555 34640
rect 29913 34582 32555 34584
rect 29913 34579 29979 34582
rect 32489 34579 32555 34582
rect 34094 34580 34100 34644
rect 34164 34642 34170 34644
rect 40309 34642 40375 34645
rect 34164 34640 40375 34642
rect 34164 34584 40314 34640
rect 40370 34584 40375 34640
rect 34164 34582 40375 34584
rect 34164 34580 34170 34582
rect 40309 34579 40375 34582
rect 7557 34506 7623 34509
rect 20529 34506 20595 34509
rect 27337 34508 27403 34509
rect 27286 34506 27292 34508
rect 7557 34504 20595 34506
rect 7557 34448 7562 34504
rect 7618 34448 20534 34504
rect 20590 34448 20595 34504
rect 7557 34446 20595 34448
rect 27246 34446 27292 34506
rect 27356 34504 27403 34508
rect 27398 34448 27403 34504
rect 7557 34443 7623 34446
rect 20529 34443 20595 34446
rect 27286 34444 27292 34446
rect 27356 34444 27403 34448
rect 36302 34444 36308 34508
rect 36372 34506 36378 34508
rect 36445 34506 36511 34509
rect 36372 34504 36511 34506
rect 36372 34448 36450 34504
rect 36506 34448 36511 34504
rect 36372 34446 36511 34448
rect 36372 34444 36378 34446
rect 27337 34443 27403 34444
rect 36445 34443 36511 34446
rect 25221 34370 25287 34373
rect 30557 34370 30623 34373
rect 34145 34370 34211 34373
rect 25221 34368 34211 34370
rect 25221 34312 25226 34368
rect 25282 34312 30562 34368
rect 30618 34312 34150 34368
rect 34206 34312 34211 34368
rect 25221 34310 34211 34312
rect 25221 34307 25287 34310
rect 30557 34307 30623 34310
rect 34145 34307 34211 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 27981 34234 28047 34237
rect 28574 34234 28580 34236
rect 27981 34232 28580 34234
rect 27981 34176 27986 34232
rect 28042 34176 28580 34232
rect 27981 34174 28580 34176
rect 27981 34171 28047 34174
rect 28574 34172 28580 34174
rect 28644 34234 28650 34236
rect 28809 34234 28875 34237
rect 28644 34232 28875 34234
rect 28644 34176 28814 34232
rect 28870 34176 28875 34232
rect 28644 34174 28875 34176
rect 28644 34172 28650 34174
rect 28809 34171 28875 34174
rect 20805 34098 20871 34101
rect 21449 34098 21515 34101
rect 39113 34098 39179 34101
rect 20805 34096 39179 34098
rect 20805 34040 20810 34096
rect 20866 34040 21454 34096
rect 21510 34040 39118 34096
rect 39174 34040 39179 34096
rect 20805 34038 39179 34040
rect 20805 34035 20871 34038
rect 21449 34035 21515 34038
rect 39113 34035 39179 34038
rect 10685 33962 10751 33965
rect 26417 33962 26483 33965
rect 10685 33960 26483 33962
rect 10685 33904 10690 33960
rect 10746 33904 26422 33960
rect 26478 33904 26483 33960
rect 10685 33902 26483 33904
rect 10685 33899 10751 33902
rect 26417 33899 26483 33902
rect 29453 33962 29519 33965
rect 33593 33962 33659 33965
rect 29453 33960 33659 33962
rect 29453 33904 29458 33960
rect 29514 33904 33598 33960
rect 33654 33904 33659 33960
rect 29453 33902 33659 33904
rect 29453 33899 29519 33902
rect 33593 33899 33659 33902
rect 35801 33962 35867 33965
rect 40033 33962 40099 33965
rect 35801 33960 40099 33962
rect 35801 33904 35806 33960
rect 35862 33904 40038 33960
rect 40094 33904 40099 33960
rect 35801 33902 40099 33904
rect 35801 33899 35867 33902
rect 40033 33899 40099 33902
rect 25221 33828 25287 33829
rect 25221 33824 25268 33828
rect 25332 33826 25338 33828
rect 26325 33826 26391 33829
rect 25221 33768 25226 33824
rect 25221 33764 25268 33768
rect 25332 33766 25378 33826
rect 26325 33824 31770 33826
rect 26325 33768 26330 33824
rect 26386 33768 31770 33824
rect 26325 33766 31770 33768
rect 25332 33764 25338 33766
rect 25221 33763 25287 33764
rect 26325 33763 26391 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 26049 33690 26115 33693
rect 30465 33690 30531 33693
rect 26049 33688 30531 33690
rect 26049 33632 26054 33688
rect 26110 33632 30470 33688
rect 30526 33632 30531 33688
rect 26049 33630 30531 33632
rect 31710 33690 31770 33766
rect 37222 33690 37228 33692
rect 31710 33630 37228 33690
rect 26049 33627 26115 33630
rect 30465 33627 30531 33630
rect 37222 33628 37228 33630
rect 37292 33690 37298 33692
rect 38009 33690 38075 33693
rect 37292 33688 38075 33690
rect 37292 33632 38014 33688
rect 38070 33632 38075 33688
rect 37292 33630 38075 33632
rect 37292 33628 37298 33630
rect 38009 33627 38075 33630
rect 19425 33554 19491 33557
rect 20253 33554 20319 33557
rect 19425 33552 20319 33554
rect 19425 33496 19430 33552
rect 19486 33496 20258 33552
rect 20314 33496 20319 33552
rect 19425 33494 20319 33496
rect 19425 33491 19491 33494
rect 20253 33491 20319 33494
rect 28993 33554 29059 33557
rect 36537 33554 36603 33557
rect 39389 33556 39455 33557
rect 39389 33554 39436 33556
rect 28993 33552 39436 33554
rect 39500 33554 39506 33556
rect 28993 33496 28998 33552
rect 29054 33496 36542 33552
rect 36598 33496 39394 33552
rect 28993 33494 39436 33496
rect 28993 33491 29059 33494
rect 36537 33491 36603 33494
rect 39389 33492 39436 33494
rect 39500 33494 39582 33554
rect 39500 33492 39506 33494
rect 39389 33491 39455 33492
rect 26182 33356 26188 33420
rect 26252 33418 26258 33420
rect 27521 33418 27587 33421
rect 26252 33416 27587 33418
rect 26252 33360 27526 33416
rect 27582 33360 27587 33416
rect 26252 33358 27587 33360
rect 26252 33356 26258 33358
rect 27521 33355 27587 33358
rect 30741 33418 30807 33421
rect 37917 33418 37983 33421
rect 30741 33416 37983 33418
rect 30741 33360 30746 33416
rect 30802 33360 37922 33416
rect 37978 33360 37983 33416
rect 30741 33358 37983 33360
rect 30741 33355 30807 33358
rect 37917 33355 37983 33358
rect 40350 33220 40356 33284
rect 40420 33282 40426 33284
rect 40861 33282 40927 33285
rect 40420 33280 40927 33282
rect 40420 33224 40866 33280
rect 40922 33224 40927 33280
rect 40420 33222 40927 33224
rect 40420 33220 40426 33222
rect 40861 33219 40927 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 23565 33146 23631 33149
rect 30373 33146 30439 33149
rect 23565 33144 30439 33146
rect 23565 33088 23570 33144
rect 23626 33088 30378 33144
rect 30434 33088 30439 33144
rect 23565 33086 30439 33088
rect 23565 33083 23631 33086
rect 30373 33083 30439 33086
rect 36261 33146 36327 33149
rect 40217 33146 40283 33149
rect 36261 33144 40283 33146
rect 36261 33088 36266 33144
rect 36322 33088 40222 33144
rect 40278 33088 40283 33144
rect 36261 33086 40283 33088
rect 36261 33083 36327 33086
rect 40217 33083 40283 33086
rect 23841 33010 23907 33013
rect 31109 33010 31175 33013
rect 23841 33008 31175 33010
rect 23841 32952 23846 33008
rect 23902 32952 31114 33008
rect 31170 32952 31175 33008
rect 23841 32950 31175 32952
rect 23841 32947 23907 32950
rect 31109 32947 31175 32950
rect 32397 33010 32463 33013
rect 32857 33010 32923 33013
rect 36629 33010 36695 33013
rect 32397 33008 36695 33010
rect 32397 32952 32402 33008
rect 32458 32952 32862 33008
rect 32918 32952 36634 33008
rect 36690 32952 36695 33008
rect 32397 32950 36695 32952
rect 32397 32947 32463 32950
rect 32857 32947 32923 32950
rect 36629 32947 36695 32950
rect 20621 32874 20687 32877
rect 33777 32874 33843 32877
rect 20621 32872 33843 32874
rect 20621 32816 20626 32872
rect 20682 32816 33782 32872
rect 33838 32816 33843 32872
rect 20621 32814 33843 32816
rect 20621 32811 20687 32814
rect 33777 32811 33843 32814
rect 29862 32676 29868 32740
rect 29932 32738 29938 32740
rect 37457 32738 37523 32741
rect 29932 32736 37523 32738
rect 29932 32680 37462 32736
rect 37518 32680 37523 32736
rect 29932 32678 37523 32680
rect 29932 32676 29938 32678
rect 37457 32675 37523 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 20529 32602 20595 32605
rect 24945 32602 25011 32605
rect 20529 32600 25011 32602
rect 20529 32544 20534 32600
rect 20590 32544 24950 32600
rect 25006 32544 25011 32600
rect 20529 32542 25011 32544
rect 20529 32539 20595 32542
rect 24945 32539 25011 32542
rect 25078 32540 25084 32604
rect 25148 32602 25154 32604
rect 25221 32602 25287 32605
rect 28165 32602 28231 32605
rect 25148 32600 28231 32602
rect 25148 32544 25226 32600
rect 25282 32544 28170 32600
rect 28226 32544 28231 32600
rect 25148 32542 28231 32544
rect 25148 32540 25154 32542
rect 25221 32539 25287 32542
rect 28165 32539 28231 32542
rect 31201 32602 31267 32605
rect 35709 32602 35775 32605
rect 38745 32602 38811 32605
rect 31201 32600 38811 32602
rect 31201 32544 31206 32600
rect 31262 32544 35714 32600
rect 35770 32544 38750 32600
rect 38806 32544 38811 32600
rect 31201 32542 38811 32544
rect 31201 32539 31267 32542
rect 35709 32539 35775 32542
rect 38745 32539 38811 32542
rect 24301 32466 24367 32469
rect 26877 32466 26943 32469
rect 35157 32466 35223 32469
rect 35382 32466 35388 32468
rect 24301 32464 35388 32466
rect 24301 32408 24306 32464
rect 24362 32408 26882 32464
rect 26938 32408 35162 32464
rect 35218 32408 35388 32464
rect 24301 32406 35388 32408
rect 24301 32403 24367 32406
rect 26877 32403 26943 32406
rect 35157 32403 35223 32406
rect 35382 32404 35388 32406
rect 35452 32404 35458 32468
rect 24669 32330 24735 32333
rect 25221 32330 25287 32333
rect 24669 32328 25287 32330
rect 24669 32272 24674 32328
rect 24730 32272 25226 32328
rect 25282 32272 25287 32328
rect 24669 32270 25287 32272
rect 24669 32267 24735 32270
rect 25221 32267 25287 32270
rect 25405 32332 25471 32333
rect 25405 32328 25452 32332
rect 25516 32330 25522 32332
rect 32121 32330 32187 32333
rect 33685 32332 33751 32333
rect 36077 32332 36143 32333
rect 37365 32332 37431 32333
rect 32438 32330 32444 32332
rect 25405 32272 25410 32328
rect 25405 32268 25452 32272
rect 25516 32270 25562 32330
rect 32121 32328 32444 32330
rect 32121 32272 32126 32328
rect 32182 32272 32444 32328
rect 32121 32270 32444 32272
rect 25516 32268 25522 32270
rect 25405 32267 25471 32268
rect 32121 32267 32187 32270
rect 32438 32268 32444 32270
rect 32508 32268 32514 32332
rect 33685 32328 33732 32332
rect 33796 32330 33802 32332
rect 33685 32272 33690 32328
rect 33685 32268 33732 32272
rect 33796 32270 33842 32330
rect 36077 32328 36124 32332
rect 36188 32330 36194 32332
rect 36077 32272 36082 32328
rect 33796 32268 33802 32270
rect 36077 32268 36124 32272
rect 36188 32270 36234 32330
rect 37365 32328 37412 32332
rect 37476 32330 37482 32332
rect 37365 32272 37370 32328
rect 36188 32268 36194 32270
rect 37365 32268 37412 32272
rect 37476 32270 37522 32330
rect 37476 32268 37482 32270
rect 33685 32267 33751 32268
rect 36077 32267 36143 32268
rect 37365 32267 37431 32268
rect 37222 32132 37228 32196
rect 37292 32194 37298 32196
rect 38193 32194 38259 32197
rect 37292 32192 38259 32194
rect 37292 32136 38198 32192
rect 38254 32136 38259 32192
rect 37292 32134 38259 32136
rect 37292 32132 37298 32134
rect 38193 32131 38259 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 32029 32058 32095 32061
rect 33961 32058 34027 32061
rect 32029 32056 34027 32058
rect 32029 32000 32034 32056
rect 32090 32000 33966 32056
rect 34022 32000 34027 32056
rect 32029 31998 34027 32000
rect 32029 31995 32095 31998
rect 33961 31995 34027 31998
rect 36997 32058 37063 32061
rect 40902 32058 40908 32060
rect 36997 32056 40908 32058
rect 36997 32000 37002 32056
rect 37058 32000 40908 32056
rect 36997 31998 40908 32000
rect 36997 31995 37063 31998
rect 40902 31996 40908 31998
rect 40972 31996 40978 32060
rect 25262 31860 25268 31924
rect 25332 31922 25338 31924
rect 25405 31922 25471 31925
rect 25332 31920 25471 31922
rect 25332 31864 25410 31920
rect 25466 31864 25471 31920
rect 25332 31862 25471 31864
rect 25332 31860 25338 31862
rect 25405 31859 25471 31862
rect 33225 31922 33291 31925
rect 34094 31922 34100 31924
rect 33225 31920 34100 31922
rect 33225 31864 33230 31920
rect 33286 31864 34100 31920
rect 33225 31862 34100 31864
rect 33225 31859 33291 31862
rect 34094 31860 34100 31862
rect 34164 31860 34170 31924
rect 34605 31922 34671 31925
rect 36813 31922 36879 31925
rect 34605 31920 36879 31922
rect 34605 31864 34610 31920
rect 34666 31864 36818 31920
rect 36874 31864 36879 31920
rect 34605 31862 36879 31864
rect 34605 31859 34671 31862
rect 36813 31859 36879 31862
rect 38745 31922 38811 31925
rect 40493 31922 40559 31925
rect 41597 31922 41663 31925
rect 38745 31920 41663 31922
rect 38745 31864 38750 31920
rect 38806 31864 40498 31920
rect 40554 31864 41602 31920
rect 41658 31864 41663 31920
rect 38745 31862 41663 31864
rect 38745 31859 38811 31862
rect 40493 31859 40559 31862
rect 41597 31859 41663 31862
rect 16481 31786 16547 31789
rect 17585 31786 17651 31789
rect 21909 31786 21975 31789
rect 16481 31784 21975 31786
rect 16481 31728 16486 31784
rect 16542 31728 17590 31784
rect 17646 31728 21914 31784
rect 21970 31728 21975 31784
rect 16481 31726 21975 31728
rect 16481 31723 16547 31726
rect 17585 31723 17651 31726
rect 21909 31723 21975 31726
rect 25129 31786 25195 31789
rect 25262 31786 25268 31788
rect 25129 31784 25268 31786
rect 25129 31728 25134 31784
rect 25190 31728 25268 31784
rect 25129 31726 25268 31728
rect 25129 31723 25195 31726
rect 25262 31724 25268 31726
rect 25332 31724 25338 31788
rect 26785 31786 26851 31789
rect 27337 31786 27403 31789
rect 28901 31786 28967 31789
rect 36997 31786 37063 31789
rect 26785 31784 37063 31786
rect 26785 31728 26790 31784
rect 26846 31728 27342 31784
rect 27398 31728 28906 31784
rect 28962 31728 37002 31784
rect 37058 31728 37063 31784
rect 26785 31726 37063 31728
rect 26785 31723 26851 31726
rect 27337 31723 27403 31726
rect 28901 31723 28967 31726
rect 36997 31723 37063 31726
rect 40309 31786 40375 31789
rect 40585 31786 40651 31789
rect 40861 31786 40927 31789
rect 40309 31784 40927 31786
rect 40309 31728 40314 31784
rect 40370 31728 40590 31784
rect 40646 31728 40866 31784
rect 40922 31728 40927 31784
rect 40309 31726 40927 31728
rect 40309 31723 40375 31726
rect 40585 31723 40651 31726
rect 40861 31723 40927 31726
rect 34053 31652 34119 31653
rect 34053 31650 34100 31652
rect 34008 31648 34100 31650
rect 34008 31592 34058 31648
rect 34008 31590 34100 31592
rect 34053 31588 34100 31590
rect 34164 31588 34170 31652
rect 43989 31650 44055 31653
rect 44200 31650 45000 31740
rect 43989 31648 45000 31650
rect 43989 31592 43994 31648
rect 44050 31592 45000 31648
rect 43989 31590 45000 31592
rect 34053 31587 34119 31588
rect 43989 31587 44055 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 44200 31500 45000 31590
rect 31845 31378 31911 31381
rect 32070 31378 32076 31380
rect 31845 31376 32076 31378
rect 31845 31320 31850 31376
rect 31906 31320 32076 31376
rect 31845 31318 32076 31320
rect 31845 31315 31911 31318
rect 32070 31316 32076 31318
rect 32140 31316 32146 31380
rect 35709 31378 35775 31381
rect 36997 31378 37063 31381
rect 35709 31376 37063 31378
rect 35709 31320 35714 31376
rect 35770 31320 37002 31376
rect 37058 31320 37063 31376
rect 35709 31318 37063 31320
rect 35709 31315 35775 31318
rect 36997 31315 37063 31318
rect 18137 31242 18203 31245
rect 42701 31242 42767 31245
rect 18137 31240 42767 31242
rect 18137 31184 18142 31240
rect 18198 31184 42706 31240
rect 42762 31184 42767 31240
rect 18137 31182 42767 31184
rect 18137 31179 18203 31182
rect 42701 31179 42767 31182
rect 18229 31106 18295 31109
rect 18781 31106 18847 31109
rect 18229 31104 18847 31106
rect 18229 31048 18234 31104
rect 18290 31048 18786 31104
rect 18842 31048 18847 31104
rect 18229 31046 18847 31048
rect 18229 31043 18295 31046
rect 18781 31043 18847 31046
rect 19977 31106 20043 31109
rect 25037 31106 25103 31109
rect 19977 31104 25103 31106
rect 19977 31048 19982 31104
rect 20038 31048 25042 31104
rect 25098 31048 25103 31104
rect 19977 31046 25103 31048
rect 19977 31043 20043 31046
rect 25037 31043 25103 31046
rect 29729 31106 29795 31109
rect 30005 31106 30071 31109
rect 29729 31104 30071 31106
rect 29729 31048 29734 31104
rect 29790 31048 30010 31104
rect 30066 31048 30071 31104
rect 29729 31046 30071 31048
rect 29729 31043 29795 31046
rect 30005 31043 30071 31046
rect 35433 31106 35499 31109
rect 36445 31106 36511 31109
rect 38101 31106 38167 31109
rect 35433 31104 38167 31106
rect 35433 31048 35438 31104
rect 35494 31048 36450 31104
rect 36506 31048 38106 31104
rect 38162 31048 38167 31104
rect 35433 31046 38167 31048
rect 35433 31043 35499 31046
rect 36445 31043 36511 31046
rect 38101 31043 38167 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 29729 30970 29795 30973
rect 33317 30970 33383 30973
rect 29729 30968 33383 30970
rect 29729 30912 29734 30968
rect 29790 30912 33322 30968
rect 33378 30912 33383 30968
rect 29729 30910 33383 30912
rect 29729 30907 29795 30910
rect 33317 30907 33383 30910
rect 24945 30836 25011 30837
rect 24894 30834 24900 30836
rect 24854 30774 24900 30834
rect 24964 30832 25011 30836
rect 25006 30776 25011 30832
rect 24894 30772 24900 30774
rect 24964 30772 25011 30776
rect 24945 30771 25011 30772
rect 35341 30834 35407 30837
rect 42793 30834 42859 30837
rect 35341 30832 42859 30834
rect 35341 30776 35346 30832
rect 35402 30776 42798 30832
rect 42854 30776 42859 30832
rect 35341 30774 42859 30776
rect 35341 30771 35407 30774
rect 42793 30771 42859 30774
rect 39389 30698 39455 30701
rect 41781 30698 41847 30701
rect 42609 30698 42675 30701
rect 39389 30696 42675 30698
rect 39389 30640 39394 30696
rect 39450 30640 41786 30696
rect 41842 30640 42614 30696
rect 42670 30640 42675 30696
rect 39389 30638 42675 30640
rect 39389 30635 39455 30638
rect 41781 30635 41847 30638
rect 42609 30635 42675 30638
rect 27889 30564 27955 30565
rect 27838 30562 27844 30564
rect 27798 30502 27844 30562
rect 27908 30560 27955 30564
rect 27950 30504 27955 30560
rect 27838 30500 27844 30502
rect 27908 30500 27955 30504
rect 28758 30500 28764 30564
rect 28828 30562 28834 30564
rect 31937 30562 32003 30565
rect 28828 30560 32003 30562
rect 28828 30504 31942 30560
rect 31998 30504 32003 30560
rect 28828 30502 32003 30504
rect 28828 30500 28834 30502
rect 27889 30499 27955 30500
rect 31937 30499 32003 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 22093 30426 22159 30429
rect 33174 30426 33180 30428
rect 22093 30424 33180 30426
rect 22093 30368 22098 30424
rect 22154 30368 33180 30424
rect 22093 30366 33180 30368
rect 22093 30363 22159 30366
rect 33174 30364 33180 30366
rect 33244 30426 33250 30428
rect 34421 30426 34487 30429
rect 33244 30424 34487 30426
rect 33244 30368 34426 30424
rect 34482 30368 34487 30424
rect 33244 30366 34487 30368
rect 33244 30364 33250 30366
rect 34421 30363 34487 30366
rect 25865 30292 25931 30293
rect 28809 30292 28875 30293
rect 25814 30228 25820 30292
rect 25884 30290 25931 30292
rect 25884 30288 25976 30290
rect 25926 30232 25976 30288
rect 25884 30230 25976 30232
rect 25884 30228 25931 30230
rect 28758 30228 28764 30292
rect 28828 30290 28875 30292
rect 34513 30290 34579 30293
rect 42885 30290 42951 30293
rect 28828 30288 28920 30290
rect 28870 30232 28920 30288
rect 28828 30230 28920 30232
rect 34513 30288 42951 30290
rect 34513 30232 34518 30288
rect 34574 30232 42890 30288
rect 42946 30232 42951 30288
rect 34513 30230 42951 30232
rect 28828 30228 28875 30230
rect 25865 30227 25931 30228
rect 28809 30227 28875 30228
rect 34513 30227 34579 30230
rect 42885 30227 42951 30230
rect 31201 30154 31267 30157
rect 36353 30154 36419 30157
rect 38469 30154 38535 30157
rect 31201 30152 38535 30154
rect 31201 30096 31206 30152
rect 31262 30096 36358 30152
rect 36414 30096 38474 30152
rect 38530 30096 38535 30152
rect 31201 30094 38535 30096
rect 31201 30091 31267 30094
rect 36353 30091 36419 30094
rect 38469 30091 38535 30094
rect 36445 30018 36511 30021
rect 38285 30018 38351 30021
rect 36445 30016 38351 30018
rect 36445 29960 36450 30016
rect 36506 29960 38290 30016
rect 38346 29960 38351 30016
rect 36445 29958 38351 29960
rect 36445 29955 36511 29958
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 18873 29610 18939 29613
rect 19149 29610 19215 29613
rect 34513 29612 34579 29613
rect 34462 29610 34468 29612
rect 18873 29608 19215 29610
rect 18873 29552 18878 29608
rect 18934 29552 19154 29608
rect 19210 29552 19215 29608
rect 18873 29550 19215 29552
rect 34422 29550 34468 29610
rect 34532 29608 34579 29612
rect 34574 29552 34579 29608
rect 18873 29547 18939 29550
rect 19149 29547 19215 29550
rect 34462 29548 34468 29550
rect 34532 29548 34579 29552
rect 34513 29547 34579 29548
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 19977 29338 20043 29341
rect 24577 29338 24643 29341
rect 19977 29336 24643 29338
rect 19977 29280 19982 29336
rect 20038 29280 24582 29336
rect 24638 29280 24643 29336
rect 19977 29278 24643 29280
rect 19977 29275 20043 29278
rect 24577 29275 24643 29278
rect 18413 29202 18479 29205
rect 20069 29202 20135 29205
rect 35617 29204 35683 29205
rect 18413 29200 20135 29202
rect 18413 29144 18418 29200
rect 18474 29144 20074 29200
rect 20130 29144 20135 29200
rect 18413 29142 20135 29144
rect 18413 29139 18479 29142
rect 20069 29139 20135 29142
rect 35566 29140 35572 29204
rect 35636 29202 35683 29204
rect 35636 29200 35728 29202
rect 35678 29144 35728 29200
rect 35636 29142 35728 29144
rect 35636 29140 35683 29142
rect 35617 29139 35683 29140
rect 18137 29066 18203 29069
rect 18965 29066 19031 29069
rect 18137 29064 19031 29066
rect 18137 29008 18142 29064
rect 18198 29008 18970 29064
rect 19026 29008 19031 29064
rect 18137 29006 19031 29008
rect 18137 29003 18203 29006
rect 18965 29003 19031 29006
rect 24393 29066 24459 29069
rect 24526 29066 24532 29068
rect 24393 29064 24532 29066
rect 24393 29008 24398 29064
rect 24454 29008 24532 29064
rect 24393 29006 24532 29008
rect 24393 29003 24459 29006
rect 24526 29004 24532 29006
rect 24596 29004 24602 29068
rect 29729 29066 29795 29069
rect 33041 29066 33107 29069
rect 36353 29066 36419 29069
rect 39021 29068 39087 29069
rect 39205 29068 39271 29069
rect 39021 29066 39068 29068
rect 29729 29064 36419 29066
rect 29729 29008 29734 29064
rect 29790 29008 33046 29064
rect 33102 29008 36358 29064
rect 36414 29008 36419 29064
rect 29729 29006 36419 29008
rect 38976 29064 39068 29066
rect 38976 29008 39026 29064
rect 38976 29006 39068 29008
rect 29729 29003 29795 29006
rect 33041 29003 33107 29006
rect 36353 29003 36419 29006
rect 39021 29004 39068 29006
rect 39132 29004 39138 29068
rect 39205 29064 39252 29068
rect 39316 29066 39322 29068
rect 39205 29008 39210 29064
rect 39205 29004 39252 29008
rect 39316 29006 39362 29066
rect 39316 29004 39322 29006
rect 39021 29003 39087 29004
rect 39205 29003 39271 29004
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 35433 28524 35499 28525
rect 35382 28522 35388 28524
rect 35342 28462 35388 28522
rect 35452 28520 35499 28524
rect 35494 28464 35499 28520
rect 35382 28460 35388 28462
rect 35452 28460 35499 28464
rect 35433 28459 35499 28460
rect 30281 28386 30347 28389
rect 37222 28386 37228 28388
rect 30281 28384 37228 28386
rect 30281 28328 30286 28384
rect 30342 28328 37228 28384
rect 30281 28326 37228 28328
rect 30281 28323 30347 28326
rect 37222 28324 37228 28326
rect 37292 28324 37298 28388
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 32438 28188 32444 28252
rect 32508 28250 32514 28252
rect 33225 28250 33291 28253
rect 32508 28248 33291 28250
rect 32508 28192 33230 28248
rect 33286 28192 33291 28248
rect 32508 28190 33291 28192
rect 32508 28188 32514 28190
rect 33225 28187 33291 28190
rect 31477 28114 31543 28117
rect 35157 28114 35223 28117
rect 31477 28112 35223 28114
rect 31477 28056 31482 28112
rect 31538 28056 35162 28112
rect 35218 28056 35223 28112
rect 31477 28054 35223 28056
rect 31477 28051 31543 28054
rect 35157 28051 35223 28054
rect 34513 27978 34579 27981
rect 37457 27978 37523 27981
rect 34513 27976 37523 27978
rect 34513 27920 34518 27976
rect 34574 27920 37462 27976
rect 37518 27920 37523 27976
rect 34513 27918 37523 27920
rect 34513 27915 34579 27918
rect 37457 27915 37523 27918
rect 43989 27978 44055 27981
rect 44200 27978 45000 28068
rect 43989 27976 45000 27978
rect 43989 27920 43994 27976
rect 44050 27920 45000 27976
rect 43989 27918 45000 27920
rect 43989 27915 44055 27918
rect 44200 27828 45000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 26693 27708 26759 27709
rect 26693 27704 26740 27708
rect 26804 27706 26810 27708
rect 26693 27648 26698 27704
rect 26693 27644 26740 27648
rect 26804 27646 26850 27706
rect 26804 27644 26810 27646
rect 35934 27644 35940 27708
rect 36004 27706 36010 27708
rect 40534 27706 40540 27708
rect 36004 27646 40540 27706
rect 36004 27644 36010 27646
rect 40534 27644 40540 27646
rect 40604 27644 40610 27708
rect 26693 27643 26759 27644
rect 29913 27570 29979 27573
rect 34513 27570 34579 27573
rect 29913 27568 34579 27570
rect 29913 27512 29918 27568
rect 29974 27512 34518 27568
rect 34574 27512 34579 27568
rect 29913 27510 34579 27512
rect 29913 27507 29979 27510
rect 34513 27507 34579 27510
rect 36353 27570 36419 27573
rect 38193 27570 38259 27573
rect 36353 27568 38259 27570
rect 36353 27512 36358 27568
rect 36414 27512 38198 27568
rect 38254 27512 38259 27568
rect 36353 27510 38259 27512
rect 36353 27507 36419 27510
rect 38193 27507 38259 27510
rect 37222 27372 37228 27436
rect 37292 27434 37298 27436
rect 38326 27434 38332 27436
rect 37292 27374 38332 27434
rect 37292 27372 37298 27374
rect 38326 27372 38332 27374
rect 38396 27372 38402 27436
rect 39021 27434 39087 27437
rect 40309 27434 40375 27437
rect 39021 27432 40375 27434
rect 39021 27376 39026 27432
rect 39082 27376 40314 27432
rect 40370 27376 40375 27432
rect 39021 27374 40375 27376
rect 39021 27371 39087 27374
rect 40309 27371 40375 27374
rect 35985 27298 36051 27301
rect 38469 27298 38535 27301
rect 35985 27296 38535 27298
rect 35985 27240 35990 27296
rect 36046 27240 38474 27296
rect 38530 27240 38535 27296
rect 35985 27238 38535 27240
rect 35985 27235 36051 27238
rect 38469 27235 38535 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 37825 27026 37891 27029
rect 38285 27026 38351 27029
rect 37825 27024 38351 27026
rect 37825 26968 37830 27024
rect 37886 26968 38290 27024
rect 38346 26968 38351 27024
rect 37825 26966 38351 26968
rect 37825 26963 37891 26966
rect 38285 26963 38351 26966
rect 34329 26890 34395 26893
rect 38101 26890 38167 26893
rect 38377 26890 38443 26893
rect 34329 26888 38443 26890
rect 34329 26832 34334 26888
rect 34390 26832 38106 26888
rect 38162 26832 38382 26888
rect 38438 26832 38443 26888
rect 34329 26830 38443 26832
rect 34329 26827 34395 26830
rect 38101 26827 38167 26830
rect 38377 26827 38443 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 24301 26346 24367 26349
rect 30649 26346 30715 26349
rect 32438 26346 32444 26348
rect 24301 26344 32444 26346
rect 24301 26288 24306 26344
rect 24362 26288 30654 26344
rect 30710 26288 32444 26344
rect 24301 26286 32444 26288
rect 24301 26283 24367 26286
rect 30649 26283 30715 26286
rect 32438 26284 32444 26286
rect 32508 26346 32514 26348
rect 33317 26346 33383 26349
rect 32508 26344 33383 26346
rect 32508 26288 33322 26344
rect 33378 26288 33383 26344
rect 32508 26286 33383 26288
rect 32508 26284 32514 26286
rect 33317 26283 33383 26286
rect 33777 26346 33843 26349
rect 35249 26346 35315 26349
rect 35382 26346 35388 26348
rect 33777 26344 35388 26346
rect 33777 26288 33782 26344
rect 33838 26288 35254 26344
rect 35310 26288 35388 26344
rect 33777 26286 35388 26288
rect 33777 26283 33843 26286
rect 35249 26283 35315 26286
rect 35382 26284 35388 26286
rect 35452 26284 35458 26348
rect 37222 26284 37228 26348
rect 37292 26346 37298 26348
rect 37917 26346 37983 26349
rect 37292 26344 37983 26346
rect 37292 26288 37922 26344
rect 37978 26288 37983 26344
rect 37292 26286 37983 26288
rect 37292 26284 37298 26286
rect 37917 26283 37983 26286
rect 34053 26212 34119 26213
rect 34053 26210 34100 26212
rect 34008 26208 34100 26210
rect 34008 26152 34058 26208
rect 34008 26150 34100 26152
rect 34053 26148 34100 26150
rect 34164 26148 34170 26212
rect 34421 26210 34487 26213
rect 37457 26210 37523 26213
rect 38469 26210 38535 26213
rect 34421 26208 38535 26210
rect 34421 26152 34426 26208
rect 34482 26152 37462 26208
rect 37518 26152 38474 26208
rect 38530 26152 38535 26208
rect 34421 26150 38535 26152
rect 34053 26147 34119 26148
rect 34421 26147 34487 26150
rect 37457 26147 37523 26150
rect 38469 26147 38535 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 20529 26074 20595 26077
rect 25446 26074 25452 26076
rect 20529 26072 25452 26074
rect 20529 26016 20534 26072
rect 20590 26016 25452 26072
rect 20529 26014 25452 26016
rect 20529 26011 20595 26014
rect 25446 26012 25452 26014
rect 25516 26012 25522 26076
rect 33041 26074 33107 26077
rect 35934 26074 35940 26076
rect 33041 26072 35940 26074
rect 33041 26016 33046 26072
rect 33102 26016 35940 26072
rect 33041 26014 35940 26016
rect 33041 26011 33107 26014
rect 35934 26012 35940 26014
rect 36004 26012 36010 26076
rect 39205 25938 39271 25941
rect 43069 25938 43135 25941
rect 39205 25936 43135 25938
rect 39205 25880 39210 25936
rect 39266 25880 43074 25936
rect 43130 25880 43135 25936
rect 39205 25878 43135 25880
rect 39205 25875 39271 25878
rect 43069 25875 43135 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 37365 25532 37431 25533
rect 37365 25530 37412 25532
rect 37320 25528 37412 25530
rect 37320 25472 37370 25528
rect 37320 25470 37412 25472
rect 37365 25468 37412 25470
rect 37476 25468 37482 25532
rect 37365 25467 37431 25468
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 32305 24850 32371 24853
rect 35985 24850 36051 24853
rect 37089 24850 37155 24853
rect 32305 24848 37155 24850
rect 32305 24792 32310 24848
rect 32366 24792 35990 24848
rect 36046 24792 37094 24848
rect 37150 24792 37155 24848
rect 32305 24790 37155 24792
rect 32305 24787 32371 24790
rect 35985 24787 36051 24790
rect 37089 24787 37155 24790
rect 32029 24714 32095 24717
rect 37549 24714 37615 24717
rect 37825 24714 37891 24717
rect 32029 24712 37891 24714
rect 32029 24656 32034 24712
rect 32090 24656 37554 24712
rect 37610 24656 37830 24712
rect 37886 24656 37891 24712
rect 32029 24654 37891 24656
rect 32029 24651 32095 24654
rect 37549 24651 37615 24654
rect 37825 24651 37891 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 37406 24380 37412 24444
rect 37476 24442 37482 24444
rect 40033 24442 40099 24445
rect 40401 24444 40467 24445
rect 37476 24440 40099 24442
rect 37476 24384 40038 24440
rect 40094 24384 40099 24440
rect 37476 24382 40099 24384
rect 37476 24380 37482 24382
rect 40033 24379 40099 24382
rect 40350 24380 40356 24444
rect 40420 24442 40467 24444
rect 40420 24440 40512 24442
rect 40462 24384 40512 24440
rect 40420 24382 40512 24384
rect 40420 24380 40467 24382
rect 40401 24379 40467 24380
rect 34237 24306 34303 24309
rect 34462 24306 34468 24308
rect 34237 24304 34468 24306
rect 34237 24248 34242 24304
rect 34298 24248 34468 24304
rect 34237 24246 34468 24248
rect 34237 24243 34303 24246
rect 34462 24244 34468 24246
rect 34532 24244 34538 24308
rect 37089 24306 37155 24309
rect 38009 24306 38075 24309
rect 37089 24304 38075 24306
rect 37089 24248 37094 24304
rect 37150 24248 38014 24304
rect 38070 24248 38075 24304
rect 37089 24246 38075 24248
rect 37089 24243 37155 24246
rect 38009 24243 38075 24246
rect 43989 24306 44055 24309
rect 44200 24306 45000 24396
rect 43989 24304 45000 24306
rect 43989 24248 43994 24304
rect 44050 24248 45000 24304
rect 43989 24246 45000 24248
rect 43989 24243 44055 24246
rect 28349 24170 28415 24173
rect 40953 24172 41019 24173
rect 40902 24170 40908 24172
rect 28349 24168 40908 24170
rect 40972 24170 41019 24172
rect 40972 24168 41064 24170
rect 28349 24112 28354 24168
rect 28410 24112 40908 24168
rect 41014 24112 41064 24168
rect 44200 24156 45000 24246
rect 28349 24110 40908 24112
rect 28349 24107 28415 24110
rect 40902 24108 40908 24110
rect 40972 24110 41064 24112
rect 40972 24108 41019 24110
rect 40953 24107 41019 24108
rect 36261 24034 36327 24037
rect 37825 24034 37891 24037
rect 36261 24032 37891 24034
rect 36261 23976 36266 24032
rect 36322 23976 37830 24032
rect 37886 23976 37891 24032
rect 36261 23974 37891 23976
rect 36261 23971 36327 23974
rect 37825 23971 37891 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 34145 23898 34211 23901
rect 34145 23896 36370 23898
rect 34145 23840 34150 23896
rect 34206 23840 36370 23896
rect 34145 23838 36370 23840
rect 34145 23835 34211 23838
rect 31845 23764 31911 23765
rect 31845 23760 31892 23764
rect 31956 23762 31962 23764
rect 32673 23762 32739 23765
rect 35566 23762 35572 23764
rect 31845 23704 31850 23760
rect 31845 23700 31892 23704
rect 31956 23702 32002 23762
rect 32673 23760 35572 23762
rect 32673 23704 32678 23760
rect 32734 23704 35572 23760
rect 32673 23702 35572 23704
rect 31956 23700 31962 23702
rect 31845 23699 31911 23700
rect 32673 23699 32739 23702
rect 35566 23700 35572 23702
rect 35636 23762 35642 23764
rect 36310 23762 36370 23838
rect 37089 23762 37155 23765
rect 38929 23762 38995 23765
rect 39389 23762 39455 23765
rect 35636 23702 36186 23762
rect 36310 23760 39455 23762
rect 36310 23704 37094 23760
rect 37150 23704 38934 23760
rect 38990 23704 39394 23760
rect 39450 23704 39455 23760
rect 36310 23702 39455 23704
rect 35636 23700 35642 23702
rect 36126 23626 36186 23702
rect 37089 23699 37155 23702
rect 38929 23699 38995 23702
rect 39389 23699 39455 23702
rect 36261 23626 36327 23629
rect 36126 23624 36327 23626
rect 36126 23568 36266 23624
rect 36322 23568 36327 23624
rect 36126 23566 36327 23568
rect 36261 23563 36327 23566
rect 36537 23626 36603 23629
rect 37825 23626 37891 23629
rect 36537 23624 37891 23626
rect 36537 23568 36542 23624
rect 36598 23568 37830 23624
rect 37886 23568 37891 23624
rect 36537 23566 37891 23568
rect 36537 23563 36603 23566
rect 37825 23563 37891 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 35433 23354 35499 23357
rect 37181 23354 37247 23357
rect 38009 23354 38075 23357
rect 35433 23352 38075 23354
rect 35433 23296 35438 23352
rect 35494 23296 37186 23352
rect 37242 23296 38014 23352
rect 38070 23296 38075 23352
rect 35433 23294 38075 23296
rect 35433 23291 35499 23294
rect 37181 23291 37247 23294
rect 38009 23291 38075 23294
rect 33133 23220 33199 23221
rect 33133 23218 33180 23220
rect 33088 23216 33180 23218
rect 33088 23160 33138 23216
rect 33088 23158 33180 23160
rect 33133 23156 33180 23158
rect 33244 23156 33250 23220
rect 33133 23155 33199 23156
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 39430 22748 39436 22812
rect 39500 22810 39506 22812
rect 39665 22810 39731 22813
rect 39500 22808 39731 22810
rect 39500 22752 39670 22808
rect 39726 22752 39731 22808
rect 39500 22750 39731 22752
rect 39500 22748 39506 22750
rect 39665 22747 39731 22750
rect 32397 22674 32463 22677
rect 36629 22674 36695 22677
rect 32397 22672 36695 22674
rect 32397 22616 32402 22672
rect 32458 22616 36634 22672
rect 36690 22616 36695 22672
rect 32397 22614 36695 22616
rect 32397 22611 32463 22614
rect 36629 22611 36695 22614
rect 36813 22674 36879 22677
rect 37222 22674 37228 22676
rect 36813 22672 37228 22674
rect 36813 22616 36818 22672
rect 36874 22616 37228 22672
rect 36813 22614 37228 22616
rect 36813 22611 36879 22614
rect 37222 22612 37228 22614
rect 37292 22612 37298 22676
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 32305 22266 32371 22269
rect 32438 22266 32444 22268
rect 32305 22264 32444 22266
rect 32305 22208 32310 22264
rect 32366 22208 32444 22264
rect 32305 22206 32444 22208
rect 32305 22203 32371 22206
rect 32438 22204 32444 22206
rect 32508 22204 32514 22268
rect 28993 22130 29059 22133
rect 32029 22130 32095 22133
rect 28993 22128 32095 22130
rect 28993 22072 28998 22128
rect 29054 22072 32034 22128
rect 32090 22072 32095 22128
rect 28993 22070 32095 22072
rect 28993 22067 29059 22070
rect 32029 22067 32095 22070
rect 39665 22130 39731 22133
rect 41321 22130 41387 22133
rect 39665 22128 41387 22130
rect 39665 22072 39670 22128
rect 39726 22072 41326 22128
rect 41382 22072 41387 22128
rect 39665 22070 41387 22072
rect 39665 22067 39731 22070
rect 41321 22067 41387 22070
rect 28809 21994 28875 21997
rect 31385 21994 31451 21997
rect 28809 21992 31451 21994
rect 28809 21936 28814 21992
rect 28870 21936 31390 21992
rect 31446 21936 31451 21992
rect 28809 21934 31451 21936
rect 28809 21931 28875 21934
rect 31385 21931 31451 21934
rect 37181 21994 37247 21997
rect 39062 21994 39068 21996
rect 37181 21992 39068 21994
rect 37181 21936 37186 21992
rect 37242 21936 39068 21992
rect 37181 21934 39068 21936
rect 37181 21931 37247 21934
rect 39062 21932 39068 21934
rect 39132 21932 39138 21996
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 41321 20772 41387 20773
rect 41270 20770 41276 20772
rect 41230 20710 41276 20770
rect 41340 20768 41387 20772
rect 41382 20712 41387 20768
rect 41270 20708 41276 20710
rect 41340 20708 41387 20712
rect 41321 20707 41387 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 27429 20634 27495 20637
rect 29729 20634 29795 20637
rect 35341 20634 35407 20637
rect 27429 20632 35407 20634
rect 27429 20576 27434 20632
rect 27490 20576 29734 20632
rect 29790 20576 35346 20632
rect 35402 20576 35407 20632
rect 27429 20574 35407 20576
rect 27429 20571 27495 20574
rect 29729 20571 29795 20574
rect 35341 20571 35407 20574
rect 43989 20634 44055 20637
rect 44200 20634 45000 20724
rect 43989 20632 45000 20634
rect 43989 20576 43994 20632
rect 44050 20576 45000 20632
rect 43989 20574 45000 20576
rect 43989 20571 44055 20574
rect 44200 20484 45000 20574
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 26141 19954 26207 19957
rect 28901 19954 28967 19957
rect 26141 19952 28967 19954
rect 26141 19896 26146 19952
rect 26202 19896 28906 19952
rect 28962 19896 28967 19952
rect 26141 19894 28967 19896
rect 26141 19891 26207 19894
rect 28901 19891 28967 19894
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 22737 19546 22803 19549
rect 25262 19546 25268 19548
rect 22737 19544 25268 19546
rect 22737 19488 22742 19544
rect 22798 19488 25268 19544
rect 22737 19486 25268 19488
rect 22737 19483 22803 19486
rect 25262 19484 25268 19486
rect 25332 19484 25338 19548
rect 33726 19348 33732 19412
rect 33796 19410 33802 19412
rect 33961 19410 34027 19413
rect 33796 19408 34027 19410
rect 33796 19352 33966 19408
rect 34022 19352 34027 19408
rect 33796 19350 34027 19352
rect 33796 19348 33802 19350
rect 33961 19347 34027 19350
rect 39665 19410 39731 19413
rect 40769 19410 40835 19413
rect 39665 19408 40835 19410
rect 39665 19352 39670 19408
rect 39726 19352 40774 19408
rect 40830 19352 40835 19408
rect 39665 19350 40835 19352
rect 39665 19347 39731 19350
rect 40769 19347 40835 19350
rect 17861 19274 17927 19277
rect 26182 19274 26188 19276
rect 17861 19272 26188 19274
rect 17861 19216 17866 19272
rect 17922 19216 26188 19272
rect 17861 19214 26188 19216
rect 17861 19211 17927 19214
rect 26182 19212 26188 19214
rect 26252 19212 26258 19276
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 39297 19004 39363 19005
rect 39246 18940 39252 19004
rect 39316 19002 39363 19004
rect 39316 19000 39408 19002
rect 39358 18944 39408 19000
rect 39316 18942 39408 18944
rect 39316 18940 39363 18942
rect 39297 18939 39363 18940
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 27981 17778 28047 17781
rect 39941 17778 40007 17781
rect 27981 17776 40007 17778
rect 27981 17720 27986 17776
rect 28042 17720 39946 17776
rect 40002 17720 40007 17776
rect 27981 17718 40007 17720
rect 27981 17715 28047 17718
rect 39941 17715 40007 17718
rect 17217 17642 17283 17645
rect 28758 17642 28764 17644
rect 17217 17640 28764 17642
rect 17217 17584 17222 17640
rect 17278 17584 28764 17640
rect 17217 17582 28764 17584
rect 17217 17579 17283 17582
rect 28758 17580 28764 17582
rect 28828 17580 28834 17644
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 43989 16962 44055 16965
rect 44200 16962 45000 17052
rect 43989 16960 45000 16962
rect 43989 16904 43994 16960
rect 44050 16904 45000 16960
rect 43989 16902 45000 16904
rect 43989 16899 44055 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 24577 16828 24643 16829
rect 24526 16764 24532 16828
rect 24596 16826 24643 16828
rect 24596 16824 24688 16826
rect 24638 16768 24688 16824
rect 44200 16812 45000 16902
rect 24596 16766 24688 16768
rect 24596 16764 24643 16766
rect 24577 16763 24643 16764
rect 27889 16554 27955 16557
rect 34145 16554 34211 16557
rect 35249 16554 35315 16557
rect 27889 16552 35315 16554
rect 27889 16496 27894 16552
rect 27950 16496 34150 16552
rect 34206 16496 35254 16552
rect 35310 16496 35315 16552
rect 27889 16494 35315 16496
rect 27889 16491 27955 16494
rect 34145 16491 34211 16494
rect 35249 16491 35315 16494
rect 32305 16418 32371 16421
rect 34881 16418 34947 16421
rect 32305 16416 34947 16418
rect 32305 16360 32310 16416
rect 32366 16360 34886 16416
rect 34942 16360 34947 16416
rect 32305 16358 34947 16360
rect 32305 16355 32371 16358
rect 34881 16355 34947 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 26601 16282 26667 16285
rect 26734 16282 26740 16284
rect 26601 16280 26740 16282
rect 26601 16224 26606 16280
rect 26662 16224 26740 16280
rect 26601 16222 26740 16224
rect 26601 16219 26667 16222
rect 26734 16220 26740 16222
rect 26804 16220 26810 16284
rect 32581 16146 32647 16149
rect 36169 16146 36235 16149
rect 37089 16146 37155 16149
rect 32581 16144 37155 16146
rect 32581 16088 32586 16144
rect 32642 16088 36174 16144
rect 36230 16088 37094 16144
rect 37150 16088 37155 16144
rect 32581 16086 37155 16088
rect 32581 16083 32647 16086
rect 36169 16083 36235 16086
rect 37089 16083 37155 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 36118 15540 36124 15604
rect 36188 15602 36194 15604
rect 39205 15602 39271 15605
rect 36188 15600 39271 15602
rect 36188 15544 39210 15600
rect 39266 15544 39271 15600
rect 36188 15542 39271 15544
rect 36188 15540 36194 15542
rect 39205 15539 39271 15542
rect 26049 15330 26115 15333
rect 27838 15330 27844 15332
rect 26049 15328 27844 15330
rect 26049 15272 26054 15328
rect 26110 15272 27844 15328
rect 26049 15270 27844 15272
rect 26049 15267 26115 15270
rect 27838 15268 27844 15270
rect 27908 15268 27914 15332
rect 32489 15330 32555 15333
rect 33501 15330 33567 15333
rect 36721 15330 36787 15333
rect 32489 15328 36787 15330
rect 32489 15272 32494 15328
rect 32550 15272 33506 15328
rect 33562 15272 36726 15328
rect 36782 15272 36787 15328
rect 32489 15270 36787 15272
rect 32489 15267 32555 15270
rect 33501 15267 33567 15270
rect 36721 15267 36787 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 28809 15194 28875 15197
rect 29177 15194 29243 15197
rect 28809 15192 29243 15194
rect 28809 15136 28814 15192
rect 28870 15136 29182 15192
rect 29238 15136 29243 15192
rect 28809 15134 29243 15136
rect 28809 15131 28875 15134
rect 29177 15131 29243 15134
rect 33317 15058 33383 15061
rect 35893 15058 35959 15061
rect 33317 15056 35959 15058
rect 33317 15000 33322 15056
rect 33378 15000 35898 15056
rect 35954 15000 35959 15056
rect 33317 14998 35959 15000
rect 33317 14995 33383 14998
rect 35893 14995 35959 14998
rect 29821 14922 29887 14925
rect 35065 14922 35131 14925
rect 35801 14922 35867 14925
rect 29821 14920 35867 14922
rect 29821 14864 29826 14920
rect 29882 14864 35070 14920
rect 35126 14864 35806 14920
rect 35862 14864 35867 14920
rect 29821 14862 35867 14864
rect 29821 14859 29887 14862
rect 35065 14859 35131 14862
rect 35801 14859 35867 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 35065 14514 35131 14517
rect 35617 14514 35683 14517
rect 38193 14514 38259 14517
rect 35065 14512 38259 14514
rect 35065 14456 35070 14512
rect 35126 14456 35622 14512
rect 35678 14456 38198 14512
rect 38254 14456 38259 14512
rect 35065 14454 38259 14456
rect 35065 14451 35131 14454
rect 35617 14451 35683 14454
rect 38193 14451 38259 14454
rect 26969 14378 27035 14381
rect 43069 14378 43135 14381
rect 26969 14376 43135 14378
rect 26969 14320 26974 14376
rect 27030 14320 43074 14376
rect 43130 14320 43135 14376
rect 26969 14318 43135 14320
rect 26969 14315 27035 14318
rect 43069 14315 43135 14318
rect 31661 14242 31727 14245
rect 33317 14242 33383 14245
rect 31661 14240 33383 14242
rect 31661 14184 31666 14240
rect 31722 14184 33322 14240
rect 33378 14184 33383 14240
rect 31661 14182 33383 14184
rect 31661 14179 31727 14182
rect 33317 14179 33383 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 41229 14108 41295 14109
rect 41229 14106 41276 14108
rect 41184 14104 41276 14106
rect 41184 14048 41234 14104
rect 41184 14046 41276 14048
rect 41229 14044 41276 14046
rect 41340 14044 41346 14108
rect 41229 14043 41295 14044
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 42793 13290 42859 13293
rect 43345 13290 43411 13293
rect 44200 13290 45000 13380
rect 42793 13288 45000 13290
rect 42793 13232 42798 13288
rect 42854 13232 43350 13288
rect 43406 13232 45000 13288
rect 42793 13230 45000 13232
rect 42793 13227 42859 13230
rect 43345 13227 43411 13230
rect 44200 13140 45000 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 31886 12004 31892 12068
rect 31956 12066 31962 12068
rect 39113 12066 39179 12069
rect 39665 12066 39731 12069
rect 31956 12064 39731 12066
rect 31956 12008 39118 12064
rect 39174 12008 39670 12064
rect 39726 12008 39731 12064
rect 31956 12006 39731 12008
rect 31956 12004 31962 12006
rect 39113 12003 39179 12006
rect 39665 12003 39731 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 38326 11868 38332 11932
rect 38396 11930 38402 11932
rect 40861 11930 40927 11933
rect 38396 11928 40927 11930
rect 38396 11872 40866 11928
rect 40922 11872 40927 11928
rect 38396 11870 40927 11872
rect 38396 11868 38402 11870
rect 40861 11867 40927 11870
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 32213 11386 32279 11389
rect 32438 11386 32444 11388
rect 32213 11384 32444 11386
rect 32213 11328 32218 11384
rect 32274 11328 32444 11384
rect 32213 11326 32444 11328
rect 32213 11323 32279 11326
rect 32438 11324 32444 11326
rect 32508 11386 32514 11388
rect 32857 11386 32923 11389
rect 32508 11384 32923 11386
rect 32508 11328 32862 11384
rect 32918 11328 32923 11384
rect 32508 11326 32923 11328
rect 32508 11324 32514 11326
rect 32857 11323 32923 11326
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 43989 9618 44055 9621
rect 44200 9618 45000 9708
rect 43989 9616 45000 9618
rect 43989 9560 43994 9616
rect 44050 9560 45000 9616
rect 43989 9558 45000 9560
rect 43989 9555 44055 9558
rect 44200 9468 45000 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 43345 5946 43411 5949
rect 44200 5946 45000 6036
rect 43345 5944 45000 5946
rect 43345 5888 43350 5944
rect 43406 5888 45000 5944
rect 43345 5886 45000 5888
rect 43345 5883 43411 5886
rect 44200 5796 45000 5886
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 43989 2274 44055 2277
rect 44200 2274 45000 2364
rect 43989 2272 45000 2274
rect 43989 2216 43994 2272
rect 44050 2216 45000 2272
rect 43989 2214 45000 2216
rect 43989 2211 44055 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 44200 2124 45000 2214
<< via3 >>
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 28764 39884 28828 39948
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 33180 39264 33244 39268
rect 33180 39208 33230 39264
rect 33230 39208 33244 39264
rect 33180 39204 33244 39208
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 27476 38992 27540 38996
rect 27476 38936 27526 38992
rect 27526 38936 27540 38992
rect 27476 38932 27540 38936
rect 40540 38932 40604 38996
rect 28764 38660 28828 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 28580 38388 28644 38452
rect 24900 38116 24964 38180
rect 35388 38116 35452 38180
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 36308 37708 36372 37772
rect 27292 37572 27356 37636
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 29868 37572 29932 37636
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 37228 37436 37292 37500
rect 25084 37300 25148 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 33180 36892 33244 36956
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 25820 36212 25884 36276
rect 37228 36212 37292 36276
rect 24900 36076 24964 36140
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 27476 35592 27540 35596
rect 27476 35536 27526 35592
rect 27526 35536 27540 35592
rect 27476 35532 27540 35536
rect 40908 35592 40972 35596
rect 40908 35536 40922 35592
rect 40922 35536 40972 35592
rect 40908 35532 40972 35536
rect 32076 35396 32140 35460
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 28764 34988 28828 35052
rect 32076 34852 32140 34916
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 34100 34580 34164 34644
rect 27292 34504 27356 34508
rect 27292 34448 27342 34504
rect 27342 34448 27356 34504
rect 27292 34444 27356 34448
rect 36308 34444 36372 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 28580 34172 28644 34236
rect 25268 33824 25332 33828
rect 25268 33768 25282 33824
rect 25282 33768 25332 33824
rect 25268 33764 25332 33768
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 37228 33628 37292 33692
rect 39436 33552 39500 33556
rect 39436 33496 39450 33552
rect 39450 33496 39500 33552
rect 39436 33492 39500 33496
rect 26188 33356 26252 33420
rect 40356 33220 40420 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 29868 32676 29932 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 25084 32540 25148 32604
rect 35388 32404 35452 32468
rect 25452 32328 25516 32332
rect 25452 32272 25466 32328
rect 25466 32272 25516 32328
rect 25452 32268 25516 32272
rect 32444 32268 32508 32332
rect 33732 32328 33796 32332
rect 33732 32272 33746 32328
rect 33746 32272 33796 32328
rect 33732 32268 33796 32272
rect 36124 32328 36188 32332
rect 36124 32272 36138 32328
rect 36138 32272 36188 32328
rect 36124 32268 36188 32272
rect 37412 32328 37476 32332
rect 37412 32272 37426 32328
rect 37426 32272 37476 32328
rect 37412 32268 37476 32272
rect 37228 32132 37292 32196
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 40908 31996 40972 32060
rect 25268 31860 25332 31924
rect 34100 31860 34164 31924
rect 25268 31724 25332 31788
rect 34100 31648 34164 31652
rect 34100 31592 34114 31648
rect 34114 31592 34164 31648
rect 34100 31588 34164 31592
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 32076 31316 32140 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 24900 30832 24964 30836
rect 24900 30776 24950 30832
rect 24950 30776 24964 30832
rect 24900 30772 24964 30776
rect 27844 30560 27908 30564
rect 27844 30504 27894 30560
rect 27894 30504 27908 30560
rect 27844 30500 27908 30504
rect 28764 30500 28828 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 33180 30364 33244 30428
rect 25820 30288 25884 30292
rect 25820 30232 25870 30288
rect 25870 30232 25884 30288
rect 25820 30228 25884 30232
rect 28764 30288 28828 30292
rect 28764 30232 28814 30288
rect 28814 30232 28828 30288
rect 28764 30228 28828 30232
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 34468 29608 34532 29612
rect 34468 29552 34518 29608
rect 34518 29552 34532 29608
rect 34468 29548 34532 29552
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 35572 29200 35636 29204
rect 35572 29144 35622 29200
rect 35622 29144 35636 29200
rect 35572 29140 35636 29144
rect 24532 29004 24596 29068
rect 39068 29064 39132 29068
rect 39068 29008 39082 29064
rect 39082 29008 39132 29064
rect 39068 29004 39132 29008
rect 39252 29064 39316 29068
rect 39252 29008 39266 29064
rect 39266 29008 39316 29064
rect 39252 29004 39316 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 35388 28520 35452 28524
rect 35388 28464 35438 28520
rect 35438 28464 35452 28520
rect 35388 28460 35452 28464
rect 37228 28324 37292 28388
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 32444 28188 32508 28252
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 26740 27704 26804 27708
rect 26740 27648 26754 27704
rect 26754 27648 26804 27704
rect 26740 27644 26804 27648
rect 35940 27644 36004 27708
rect 40540 27644 40604 27708
rect 37228 27372 37292 27436
rect 38332 27372 38396 27436
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 32444 26284 32508 26348
rect 35388 26284 35452 26348
rect 37228 26284 37292 26348
rect 34100 26208 34164 26212
rect 34100 26152 34114 26208
rect 34114 26152 34164 26208
rect 34100 26148 34164 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 25452 26012 25516 26076
rect 35940 26012 36004 26076
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 37412 25528 37476 25532
rect 37412 25472 37426 25528
rect 37426 25472 37476 25528
rect 37412 25468 37476 25472
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 37412 24380 37476 24444
rect 40356 24440 40420 24444
rect 40356 24384 40406 24440
rect 40406 24384 40420 24440
rect 40356 24380 40420 24384
rect 34468 24244 34532 24308
rect 40908 24168 40972 24172
rect 40908 24112 40958 24168
rect 40958 24112 40972 24168
rect 40908 24108 40972 24112
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 31892 23760 31956 23764
rect 31892 23704 31906 23760
rect 31906 23704 31956 23760
rect 31892 23700 31956 23704
rect 35572 23700 35636 23764
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 33180 23216 33244 23220
rect 33180 23160 33194 23216
rect 33194 23160 33244 23216
rect 33180 23156 33244 23160
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 39436 22748 39500 22812
rect 37228 22612 37292 22676
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 32444 22204 32508 22268
rect 39068 21932 39132 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 41276 20768 41340 20772
rect 41276 20712 41326 20768
rect 41326 20712 41340 20768
rect 41276 20708 41340 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 25268 19484 25332 19548
rect 33732 19348 33796 19412
rect 26188 19212 26252 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 39252 19000 39316 19004
rect 39252 18944 39302 19000
rect 39302 18944 39316 19000
rect 39252 18940 39316 18944
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 28764 17580 28828 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 24532 16824 24596 16828
rect 24532 16768 24582 16824
rect 24582 16768 24596 16824
rect 24532 16764 24596 16768
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 26740 16220 26804 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 36124 15540 36188 15604
rect 27844 15268 27908 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 41276 14104 41340 14108
rect 41276 14048 41290 14104
rect 41290 14048 41340 14104
rect 41276 14044 41340 14048
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 31892 12004 31956 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 38332 11868 38396 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 32444 11324 32508 11388
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 41920 4528 42480
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 42464 19888 42480
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 34928 41920 35248 42480
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 28763 39948 28829 39949
rect 28763 39884 28764 39948
rect 28828 39884 28829 39948
rect 28763 39883 28829 39884
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 27475 38996 27541 38997
rect 27475 38932 27476 38996
rect 27540 38932 27541 38996
rect 27475 38931 27541 38932
rect 24899 38180 24965 38181
rect 24899 38116 24900 38180
rect 24964 38116 24965 38180
rect 24899 38115 24965 38116
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 24902 36141 24962 38115
rect 27291 37636 27357 37637
rect 27291 37572 27292 37636
rect 27356 37572 27357 37636
rect 27291 37571 27357 37572
rect 25083 37364 25149 37365
rect 25083 37300 25084 37364
rect 25148 37300 25149 37364
rect 25083 37299 25149 37300
rect 24899 36140 24965 36141
rect 24899 36076 24900 36140
rect 24964 36076 24965 36140
rect 24899 36075 24965 36076
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 24902 30837 24962 36075
rect 25086 32605 25146 37299
rect 25819 36276 25885 36277
rect 25819 36212 25820 36276
rect 25884 36212 25885 36276
rect 25819 36211 25885 36212
rect 25267 33828 25333 33829
rect 25267 33764 25268 33828
rect 25332 33764 25333 33828
rect 25267 33763 25333 33764
rect 25083 32604 25149 32605
rect 25083 32540 25084 32604
rect 25148 32540 25149 32604
rect 25083 32539 25149 32540
rect 25270 31925 25330 33763
rect 25451 32332 25517 32333
rect 25451 32268 25452 32332
rect 25516 32268 25517 32332
rect 25451 32267 25517 32268
rect 25267 31924 25333 31925
rect 25267 31860 25268 31924
rect 25332 31860 25333 31924
rect 25267 31859 25333 31860
rect 25267 31788 25333 31789
rect 25267 31724 25268 31788
rect 25332 31724 25333 31788
rect 25267 31723 25333 31724
rect 24899 30836 24965 30837
rect 24899 30772 24900 30836
rect 24964 30772 24965 30836
rect 24899 30771 24965 30772
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 24531 29068 24597 29069
rect 24531 29004 24532 29068
rect 24596 29004 24597 29068
rect 24531 29003 24597 29004
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 24534 16829 24594 29003
rect 25270 19549 25330 31723
rect 25454 26077 25514 32267
rect 25822 30293 25882 36211
rect 27294 34509 27354 37571
rect 27478 35597 27538 38931
rect 28766 38725 28826 39883
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 33179 39268 33245 39269
rect 33179 39204 33180 39268
rect 33244 39204 33245 39268
rect 33179 39203 33245 39204
rect 28763 38724 28829 38725
rect 28763 38660 28764 38724
rect 28828 38660 28829 38724
rect 28763 38659 28829 38660
rect 28579 38452 28645 38453
rect 28579 38388 28580 38452
rect 28644 38388 28645 38452
rect 28579 38387 28645 38388
rect 27475 35596 27541 35597
rect 27475 35532 27476 35596
rect 27540 35532 27541 35596
rect 27475 35531 27541 35532
rect 27291 34508 27357 34509
rect 27291 34444 27292 34508
rect 27356 34444 27357 34508
rect 27291 34443 27357 34444
rect 28582 34237 28642 38387
rect 28766 35053 28826 38659
rect 29867 37636 29933 37637
rect 29867 37572 29868 37636
rect 29932 37572 29933 37636
rect 29867 37571 29933 37572
rect 28763 35052 28829 35053
rect 28763 34988 28764 35052
rect 28828 34988 28829 35052
rect 28763 34987 28829 34988
rect 28579 34236 28645 34237
rect 28579 34172 28580 34236
rect 28644 34172 28645 34236
rect 28579 34171 28645 34172
rect 26187 33420 26253 33421
rect 26187 33356 26188 33420
rect 26252 33356 26253 33420
rect 26187 33355 26253 33356
rect 25819 30292 25885 30293
rect 25819 30228 25820 30292
rect 25884 30228 25885 30292
rect 25819 30227 25885 30228
rect 25451 26076 25517 26077
rect 25451 26012 25452 26076
rect 25516 26012 25517 26076
rect 25451 26011 25517 26012
rect 25267 19548 25333 19549
rect 25267 19484 25268 19548
rect 25332 19484 25333 19548
rect 25267 19483 25333 19484
rect 26190 19277 26250 33355
rect 28766 30565 28826 34987
rect 29870 32741 29930 37571
rect 33182 36957 33242 39203
rect 34928 38656 35248 39680
rect 40539 38996 40605 38997
rect 40539 38932 40540 38996
rect 40604 38932 40605 38996
rect 40539 38931 40605 38932
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 35387 38180 35453 38181
rect 35387 38116 35388 38180
rect 35452 38116 35453 38180
rect 35387 38115 35453 38116
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 33179 36956 33245 36957
rect 33179 36892 33180 36956
rect 33244 36892 33245 36956
rect 33179 36891 33245 36892
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 32075 35460 32141 35461
rect 32075 35396 32076 35460
rect 32140 35396 32141 35460
rect 32075 35395 32141 35396
rect 32078 34917 32138 35395
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 32075 34916 32141 34917
rect 32075 34852 32076 34916
rect 32140 34852 32141 34916
rect 32075 34851 32141 34852
rect 29867 32740 29933 32741
rect 29867 32676 29868 32740
rect 29932 32676 29933 32740
rect 29867 32675 29933 32676
rect 32078 31381 32138 34851
rect 34099 34644 34165 34645
rect 34099 34580 34100 34644
rect 34164 34580 34165 34644
rect 34099 34579 34165 34580
rect 32443 32332 32509 32333
rect 32443 32268 32444 32332
rect 32508 32268 32509 32332
rect 32443 32267 32509 32268
rect 33731 32332 33797 32333
rect 33731 32268 33732 32332
rect 33796 32268 33797 32332
rect 33731 32267 33797 32268
rect 32075 31380 32141 31381
rect 32075 31316 32076 31380
rect 32140 31316 32141 31380
rect 32075 31315 32141 31316
rect 27843 30564 27909 30565
rect 27843 30500 27844 30564
rect 27908 30500 27909 30564
rect 27843 30499 27909 30500
rect 28763 30564 28829 30565
rect 28763 30500 28764 30564
rect 28828 30500 28829 30564
rect 28763 30499 28829 30500
rect 26739 27708 26805 27709
rect 26739 27644 26740 27708
rect 26804 27644 26805 27708
rect 26739 27643 26805 27644
rect 26187 19276 26253 19277
rect 26187 19212 26188 19276
rect 26252 19212 26253 19276
rect 26187 19211 26253 19212
rect 24531 16828 24597 16829
rect 24531 16764 24532 16828
rect 24596 16764 24597 16828
rect 24531 16763 24597 16764
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 26742 16285 26802 27643
rect 26739 16284 26805 16285
rect 26739 16220 26740 16284
rect 26804 16220 26805 16284
rect 26739 16219 26805 16220
rect 27846 15333 27906 30499
rect 28766 30293 28826 30499
rect 28763 30292 28829 30293
rect 28763 30228 28764 30292
rect 28828 30228 28829 30292
rect 28763 30227 28829 30228
rect 28766 17645 28826 30227
rect 32446 28253 32506 32267
rect 33179 30428 33245 30429
rect 33179 30364 33180 30428
rect 33244 30364 33245 30428
rect 33179 30363 33245 30364
rect 32443 28252 32509 28253
rect 32443 28188 32444 28252
rect 32508 28188 32509 28252
rect 32443 28187 32509 28188
rect 32446 26349 32506 28187
rect 32443 26348 32509 26349
rect 32443 26284 32444 26348
rect 32508 26284 32509 26348
rect 32443 26283 32509 26284
rect 31891 23764 31957 23765
rect 31891 23700 31892 23764
rect 31956 23700 31957 23764
rect 31891 23699 31957 23700
rect 28763 17644 28829 17645
rect 28763 17580 28764 17644
rect 28828 17580 28829 17644
rect 28763 17579 28829 17580
rect 27843 15332 27909 15333
rect 27843 15268 27844 15332
rect 27908 15268 27909 15332
rect 27843 15267 27909 15268
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 31894 12069 31954 23699
rect 33182 23221 33242 30363
rect 33179 23220 33245 23221
rect 33179 23156 33180 23220
rect 33244 23156 33245 23220
rect 33179 23155 33245 23156
rect 32443 22268 32509 22269
rect 32443 22204 32444 22268
rect 32508 22204 32509 22268
rect 32443 22203 32509 22204
rect 31891 12068 31957 12069
rect 31891 12004 31892 12068
rect 31956 12004 31957 12068
rect 31891 12003 31957 12004
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 32446 11389 32506 22203
rect 33734 19413 33794 32267
rect 34102 31925 34162 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 35390 32469 35450 38115
rect 36307 37772 36373 37773
rect 36307 37708 36308 37772
rect 36372 37708 36373 37772
rect 36307 37707 36373 37708
rect 36310 34509 36370 37707
rect 37227 37500 37293 37501
rect 37227 37436 37228 37500
rect 37292 37436 37293 37500
rect 37227 37435 37293 37436
rect 37230 36277 37290 37435
rect 37227 36276 37293 36277
rect 37227 36212 37228 36276
rect 37292 36212 37293 36276
rect 37227 36211 37293 36212
rect 36307 34508 36373 34509
rect 36307 34444 36308 34508
rect 36372 34444 36373 34508
rect 36307 34443 36373 34444
rect 37230 33693 37290 36211
rect 37227 33692 37293 33693
rect 37227 33628 37228 33692
rect 37292 33628 37293 33692
rect 37227 33627 37293 33628
rect 39435 33556 39501 33557
rect 39435 33492 39436 33556
rect 39500 33492 39501 33556
rect 39435 33491 39501 33492
rect 35387 32468 35453 32469
rect 35387 32404 35388 32468
rect 35452 32404 35453 32468
rect 35387 32403 35453 32404
rect 36123 32332 36189 32333
rect 36123 32268 36124 32332
rect 36188 32268 36189 32332
rect 36123 32267 36189 32268
rect 37411 32332 37477 32333
rect 37411 32268 37412 32332
rect 37476 32268 37477 32332
rect 37411 32267 37477 32268
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34099 31924 34165 31925
rect 34099 31860 34100 31924
rect 34164 31860 34165 31924
rect 34099 31859 34165 31860
rect 34099 31652 34165 31653
rect 34099 31588 34100 31652
rect 34164 31588 34165 31652
rect 34099 31587 34165 31588
rect 34102 26213 34162 31587
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34467 29612 34533 29613
rect 34467 29548 34468 29612
rect 34532 29548 34533 29612
rect 34467 29547 34533 29548
rect 34099 26212 34165 26213
rect 34099 26148 34100 26212
rect 34164 26148 34165 26212
rect 34099 26147 34165 26148
rect 34470 24309 34530 29547
rect 34928 28864 35248 29888
rect 35571 29204 35637 29205
rect 35571 29140 35572 29204
rect 35636 29140 35637 29204
rect 35571 29139 35637 29140
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 35387 28524 35453 28525
rect 35387 28460 35388 28524
rect 35452 28460 35453 28524
rect 35387 28459 35453 28460
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 35390 26349 35450 28459
rect 35387 26348 35453 26349
rect 35387 26284 35388 26348
rect 35452 26284 35453 26348
rect 35387 26283 35453 26284
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34467 24308 34533 24309
rect 34467 24244 34468 24308
rect 34532 24244 34533 24308
rect 34467 24243 34533 24244
rect 34928 23424 35248 24448
rect 35574 23765 35634 29139
rect 35939 27708 36005 27709
rect 35939 27644 35940 27708
rect 36004 27644 36005 27708
rect 35939 27643 36005 27644
rect 35942 26077 36002 27643
rect 35939 26076 36005 26077
rect 35939 26012 35940 26076
rect 36004 26012 36005 26076
rect 35939 26011 36005 26012
rect 35571 23764 35637 23765
rect 35571 23700 35572 23764
rect 35636 23700 35637 23764
rect 35571 23699 35637 23700
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 33731 19412 33797 19413
rect 33731 19348 33732 19412
rect 33796 19348 33797 19412
rect 33731 19347 33797 19348
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 36126 15605 36186 32267
rect 37227 32196 37293 32197
rect 37227 32132 37228 32196
rect 37292 32132 37293 32196
rect 37227 32131 37293 32132
rect 37230 28389 37290 32131
rect 37227 28388 37293 28389
rect 37227 28324 37228 28388
rect 37292 28324 37293 28388
rect 37227 28323 37293 28324
rect 37230 27437 37290 28323
rect 37227 27436 37293 27437
rect 37227 27372 37228 27436
rect 37292 27372 37293 27436
rect 37227 27371 37293 27372
rect 37227 26348 37293 26349
rect 37227 26284 37228 26348
rect 37292 26284 37293 26348
rect 37227 26283 37293 26284
rect 37230 22677 37290 26283
rect 37414 25533 37474 32267
rect 39067 29068 39133 29069
rect 39067 29004 39068 29068
rect 39132 29004 39133 29068
rect 39067 29003 39133 29004
rect 39251 29068 39317 29069
rect 39251 29004 39252 29068
rect 39316 29004 39317 29068
rect 39251 29003 39317 29004
rect 38331 27436 38397 27437
rect 38331 27372 38332 27436
rect 38396 27372 38397 27436
rect 38331 27371 38397 27372
rect 37411 25532 37477 25533
rect 37411 25468 37412 25532
rect 37476 25468 37477 25532
rect 37411 25467 37477 25468
rect 37414 24445 37474 25467
rect 37411 24444 37477 24445
rect 37411 24380 37412 24444
rect 37476 24380 37477 24444
rect 37411 24379 37477 24380
rect 37227 22676 37293 22677
rect 37227 22612 37228 22676
rect 37292 22612 37293 22676
rect 37227 22611 37293 22612
rect 36123 15604 36189 15605
rect 36123 15540 36124 15604
rect 36188 15540 36189 15604
rect 36123 15539 36189 15540
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 38334 11933 38394 27371
rect 39070 21997 39130 29003
rect 39067 21996 39133 21997
rect 39067 21932 39068 21996
rect 39132 21932 39133 21996
rect 39067 21931 39133 21932
rect 39254 19005 39314 29003
rect 39438 22813 39498 33491
rect 40355 33284 40421 33285
rect 40355 33220 40356 33284
rect 40420 33220 40421 33284
rect 40355 33219 40421 33220
rect 40358 24445 40418 33219
rect 40542 27709 40602 38931
rect 40907 35596 40973 35597
rect 40907 35532 40908 35596
rect 40972 35532 40973 35596
rect 40907 35531 40973 35532
rect 40910 32061 40970 35531
rect 40907 32060 40973 32061
rect 40907 31996 40908 32060
rect 40972 31996 40973 32060
rect 40907 31995 40973 31996
rect 40539 27708 40605 27709
rect 40539 27644 40540 27708
rect 40604 27644 40605 27708
rect 40539 27643 40605 27644
rect 40355 24444 40421 24445
rect 40355 24380 40356 24444
rect 40420 24380 40421 24444
rect 40355 24379 40421 24380
rect 40910 24173 40970 31995
rect 40907 24172 40973 24173
rect 40907 24108 40908 24172
rect 40972 24108 40973 24172
rect 40907 24107 40973 24108
rect 39435 22812 39501 22813
rect 39435 22748 39436 22812
rect 39500 22748 39501 22812
rect 39435 22747 39501 22748
rect 41275 20772 41341 20773
rect 41275 20708 41276 20772
rect 41340 20708 41341 20772
rect 41275 20707 41341 20708
rect 39251 19004 39317 19005
rect 39251 18940 39252 19004
rect 39316 18940 39317 19004
rect 39251 18939 39317 18940
rect 41278 14109 41338 20707
rect 41275 14108 41341 14109
rect 41275 14044 41276 14108
rect 41340 14044 41341 14108
rect 41275 14043 41341 14044
rect 38331 11932 38397 11933
rect 38331 11868 38332 11932
rect 38396 11868 38397 11932
rect 38331 11867 38397 11868
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 32443 11388 32509 11389
rect 32443 11324 32444 11388
rect 32508 11324 32509 11388
rect 32443 11323 32509 11324
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A0
timestamp 1676037725
transform -1 0 43424 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A0
timestamp 1676037725
transform -1 0 40940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A0
timestamp 1676037725
transform 1 0 41308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 1676037725
transform -1 0 39008 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B
timestamp 1676037725
transform 1 0 36616 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B
timestamp 1676037725
transform 1 0 31464 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1676037725
transform -1 0 43424 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1676037725
transform -1 0 41032 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1676037725
transform 1 0 14996 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1676037725
transform -1 0 38640 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B2
timestamp 1676037725
transform 1 0 28888 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A1
timestamp 1676037725
transform -1 0 43424 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B2
timestamp 1676037725
transform -1 0 37628 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__C1
timestamp 1676037725
transform 1 0 38180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__D
timestamp 1676037725
transform 1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A2
timestamp 1676037725
transform -1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A2
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__B
timestamp 1676037725
transform -1 0 30728 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B2
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A1
timestamp 1676037725
transform 1 0 39376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B
timestamp 1676037725
transform -1 0 34408 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1676037725
transform 1 0 29716 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B2
timestamp 1676037725
transform 1 0 36708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A1
timestamp 1676037725
transform 1 0 36984 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A1
timestamp 1676037725
transform -1 0 42596 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1676037725
transform 1 0 36616 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A2
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B2
timestamp 1676037725
transform 1 0 25944 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A1
timestamp 1676037725
transform 1 0 39284 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1676037725
transform 1 0 33304 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A2
timestamp 1676037725
transform -1 0 23828 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B2
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1676037725
transform 1 0 14720 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B2
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1676037725
transform 1 0 38548 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A1
timestamp 1676037725
transform 1 0 39928 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A1
timestamp 1676037725
transform 1 0 38180 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1676037725
transform 1 0 23828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A
timestamp 1676037725
transform 1 0 35696 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 1676037725
transform -1 0 40480 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1676037725
transform 1 0 36800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__B2
timestamp 1676037725
transform 1 0 25852 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A1
timestamp 1676037725
transform 1 0 39376 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__A1
timestamp 1676037725
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A2
timestamp 1676037725
transform -1 0 26036 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B2
timestamp 1676037725
transform 1 0 24380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1
timestamp 1676037725
transform -1 0 11500 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A1
timestamp 1676037725
transform 1 0 12144 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B
timestamp 1676037725
transform 1 0 31924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A1
timestamp 1676037725
transform 1 0 42964 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1676037725
transform 1 0 33304 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__B2
timestamp 1676037725
transform 1 0 27140 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A
timestamp 1676037725
transform -1 0 15456 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__B2
timestamp 1676037725
transform 1 0 31648 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1676037725
transform 1 0 17204 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A
timestamp 1676037725
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1676037725
transform -1 0 37628 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B
timestamp 1676037725
transform -1 0 42780 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A1
timestamp 1676037725
transform 1 0 35880 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A2
timestamp 1676037725
transform 1 0 37444 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1676037725
transform -1 0 38180 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B
timestamp 1676037725
transform -1 0 42136 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1676037725
transform 1 0 33856 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__B
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__B
timestamp 1676037725
transform -1 0 43424 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__B2
timestamp 1676037725
transform -1 0 43332 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B1
timestamp 1676037725
transform -1 0 38180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1676037725
transform 1 0 26128 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A1
timestamp 1676037725
transform 1 0 38456 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A1
timestamp 1676037725
transform 1 0 23736 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__C1
timestamp 1676037725
transform 1 0 26496 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A1
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__C1
timestamp 1676037725
transform -1 0 26128 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__A1
timestamp 1676037725
transform -1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__C1
timestamp 1676037725
transform -1 0 27968 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1676037725
transform 1 0 32292 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__C1
timestamp 1676037725
transform -1 0 29900 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A
timestamp 1676037725
transform -1 0 42044 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__A1
timestamp 1676037725
transform -1 0 34408 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A
timestamp 1676037725
transform 1 0 38088 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__B
timestamp 1676037725
transform -1 0 38732 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A1
timestamp 1676037725
transform -1 0 42780 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A1
timestamp 1676037725
transform -1 0 41952 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A1
timestamp 1676037725
transform -1 0 39284 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A1
timestamp 1676037725
transform -1 0 17848 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__A1
timestamp 1676037725
transform -1 0 41492 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A1
timestamp 1676037725
transform -1 0 15272 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__A1
timestamp 1676037725
transform -1 0 40204 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A1
timestamp 1676037725
transform -1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__B2
timestamp 1676037725
transform -1 0 15088 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__A1
timestamp 1676037725
transform -1 0 42780 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A1
timestamp 1676037725
transform -1 0 14720 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A1
timestamp 1676037725
transform -1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1676037725
transform -1 0 15824 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A1
timestamp 1676037725
transform -1 0 41400 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__B2
timestamp 1676037725
transform -1 0 43332 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A1
timestamp 1676037725
transform -1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__B2
timestamp 1676037725
transform -1 0 14076 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A1
timestamp 1676037725
transform -1 0 42780 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1676037725
transform -1 0 14628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A1
timestamp 1676037725
transform 1 0 17296 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B2
timestamp 1676037725
transform 1 0 38088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A0
timestamp 1676037725
transform 1 0 41860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A
timestamp 1676037725
transform -1 0 40204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A0
timestamp 1676037725
transform 1 0 40112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A
timestamp 1676037725
transform -1 0 37904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A0
timestamp 1676037725
transform 1 0 41308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A0
timestamp 1676037725
transform -1 0 43424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__A0
timestamp 1676037725
transform -1 0 43424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A1
timestamp 1676037725
transform -1 0 43424 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B1
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A2
timestamp 1676037725
transform 1 0 40204 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__A1
timestamp 1676037725
transform 1 0 34684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__A2
timestamp 1676037725
transform 1 0 36432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1676037725
transform 1 0 36800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A
timestamp 1676037725
transform -1 0 35880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__A
timestamp 1676037725
transform -1 0 41400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1676037725
transform 1 0 41584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__A
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__A
timestamp 1676037725
transform -1 0 33580 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A
timestamp 1676037725
transform 1 0 38180 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__A
timestamp 1676037725
transform 1 0 36800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A
timestamp 1676037725
transform -1 0 38180 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__A
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__D1
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A
timestamp 1676037725
transform 1 0 41676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A
timestamp 1676037725
transform -1 0 35052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__C
timestamp 1676037725
transform -1 0 41308 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__B2
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__A1_N
timestamp 1676037725
transform -1 0 40848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__C
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__A
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__B1
timestamp 1676037725
transform -1 0 43332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__A1
timestamp 1676037725
transform 1 0 39652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__A
timestamp 1676037725
transform -1 0 41584 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__B
timestamp 1676037725
transform 1 0 40756 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__A
timestamp 1676037725
transform -1 0 40388 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__A1
timestamp 1676037725
transform 1 0 41952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__A1
timestamp 1676037725
transform -1 0 20884 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__A2
timestamp 1676037725
transform 1 0 21344 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__B2
timestamp 1676037725
transform 1 0 25668 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__B
timestamp 1676037725
transform -1 0 20976 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__B
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__B2
timestamp 1676037725
transform 1 0 21344 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__C1
timestamp 1676037725
transform 1 0 22172 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__B1
timestamp 1676037725
transform 1 0 21344 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__B2
timestamp 1676037725
transform 1 0 18768 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__B2
timestamp 1676037725
transform 1 0 22080 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__C1
timestamp 1676037725
transform -1 0 22448 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__A1_N
timestamp 1676037725
transform -1 0 19780 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__B1
timestamp 1676037725
transform 1 0 21252 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__B2
timestamp 1676037725
transform 1 0 20792 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__B2
timestamp 1676037725
transform -1 0 21620 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__A1_N
timestamp 1676037725
transform 1 0 18768 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__B1
timestamp 1676037725
transform 1 0 23092 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__B2
timestamp 1676037725
transform 1 0 20240 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__B2
timestamp 1676037725
transform 1 0 20792 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__A1_N
timestamp 1676037725
transform -1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__B1
timestamp 1676037725
transform -1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__B2
timestamp 1676037725
transform 1 0 19872 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__B2
timestamp 1676037725
transform -1 0 27048 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A1_N
timestamp 1676037725
transform 1 0 27140 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__B1
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__B2
timestamp 1676037725
transform 1 0 27692 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__B2
timestamp 1676037725
transform -1 0 28520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__A1_N
timestamp 1676037725
transform -1 0 29164 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__B1
timestamp 1676037725
transform 1 0 29072 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__B2
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__B2
timestamp 1676037725
transform -1 0 29256 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__A1_N
timestamp 1676037725
transform -1 0 32476 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__B1
timestamp 1676037725
transform -1 0 30268 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__B2
timestamp 1676037725
transform 1 0 29532 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1593__A1
timestamp 1676037725
transform -1 0 33304 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__A
timestamp 1676037725
transform -1 0 39836 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__A1
timestamp 1676037725
transform -1 0 20056 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__A2
timestamp 1676037725
transform -1 0 43332 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__A1
timestamp 1676037725
transform -1 0 36800 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A1
timestamp 1676037725
transform -1 0 37628 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A1
timestamp 1676037725
transform -1 0 36248 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__B2
timestamp 1676037725
transform -1 0 33856 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__A2
timestamp 1676037725
transform 1 0 42596 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__A1
timestamp 1676037725
transform 1 0 16928 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__B2
timestamp 1676037725
transform 1 0 17940 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A1
timestamp 1676037725
transform 1 0 17388 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A2
timestamp 1676037725
transform 1 0 18216 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__A1
timestamp 1676037725
transform 1 0 16192 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__B2
timestamp 1676037725
transform 1 0 17112 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1606__A2
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1607__A1
timestamp 1676037725
transform 1 0 17112 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1607__B2
timestamp 1676037725
transform -1 0 41860 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1608__A2
timestamp 1676037725
transform 1 0 16008 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__A1
timestamp 1676037725
transform 1 0 16560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__B2
timestamp 1676037725
transform 1 0 17664 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__A1
timestamp 1676037725
transform 1 0 16836 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__A2
timestamp 1676037725
transform 1 0 17664 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__B2
timestamp 1676037725
transform -1 0 16560 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__A1
timestamp 1676037725
transform 1 0 15456 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__B2
timestamp 1676037725
transform -1 0 15272 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__A2
timestamp 1676037725
transform -1 0 15824 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1613__B
timestamp 1676037725
transform 1 0 30728 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1614__A1
timestamp 1676037725
transform -1 0 34868 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A1
timestamp 1676037725
transform -1 0 39192 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__B1_N
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1617__B2
timestamp 1676037725
transform 1 0 25576 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1621__B2
timestamp 1676037725
transform 1 0 26312 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1624__B2
timestamp 1676037725
transform 1 0 34868 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1625__B
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1627__B2
timestamp 1676037725
transform -1 0 30452 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1628__B2
timestamp 1676037725
transform 1 0 30360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1676037725
transform 1 0 17296 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1630__A2
timestamp 1676037725
transform -1 0 38732 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1630__B1
timestamp 1676037725
transform -1 0 35696 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1632__A1
timestamp 1676037725
transform 1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1634__A2
timestamp 1676037725
transform -1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1635__B
timestamp 1676037725
transform -1 0 29900 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1636__A2
timestamp 1676037725
transform 1 0 32108 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1636__B1
timestamp 1676037725
transform 1 0 30820 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1639__A
timestamp 1676037725
transform -1 0 10488 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A1
timestamp 1676037725
transform -1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B2
timestamp 1676037725
transform 1 0 27324 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1642__A2_N
timestamp 1676037725
transform 1 0 29808 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__A2_N
timestamp 1676037725
transform -1 0 27876 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__B2
timestamp 1676037725
transform 1 0 29716 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__A
timestamp 1676037725
transform -1 0 41584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1647__A
timestamp 1676037725
transform 1 0 41308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1648__A
timestamp 1676037725
transform 1 0 41032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1649__A
timestamp 1676037725
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1650__A
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1651__A
timestamp 1676037725
transform -1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1653__A0
timestamp 1676037725
transform -1 0 24196 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1653__A1
timestamp 1676037725
transform 1 0 23460 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1658__S
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1663__A
timestamp 1676037725
transform -1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1664__B1
timestamp 1676037725
transform 1 0 20148 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1666__A1
timestamp 1676037725
transform 1 0 23644 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1667__S
timestamp 1676037725
transform -1 0 24012 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1669__A
timestamp 1676037725
transform 1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1670__A
timestamp 1676037725
transform -1 0 19596 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1673__B1
timestamp 1676037725
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1674__S
timestamp 1676037725
transform -1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1677__A
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1679__A1
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1680__S
timestamp 1676037725
transform -1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1682__A0
timestamp 1676037725
transform 1 0 20332 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1682__A1
timestamp 1676037725
transform 1 0 19504 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1683__S
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1685__A
timestamp 1676037725
transform 1 0 21620 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1686__A
timestamp 1676037725
transform 1 0 21344 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__B1
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__A
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1690__A1
timestamp 1676037725
transform 1 0 25852 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1691__S
timestamp 1676037725
transform 1 0 13616 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__A
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1694__A
timestamp 1676037725
transform 1 0 23000 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1697__B1
timestamp 1676037725
transform 1 0 25760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1698__S
timestamp 1676037725
transform -1 0 17020 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1701__A
timestamp 1676037725
transform 1 0 20884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1704__A1
timestamp 1676037725
transform 1 0 28244 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1704__A2
timestamp 1676037725
transform 1 0 29072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1704__A3
timestamp 1676037725
transform -1 0 27324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1705__A1
timestamp 1676037725
transform -1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1705__S
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1723__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1728__A
timestamp 1676037725
transform -1 0 40296 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1729__B
timestamp 1676037725
transform 1 0 36248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1735__B
timestamp 1676037725
transform -1 0 42780 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1738__S
timestamp 1676037725
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1740__S
timestamp 1676037725
transform -1 0 18400 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1742__S
timestamp 1676037725
transform 1 0 18768 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1744__S
timestamp 1676037725
transform 1 0 20148 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__S
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1748__S
timestamp 1676037725
transform -1 0 24104 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1750__S
timestamp 1676037725
transform -1 0 23552 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1752__S
timestamp 1676037725
transform -1 0 22172 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1755__A1
timestamp 1676037725
transform -1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1757__A1
timestamp 1676037725
transform 1 0 29808 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1758__A0
timestamp 1676037725
transform 1 0 31648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1761__A2_N
timestamp 1676037725
transform 1 0 32476 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1761__B1
timestamp 1676037725
transform -1 0 33212 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__A
timestamp 1676037725
transform 1 0 30452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__B
timestamp 1676037725
transform 1 0 25576 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__C
timestamp 1676037725
transform 1 0 24932 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__D
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__A
timestamp 1676037725
transform 1 0 26772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__B
timestamp 1676037725
transform 1 0 26036 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__C
timestamp 1676037725
transform 1 0 26220 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__D
timestamp 1676037725
transform 1 0 25668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__A0
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__A1
timestamp 1676037725
transform 1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1770__B1_N
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1777__A0
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1777__A1
timestamp 1676037725
transform 1 0 29072 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1778__B1
timestamp 1676037725
transform 1 0 28520 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1779__A1
timestamp 1676037725
transform 1 0 27968 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1783__A1
timestamp 1676037725
transform 1 0 26404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1784__A0
timestamp 1676037725
transform 1 0 26496 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1785__A
timestamp 1676037725
transform 1 0 34592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1787__A1
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1791__A0
timestamp 1676037725
transform 1 0 31648 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1792__A0
timestamp 1676037725
transform 1 0 33396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1794__A2
timestamp 1676037725
transform 1 0 35144 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1796__A
timestamp 1676037725
transform 1 0 31188 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__A
timestamp 1676037725
transform 1 0 20700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__B
timestamp 1676037725
transform 1 0 20148 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__A2
timestamp 1676037725
transform 1 0 26404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__C1
timestamp 1676037725
transform 1 0 28060 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__A1
timestamp 1676037725
transform 1 0 28244 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__A2
timestamp 1676037725
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1804__A4
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1807__A
timestamp 1676037725
transform 1 0 41952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1807__B
timestamp 1676037725
transform -1 0 41952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1809__A0
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__A0
timestamp 1676037725
transform 1 0 41860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1813__A0
timestamp 1676037725
transform -1 0 42872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1815__A0
timestamp 1676037725
transform -1 0 42872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A0
timestamp 1676037725
transform -1 0 42228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1819__A0
timestamp 1676037725
transform -1 0 41768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1821__A0
timestamp 1676037725
transform -1 0 43424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1823__A0
timestamp 1676037725
transform 1 0 32016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1825__A
timestamp 1676037725
transform 1 0 42320 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1827__A1
timestamp 1676037725
transform -1 0 43240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1827__B1
timestamp 1676037725
transform 1 0 41952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1845__A
timestamp 1676037725
transform 1 0 26496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__A
timestamp 1676037725
transform -1 0 40756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__A2
timestamp 1676037725
transform -1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__B1
timestamp 1676037725
transform 1 0 21344 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__B1
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1874__S
timestamp 1676037725
transform 1 0 35052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__A0
timestamp 1676037725
transform -1 0 35788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__S
timestamp 1676037725
transform 1 0 33856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1879__B
timestamp 1676037725
transform 1 0 31648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1881__A0
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1881__S
timestamp 1676037725
transform 1 0 29072 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1885__A2
timestamp 1676037725
transform 1 0 30728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1889__B
timestamp 1676037725
transform 1 0 31096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1890__A2
timestamp 1676037725
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1895__A2
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1897__S
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1899__A2
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1900__C
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1910__S
timestamp 1676037725
transform 1 0 26496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1914__A2
timestamp 1676037725
transform 1 0 27508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1915__S
timestamp 1676037725
transform 1 0 28520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1918__B2
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1921__A2
timestamp 1676037725
transform 1 0 36064 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1923__A2
timestamp 1676037725
transform 1 0 30636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__A2
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1928__A1
timestamp 1676037725
transform -1 0 35880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1931__A2
timestamp 1676037725
transform -1 0 42044 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1932__S
timestamp 1676037725
transform -1 0 43332 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1934__S
timestamp 1676037725
transform -1 0 40756 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1944__A0
timestamp 1676037725
transform 1 0 18768 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1950__S
timestamp 1676037725
transform -1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1952__S
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1954__S
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1956__S
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1958__S
timestamp 1676037725
transform 1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1960__S
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1962__S
timestamp 1676037725
transform -1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1964__A1
timestamp 1676037725
transform -1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1964__S
timestamp 1676037725
transform -1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1982__A1
timestamp 1676037725
transform -1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1988__CLK
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1989__CLK
timestamp 1676037725
transform 1 0 22264 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2018__CLK
timestamp 1676037725
transform -1 0 31556 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2022__CLK
timestamp 1676037725
transform -1 0 24840 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2025__CLK
timestamp 1676037725
transform 1 0 39284 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2041__CLK
timestamp 1676037725
transform -1 0 41308 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2042__CLK
timestamp 1676037725
transform -1 0 29440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2044__CLK
timestamp 1676037725
transform 1 0 26404 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2044__D
timestamp 1676037725
transform 1 0 30176 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2045__CLK
timestamp 1676037725
transform -1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2046__CLK
timestamp 1676037725
transform -1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2048__CLK
timestamp 1676037725
transform 1 0 36340 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2071__CLK
timestamp 1676037725
transform -1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2075__CLK
timestamp 1676037725
transform -1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2090__CLK
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2093__CLK
timestamp 1676037725
transform -1 0 12788 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2094__CLK
timestamp 1676037725
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2095__CLK
timestamp 1676037725
transform -1 0 19780 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2096__CLK
timestamp 1676037725
transform -1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1676037725
transform -1 0 33028 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1676037725
transform 1 0 23828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1676037725
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1676037725
transform 1 0 31464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1676037725
transform 1 0 30084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1676037725
transform 1 0 33488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1676037725
transform 1 0 23184 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1676037725
transform 1 0 27140 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1676037725
transform 1 0 26496 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1676037725
transform 1 0 30912 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1676037725
transform 1 0 39284 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1676037725
transform -1 0 39284 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1676037725
transform -1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1676037725
transform 1 0 37444 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform -1 0 43424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 43424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 43424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 42872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 42780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 43424 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 43424 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform -1 0 18216 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform -1 0 14168 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform -1 0 20056 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_453
timestamp 1676037725
transform 1 0 42780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_460 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43424 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_449 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_457
timestamp 1676037725
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_460
timestamp 1676037725
transform 1 0 43424 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_461
timestamp 1676037725
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_461
timestamp 1676037725
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_460
timestamp 1676037725
transform 1 0 43424 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_453
timestamp 1676037725
transform 1 0 42780 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_460
timestamp 1676037725
transform 1 0 43424 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_461
timestamp 1676037725
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_460
timestamp 1676037725
transform 1 0 43424 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_454
timestamp 1676037725
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_460
timestamp 1676037725
transform 1 0 43424 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_451
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_454
timestamp 1676037725
transform 1 0 42872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_460
timestamp 1676037725
transform 1 0 43424 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_423
timestamp 1676037725
transform 1 0 40020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_426
timestamp 1676037725
transform 1 0 40296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_430
timestamp 1676037725
transform 1 0 40664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_433
timestamp 1676037725
transform 1 0 40940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_439
timestamp 1676037725
transform 1 0 41492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_442
timestamp 1676037725
transform 1 0 41768 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_454
timestamp 1676037725
transform 1 0 42872 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_460
timestamp 1676037725
transform 1 0 43424 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_317
timestamp 1676037725
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_326
timestamp 1676037725
transform 1 0 31096 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_350
timestamp 1676037725
transform 1 0 33304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_397
timestamp 1676037725
transform 1 0 37628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_400
timestamp 1676037725
transform 1 0 37904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_412
timestamp 1676037725
transform 1 0 39008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 1676037725
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_425
timestamp 1676037725
transform 1 0 40204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_429
timestamp 1676037725
transform 1 0 40572 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_439
timestamp 1676037725
transform 1 0 41492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_447
timestamp 1676037725
transform 1 0 42228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_453
timestamp 1676037725
transform 1 0 42780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_460
timestamp 1676037725
transform 1 0 43424 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_314
timestamp 1676037725
transform 1 0 29992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_348
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_358
timestamp 1676037725
transform 1 0 34040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_371
timestamp 1676037725
transform 1 0 35236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_377
timestamp 1676037725
transform 1 0 35788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_403
timestamp 1676037725
transform 1 0 38180 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_425
timestamp 1676037725
transform 1 0 40204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1676037725
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_453
timestamp 1676037725
transform 1 0 42780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_457
timestamp 1676037725
transform 1 0 43148 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_460
timestamp 1676037725
transform 1 0 43424 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_287
timestamp 1676037725
transform 1 0 27508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_327
timestamp 1676037725
transform 1 0 31188 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_335
timestamp 1676037725
transform 1 0 31924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_354
timestamp 1676037725
transform 1 0 33672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_358
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_369
timestamp 1676037725
transform 1 0 35052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_386
timestamp 1676037725
transform 1 0 36616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_393
timestamp 1676037725
transform 1 0 37260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_405
timestamp 1676037725
transform 1 0 38364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_443
timestamp 1676037725
transform 1 0 41860 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_447
timestamp 1676037725
transform 1 0 42228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_461
timestamp 1676037725
transform 1 0 43516 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1676037725
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_312
timestamp 1676037725
transform 1 0 29808 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_327
timestamp 1676037725
transform 1 0 31188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1676037725
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_358
timestamp 1676037725
transform 1 0 34040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_369
timestamp 1676037725
transform 1 0 35052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_379
timestamp 1676037725
transform 1 0 35972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_400
timestamp 1676037725
transform 1 0 37904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_409
timestamp 1676037725
transform 1 0 38732 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_424
timestamp 1676037725
transform 1 0 40112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_437
timestamp 1676037725
transform 1 0 41308 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1676037725
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_460
timestamp 1676037725
transform 1 0 43424 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_229
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_235
timestamp 1676037725
transform 1 0 22724 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1676037725
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_300
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1676037725
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_325
timestamp 1676037725
transform 1 0 31004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_344
timestamp 1676037725
transform 1 0 32752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_352
timestamp 1676037725
transform 1 0 33488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1676037725
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_372
timestamp 1676037725
transform 1 0 35328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_378
timestamp 1676037725
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_396
timestamp 1676037725
transform 1 0 37536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_410
timestamp 1676037725
transform 1 0 38824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1676037725
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_425
timestamp 1676037725
transform 1 0 40204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_431
timestamp 1676037725
transform 1 0 40756 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_437
timestamp 1676037725
transform 1 0 41308 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_440
timestamp 1676037725
transform 1 0 41584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_460
timestamp 1676037725
transform 1 0 43424 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_216
timestamp 1676037725
transform 1 0 20976 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_255
timestamp 1676037725
transform 1 0 24564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_269
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_275
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_286
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_294
timestamp 1676037725
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_313
timestamp 1676037725
transform 1 0 29900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_327
timestamp 1676037725
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_347
timestamp 1676037725
transform 1 0 33028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_356
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_366
timestamp 1676037725
transform 1 0 34776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_372
timestamp 1676037725
transform 1 0 35328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_378
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_404
timestamp 1676037725
transform 1 0 38272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_413
timestamp 1676037725
transform 1 0 39100 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_421
timestamp 1676037725
transform 1 0 39836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_431
timestamp 1676037725
transform 1 0 40756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_439
timestamp 1676037725
transform 1 0 41492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1676037725
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_460
timestamp 1676037725
transform 1 0 43424 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_175
timestamp 1676037725
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_202
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_271
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_287
timestamp 1676037725
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_293
timestamp 1676037725
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1676037725
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1676037725
transform 1 0 31372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_340
timestamp 1676037725
transform 1 0 32384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_371
timestamp 1676037725
transform 1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_375
timestamp 1676037725
transform 1 0 35604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_383
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_396
timestamp 1676037725
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_410
timestamp 1676037725
transform 1 0 38824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_414
timestamp 1676037725
transform 1 0 39192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_439
timestamp 1676037725
transform 1 0 41492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_459
timestamp 1676037725
transform 1 0 43332 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1676037725
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_162
timestamp 1676037725
transform 1 0 16008 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1676037725
transform 1 0 18032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_204
timestamp 1676037725
transform 1 0 19872 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_241
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_267
timestamp 1676037725
transform 1 0 25668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1676037725
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1676037725
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_321
timestamp 1676037725
transform 1 0 30636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_344
timestamp 1676037725
transform 1 0 32752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_348
timestamp 1676037725
transform 1 0 33120 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_354
timestamp 1676037725
transform 1 0 33672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1676037725
transform 1 0 34408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_368
timestamp 1676037725
transform 1 0 34960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_375
timestamp 1676037725
transform 1 0 35604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_383
timestamp 1676037725
transform 1 0 36340 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_387
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_406
timestamp 1676037725
transform 1 0 38456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_413
timestamp 1676037725
transform 1 0 39100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_427
timestamp 1676037725
transform 1 0 40388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_440
timestamp 1676037725
transform 1 0 41584 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_446
timestamp 1676037725
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_460
timestamp 1676037725
transform 1 0 43424 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1676037725
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_190
timestamp 1676037725
transform 1 0 18584 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_227
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_232
timestamp 1676037725
transform 1 0 22448 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1676037725
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_263
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_285
timestamp 1676037725
transform 1 0 27324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_297
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_318
timestamp 1676037725
transform 1 0 30360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_324
timestamp 1676037725
transform 1 0 30912 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_337
timestamp 1676037725
transform 1 0 32108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1676037725
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp 1676037725
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1676037725
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_372
timestamp 1676037725
transform 1 0 35328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_384
timestamp 1676037725
transform 1 0 36432 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_393
timestamp 1676037725
transform 1 0 37260 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_397
timestamp 1676037725
transform 1 0 37628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_402
timestamp 1676037725
transform 1 0 38088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_409
timestamp 1676037725
transform 1 0 38732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_432
timestamp 1676037725
transform 1 0 40848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_438
timestamp 1676037725
transform 1 0 41400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_444
timestamp 1676037725
transform 1 0 41952 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_450
timestamp 1676037725
transform 1 0 42504 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_460
timestamp 1676037725
transform 1 0 43424 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1676037725
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1676037725
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_249
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1676037725
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_294
timestamp 1676037725
transform 1 0 28152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_304
timestamp 1676037725
transform 1 0 29072 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1676037725
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1676037725
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_341
timestamp 1676037725
transform 1 0 32476 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_347
timestamp 1676037725
transform 1 0 33028 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_355
timestamp 1676037725
transform 1 0 33764 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_371
timestamp 1676037725
transform 1 0 35236 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1676037725
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_400
timestamp 1676037725
transform 1 0 37904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_409
timestamp 1676037725
transform 1 0 38732 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_415
timestamp 1676037725
transform 1 0 39284 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_421
timestamp 1676037725
transform 1 0 39836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_440
timestamp 1676037725
transform 1 0 41584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_454
timestamp 1676037725
transform 1 0 42872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_460
timestamp 1676037725
transform 1 0 43424 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_175
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_181
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1676037725
transform 1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1676037725
transform 1 0 20424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1676037725
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_272
timestamp 1676037725
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_278
timestamp 1676037725
transform 1 0 26680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1676037725
transform 1 0 27600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1676037725
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1676037725
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_322
timestamp 1676037725
transform 1 0 30728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1676037725
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_334
timestamp 1676037725
transform 1 0 31832 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_340
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_348
timestamp 1676037725
transform 1 0 33120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_355
timestamp 1676037725
transform 1 0 33764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1676037725
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_372
timestamp 1676037725
transform 1 0 35328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_378
timestamp 1676037725
transform 1 0 35880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_382
timestamp 1676037725
transform 1 0 36248 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_390
timestamp 1676037725
transform 1 0 36984 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_396
timestamp 1676037725
transform 1 0 37536 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_404
timestamp 1676037725
transform 1 0 38272 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1676037725
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_427
timestamp 1676037725
transform 1 0 40388 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_437
timestamp 1676037725
transform 1 0 41308 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_443
timestamp 1676037725
transform 1 0 41860 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_460
timestamp 1676037725
transform 1 0 43424 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_156
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_173
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1676037725
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1676037725
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_255
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_294
timestamp 1676037725
transform 1 0 28152 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_300
timestamp 1676037725
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1676037725
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_308
timestamp 1676037725
transform 1 0 29440 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_325
timestamp 1676037725
transform 1 0 31004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_344
timestamp 1676037725
transform 1 0 32752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_352
timestamp 1676037725
transform 1 0 33488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_365
timestamp 1676037725
transform 1 0 34684 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_375
timestamp 1676037725
transform 1 0 35604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_384
timestamp 1676037725
transform 1 0 36432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_397
timestamp 1676037725
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1676037725
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_409
timestamp 1676037725
transform 1 0 38732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_419
timestamp 1676037725
transform 1 0 39652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_425
timestamp 1676037725
transform 1 0 40204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1676037725
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_460
timestamp 1676037725
transform 1 0 43424 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_152
timestamp 1676037725
transform 1 0 15088 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1676037725
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1676037725
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1676037725
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_211
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_218
timestamp 1676037725
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_225
timestamp 1676037725
transform 1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_238
timestamp 1676037725
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_281
timestamp 1676037725
transform 1 0 26956 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_294
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1676037725
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1676037725
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_323
timestamp 1676037725
transform 1 0 30820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_336
timestamp 1676037725
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1676037725
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1676037725
transform 1 0 35420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_383
timestamp 1676037725
transform 1 0 36340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_396
timestamp 1676037725
transform 1 0 37536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_406
timestamp 1676037725
transform 1 0 38456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_415
timestamp 1676037725
transform 1 0 39284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_429
timestamp 1676037725
transform 1 0 40572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_443
timestamp 1676037725
transform 1 0 41860 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_456
timestamp 1676037725
transform 1 0 43056 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1676037725
transform 1 0 13064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_187
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_195
timestamp 1676037725
transform 1 0 19044 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_212
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_299
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_307
timestamp 1676037725
transform 1 0 29348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_311
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_323
timestamp 1676037725
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_327
timestamp 1676037725
transform 1 0 31188 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_355
timestamp 1676037725
transform 1 0 33764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_365
timestamp 1676037725
transform 1 0 34684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_369
timestamp 1676037725
transform 1 0 35052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_401
timestamp 1676037725
transform 1 0 37996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_407
timestamp 1676037725
transform 1 0 38548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_414
timestamp 1676037725
transform 1 0 39192 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_425
timestamp 1676037725
transform 1 0 40204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_433
timestamp 1676037725
transform 1 0 40940 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_436
timestamp 1676037725
transform 1 0 41216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_460
timestamp 1676037725
transform 1 0 43424 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_207
timestamp 1676037725
transform 1 0 20148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_220
timestamp 1676037725
transform 1 0 21344 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_226
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_231
timestamp 1676037725
transform 1 0 22356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1676037725
transform 1 0 23184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_283
timestamp 1676037725
transform 1 0 27140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1676037725
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_319
timestamp 1676037725
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_326
timestamp 1676037725
transform 1 0 31096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1676037725
transform 1 0 31648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_338
timestamp 1676037725
transform 1 0 32200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_348
timestamp 1676037725
transform 1 0 33120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_354
timestamp 1676037725
transform 1 0 33672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_358
timestamp 1676037725
transform 1 0 34040 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_372
timestamp 1676037725
transform 1 0 35328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_378
timestamp 1676037725
transform 1 0 35880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_391
timestamp 1676037725
transform 1 0 37076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_404
timestamp 1676037725
transform 1 0 38272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1676037725
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_427
timestamp 1676037725
transform 1 0 40388 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_439
timestamp 1676037725
transform 1 0 41492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_443
timestamp 1676037725
transform 1 0 41860 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_460
timestamp 1676037725
transform 1 0 43424 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_202
timestamp 1676037725
transform 1 0 19688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1676037725
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_250
timestamp 1676037725
transform 1 0 24104 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1676037725
transform 1 0 24840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_289
timestamp 1676037725
transform 1 0 27692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_304
timestamp 1676037725
transform 1 0 29072 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1676037725
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_346
timestamp 1676037725
transform 1 0 32936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1676037725
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_365
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_371
timestamp 1676037725
transform 1 0 35236 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_384
timestamp 1676037725
transform 1 0 36432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1676037725
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_415
timestamp 1676037725
transform 1 0 39284 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_424
timestamp 1676037725
transform 1 0 40112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_428
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1676037725
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_460
timestamp 1676037725
transform 1 0 43424 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_149
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_154
timestamp 1676037725
transform 1 0 15272 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1676037725
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1676037725
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1676037725
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_234
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_257
timestamp 1676037725
transform 1 0 24748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_269
timestamp 1676037725
transform 1 0 25852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1676037725
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_327
timestamp 1676037725
transform 1 0 31188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_331
timestamp 1676037725
transform 1 0 31556 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_348
timestamp 1676037725
transform 1 0 33120 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1676037725
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_369
timestamp 1676037725
transform 1 0 35052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_376
timestamp 1676037725
transform 1 0 35696 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_384
timestamp 1676037725
transform 1 0 36432 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_390
timestamp 1676037725
transform 1 0 36984 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_397
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_403
timestamp 1676037725
transform 1 0 38180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1676037725
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_427
timestamp 1676037725
transform 1 0 40388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_436
timestamp 1676037725
transform 1 0 41216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_442
timestamp 1676037725
transform 1 0 41768 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_448
timestamp 1676037725
transform 1 0 42320 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_452
timestamp 1676037725
transform 1 0 42688 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_458
timestamp 1676037725
transform 1 0 43240 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_257
timestamp 1676037725
transform 1 0 24748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_299
timestamp 1676037725
transform 1 0 28612 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_314
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_323
timestamp 1676037725
transform 1 0 30820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_351
timestamp 1676037725
transform 1 0 33396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_372
timestamp 1676037725
transform 1 0 35328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_376
timestamp 1676037725
transform 1 0 35696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_381
timestamp 1676037725
transform 1 0 36156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1676037725
transform 1 0 37904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_409
timestamp 1676037725
transform 1 0 38732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_424
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_434
timestamp 1676037725
transform 1 0 41032 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1676037725
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_453
timestamp 1676037725
transform 1 0 42780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_459
timestamp 1676037725
transform 1 0 43332 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1676037725
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1676037725
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_270
timestamp 1676037725
transform 1 0 25944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_278
timestamp 1676037725
transform 1 0 26680 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_285
timestamp 1676037725
transform 1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1676037725
transform 1 0 28336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1676037725
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_313
timestamp 1676037725
transform 1 0 29900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_317
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_325
timestamp 1676037725
transform 1 0 31004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_349
timestamp 1676037725
transform 1 0 33212 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_355
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1676037725
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_387
timestamp 1676037725
transform 1 0 36708 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_395
timestamp 1676037725
transform 1 0 37444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_403
timestamp 1676037725
transform 1 0 38180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1676037725
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_426
timestamp 1676037725
transform 1 0 40296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_432
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_438
timestamp 1676037725
transform 1 0 41400 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_460
timestamp 1676037725
transform 1 0 43424 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_132
timestamp 1676037725
transform 1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1676037725
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_202
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1676037725
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1676037725
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1676037725
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1676037725
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_290
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_308
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_327
timestamp 1676037725
transform 1 0 31188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_331
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_346
timestamp 1676037725
transform 1 0 32936 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_352
timestamp 1676037725
transform 1 0 33488 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_369
timestamp 1676037725
transform 1 0 35052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_380
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_402
timestamp 1676037725
transform 1 0 38088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_416
timestamp 1676037725
transform 1 0 39376 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_424
timestamp 1676037725
transform 1 0 40112 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1676037725
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_456
timestamp 1676037725
transform 1 0 43056 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1676037725
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_180
timestamp 1676037725
transform 1 0 17664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_220
timestamp 1676037725
transform 1 0 21344 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1676037725
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1676037725
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_300
timestamp 1676037725
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1676037725
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_331
timestamp 1676037725
transform 1 0 31556 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_339
timestamp 1676037725
transform 1 0 32292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_348
timestamp 1676037725
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_354
timestamp 1676037725
transform 1 0 33672 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_376
timestamp 1676037725
transform 1 0 35696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1676037725
transform 1 0 36248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_386
timestamp 1676037725
transform 1 0 36616 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_392
timestamp 1676037725
transform 1 0 37168 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_402
timestamp 1676037725
transform 1 0 38088 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_408
timestamp 1676037725
transform 1 0 38640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1676037725
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_431
timestamp 1676037725
transform 1 0 40756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_437
timestamp 1676037725
transform 1 0 41308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_443
timestamp 1676037725
transform 1 0 41860 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_449
timestamp 1676037725
transform 1 0 42412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_453
timestamp 1676037725
transform 1 0 42780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_460
timestamp 1676037725
transform 1 0 43424 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_162
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1676037725
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_259
timestamp 1676037725
transform 1 0 24932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_314
timestamp 1676037725
transform 1 0 29992 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_324
timestamp 1676037725
transform 1 0 30912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_360
timestamp 1676037725
transform 1 0 34224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_364
timestamp 1676037725
transform 1 0 34592 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_367
timestamp 1676037725
transform 1 0 34868 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_380
timestamp 1676037725
transform 1 0 36064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1676037725
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_401
timestamp 1676037725
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_410
timestamp 1676037725
transform 1 0 38824 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_422
timestamp 1676037725
transform 1 0 39928 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_454
timestamp 1676037725
transform 1 0 42872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_460
timestamp 1676037725
transform 1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1676037725
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_156
timestamp 1676037725
transform 1 0 15456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_181
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_220
timestamp 1676037725
transform 1 0 21344 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1676037725
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_235
timestamp 1676037725
transform 1 0 22724 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_271
timestamp 1676037725
transform 1 0 26036 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1676037725
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_326
timestamp 1676037725
transform 1 0 31096 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_352
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_358
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_373
timestamp 1676037725
transform 1 0 35420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_390
timestamp 1676037725
transform 1 0 36984 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_396
timestamp 1676037725
transform 1 0 37536 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1676037725
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_410
timestamp 1676037725
transform 1 0 38824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1676037725
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_426
timestamp 1676037725
transform 1 0 40296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_437
timestamp 1676037725
transform 1 0 41308 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_459
timestamp 1676037725
transform 1 0 43332 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_131
timestamp 1676037725
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_156
timestamp 1676037725
transform 1 0 15456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1676037725
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_199
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1676037725
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1676037725
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_229
timestamp 1676037725
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_239
timestamp 1676037725
transform 1 0 23092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1676037725
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_251
timestamp 1676037725
transform 1 0 24196 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_271
timestamp 1676037725
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_275
timestamp 1676037725
transform 1 0 26404 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_285
timestamp 1676037725
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_291
timestamp 1676037725
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_297
timestamp 1676037725
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_308
timestamp 1676037725
transform 1 0 29440 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_314
timestamp 1676037725
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_327
timestamp 1676037725
transform 1 0 31188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_346
timestamp 1676037725
transform 1 0 32936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_360
timestamp 1676037725
transform 1 0 34224 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_366
timestamp 1676037725
transform 1 0 34776 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_381
timestamp 1676037725
transform 1 0 36156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1676037725
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_398
timestamp 1676037725
transform 1 0 37720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_404
timestamp 1676037725
transform 1 0 38272 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1676037725
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_421
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_427
timestamp 1676037725
transform 1 0 40388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_431
timestamp 1676037725
transform 1 0 40756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_435
timestamp 1676037725
transform 1 0 41124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1676037725
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_459
timestamp 1676037725
transform 1 0 43332 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1676037725
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1676037725
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1676037725
transform 1 0 15824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_164
timestamp 1676037725
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1676037725
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1676037725
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_217
timestamp 1676037725
transform 1 0 21068 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_227
timestamp 1676037725
transform 1 0 21988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_263
timestamp 1676037725
transform 1 0 25300 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_269
timestamp 1676037725
transform 1 0 25852 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_279
timestamp 1676037725
transform 1 0 26772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1676037725
transform 1 0 28244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_299
timestamp 1676037725
transform 1 0 28612 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1676037725
transform 1 0 31188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1676037725
transform 1 0 32660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1676037725
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1676037725
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_373
timestamp 1676037725
transform 1 0 35420 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_379
timestamp 1676037725
transform 1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_387
timestamp 1676037725
transform 1 0 36708 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_394
timestamp 1676037725
transform 1 0 37352 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_406
timestamp 1676037725
transform 1 0 38456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1676037725
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_429
timestamp 1676037725
transform 1 0 40572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_435
timestamp 1676037725
transform 1 0 41124 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_449
timestamp 1676037725
transform 1 0 42412 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_456
timestamp 1676037725
transform 1 0 43056 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_133
timestamp 1676037725
transform 1 0 13340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_150
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1676037725
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_177
timestamp 1676037725
transform 1 0 17388 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_201
timestamp 1676037725
transform 1 0 19596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_209
timestamp 1676037725
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_218
timestamp 1676037725
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_234
timestamp 1676037725
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_241
timestamp 1676037725
transform 1 0 23276 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_247
timestamp 1676037725
transform 1 0 23828 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_292
timestamp 1676037725
transform 1 0 27968 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_328
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_343
timestamp 1676037725
transform 1 0 32660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_351
timestamp 1676037725
transform 1 0 33396 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_356
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_363
timestamp 1676037725
transform 1 0 34500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_372
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_384
timestamp 1676037725
transform 1 0 36432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_403
timestamp 1676037725
transform 1 0 38180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_411
timestamp 1676037725
transform 1 0 38916 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_420
timestamp 1676037725
transform 1 0 39744 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_428
timestamp 1676037725
transform 1 0 40480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_433
timestamp 1676037725
transform 1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_457
timestamp 1676037725
transform 1 0 43148 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1676037725
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_158
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1676037725
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_178
timestamp 1676037725
transform 1 0 17480 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_204
timestamp 1676037725
transform 1 0 19872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_216
timestamp 1676037725
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_227
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_234
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_240
timestamp 1676037725
transform 1 0 23184 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_262
timestamp 1676037725
transform 1 0 25208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_270
timestamp 1676037725
transform 1 0 25944 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1676037725
transform 1 0 26496 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1676037725
transform 1 0 27324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_296
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_320
timestamp 1676037725
transform 1 0 30544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_332
timestamp 1676037725
transform 1 0 31648 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_336
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_341
timestamp 1676037725
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_347
timestamp 1676037725
transform 1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_351
timestamp 1676037725
transform 1 0 33396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_374
timestamp 1676037725
transform 1 0 35512 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_382
timestamp 1676037725
transform 1 0 36248 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_388
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_407
timestamp 1676037725
transform 1 0 38548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1676037725
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_428
timestamp 1676037725
transform 1 0 40480 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_434
timestamp 1676037725
transform 1 0 41032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_439
timestamp 1676037725
transform 1 0 41492 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_447
timestamp 1676037725
transform 1 0 42228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_453
timestamp 1676037725
transform 1 0 42780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_460
timestamp 1676037725
transform 1 0 43424 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_131
timestamp 1676037725
transform 1 0 13156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_151
timestamp 1676037725
transform 1 0 14996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_191
timestamp 1676037725
transform 1 0 18676 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1676037725
transform 1 0 20240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1676037725
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_232
timestamp 1676037725
transform 1 0 22448 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_241
timestamp 1676037725
transform 1 0 23276 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_253
timestamp 1676037725
transform 1 0 24380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1676037725
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_274
timestamp 1676037725
transform 1 0 26312 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1676037725
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_285
timestamp 1676037725
transform 1 0 27324 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_289
timestamp 1676037725
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_306
timestamp 1676037725
transform 1 0 29256 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_310
timestamp 1676037725
transform 1 0 29624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_318
timestamp 1676037725
transform 1 0 30360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_325
timestamp 1676037725
transform 1 0 31004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1676037725
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_347
timestamp 1676037725
transform 1 0 33028 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_353
timestamp 1676037725
transform 1 0 33580 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_357
timestamp 1676037725
transform 1 0 33948 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_366
timestamp 1676037725
transform 1 0 34776 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_372
timestamp 1676037725
transform 1 0 35328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_380
timestamp 1676037725
transform 1 0 36064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_401
timestamp 1676037725
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_408
timestamp 1676037725
transform 1 0 38640 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_412
timestamp 1676037725
transform 1 0 39008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_420
timestamp 1676037725
transform 1 0 39744 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_427
timestamp 1676037725
transform 1 0 40388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_434
timestamp 1676037725
transform 1 0 41032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1676037725
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_459
timestamp 1676037725
transform 1 0 43332 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_146
timestamp 1676037725
transform 1 0 14536 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_170
timestamp 1676037725
transform 1 0 16744 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_181
timestamp 1676037725
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1676037725
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_203
timestamp 1676037725
transform 1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_218
timestamp 1676037725
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_222
timestamp 1676037725
transform 1 0 21528 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_231
timestamp 1676037725
transform 1 0 22356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_240
timestamp 1676037725
transform 1 0 23184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_244
timestamp 1676037725
transform 1 0 23552 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1676037725
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1676037725
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_275
timestamp 1676037725
transform 1 0 26404 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_281
timestamp 1676037725
transform 1 0 26956 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_295
timestamp 1676037725
transform 1 0 28244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_302
timestamp 1676037725
transform 1 0 28888 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_319
timestamp 1676037725
transform 1 0 30452 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_334
timestamp 1676037725
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_341
timestamp 1676037725
transform 1 0 32476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_348
timestamp 1676037725
transform 1 0 33120 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1676037725
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_371
timestamp 1676037725
transform 1 0 35236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_378
timestamp 1676037725
transform 1 0 35880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_384
timestamp 1676037725
transform 1 0 36432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_390
timestamp 1676037725
transform 1 0 36984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_396
timestamp 1676037725
transform 1 0 37536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_402
timestamp 1676037725
transform 1 0 38088 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_406
timestamp 1676037725
transform 1 0 38456 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_410
timestamp 1676037725
transform 1 0 38824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1676037725
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_426
timestamp 1676037725
transform 1 0 40296 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_444
timestamp 1676037725
transform 1 0 41952 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_456
timestamp 1676037725
transform 1 0 43056 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_133
timestamp 1676037725
transform 1 0 13340 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_194
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1676037725
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_215
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_233
timestamp 1676037725
transform 1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_247
timestamp 1676037725
transform 1 0 23828 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1676037725
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_292
timestamp 1676037725
transform 1 0 27968 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_316
timestamp 1676037725
transform 1 0 30176 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_324
timestamp 1676037725
transform 1 0 30912 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1676037725
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_344
timestamp 1676037725
transform 1 0 32752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_352
timestamp 1676037725
transform 1 0 33488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_366
timestamp 1676037725
transform 1 0 34776 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_372
timestamp 1676037725
transform 1 0 35328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_382
timestamp 1676037725
transform 1 0 36248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1676037725
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_399
timestamp 1676037725
transform 1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_415
timestamp 1676037725
transform 1 0 39284 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_421
timestamp 1676037725
transform 1 0 39836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_429
timestamp 1676037725
transform 1 0 40572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_437
timestamp 1676037725
transform 1 0 41308 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1676037725
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_456
timestamp 1676037725
transform 1 0 43056 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_159
timestamp 1676037725
transform 1 0 15732 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_171
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1676037725
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_207
timestamp 1676037725
transform 1 0 20148 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_217
timestamp 1676037725
transform 1 0 21068 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_226
timestamp 1676037725
transform 1 0 21896 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_235
timestamp 1676037725
transform 1 0 22724 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_262
timestamp 1676037725
transform 1 0 25208 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1676037725
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_287
timestamp 1676037725
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_300
timestamp 1676037725
transform 1 0 28704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1676037725
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_314
timestamp 1676037725
transform 1 0 29992 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1676037725
transform 1 0 31372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_335
timestamp 1676037725
transform 1 0 31924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_343
timestamp 1676037725
transform 1 0 32660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_349
timestamp 1676037725
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1676037725
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_372
timestamp 1676037725
transform 1 0 35328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_378
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_390
timestamp 1676037725
transform 1 0 36984 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_399
timestamp 1676037725
transform 1 0 37812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_405
timestamp 1676037725
transform 1 0 38364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_417
timestamp 1676037725
transform 1 0 39468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_431
timestamp 1676037725
transform 1 0 40756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_435
timestamp 1676037725
transform 1 0 41124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_455
timestamp 1676037725
transform 1 0 42964 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_461
timestamp 1676037725
transform 1 0 43516 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_145
timestamp 1676037725
transform 1 0 14444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1676037725
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_195
timestamp 1676037725
transform 1 0 19044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_211
timestamp 1676037725
transform 1 0 20516 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1676037725
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1676037725
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_236
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_239
timestamp 1676037725
transform 1 0 23092 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_248
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1676037725
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1676037725
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_290
timestamp 1676037725
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_298
timestamp 1676037725
transform 1 0 28520 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_304
timestamp 1676037725
transform 1 0 29072 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_313
timestamp 1676037725
transform 1 0 29900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_320
timestamp 1676037725
transform 1 0 30544 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_328
timestamp 1676037725
transform 1 0 31280 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1676037725
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_342
timestamp 1676037725
transform 1 0 32568 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_351
timestamp 1676037725
transform 1 0 33396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_355
timestamp 1676037725
transform 1 0 33764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_374
timestamp 1676037725
transform 1 0 35512 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1676037725
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1676037725
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_412
timestamp 1676037725
transform 1 0 39008 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_424
timestamp 1676037725
transform 1 0 40112 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_432
timestamp 1676037725
transform 1 0 40848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1676037725
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_457
timestamp 1676037725
transform 1 0 43148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_162
timestamp 1676037725
transform 1 0 16008 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_174
timestamp 1676037725
transform 1 0 17112 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1676037725
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_205
timestamp 1676037725
transform 1 0 19964 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1676037725
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_219
timestamp 1676037725
transform 1 0 21252 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_237
timestamp 1676037725
transform 1 0 22908 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1676037725
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_261
timestamp 1676037725
transform 1 0 25116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_268
timestamp 1676037725
transform 1 0 25760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_272
timestamp 1676037725
transform 1 0 26128 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_279
timestamp 1676037725
transform 1 0 26772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_291
timestamp 1676037725
transform 1 0 27876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_297
timestamp 1676037725
transform 1 0 28428 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1676037725
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_315
timestamp 1676037725
transform 1 0 30084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1676037725
transform 1 0 31648 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_343
timestamp 1676037725
transform 1 0 32660 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_349
timestamp 1676037725
transform 1 0 33212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_355
timestamp 1676037725
transform 1 0 33764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1676037725
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_371
timestamp 1676037725
transform 1 0 35236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_378
timestamp 1676037725
transform 1 0 35880 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_382
timestamp 1676037725
transform 1 0 36248 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_387
timestamp 1676037725
transform 1 0 36708 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_395
timestamp 1676037725
transform 1 0 37444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_409
timestamp 1676037725
transform 1 0 38732 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1676037725
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_429
timestamp 1676037725
transform 1 0 40572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_441
timestamp 1676037725
transform 1 0 41676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_451
timestamp 1676037725
transform 1 0 42596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_460
timestamp 1676037725
transform 1 0 43424 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_132
timestamp 1676037725
transform 1 0 13248 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_144
timestamp 1676037725
transform 1 0 14352 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_148
timestamp 1676037725
transform 1 0 14720 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_156
timestamp 1676037725
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_173
timestamp 1676037725
transform 1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_191
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_203
timestamp 1676037725
transform 1 0 19780 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_216
timestamp 1676037725
transform 1 0 20976 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1676037725
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_232
timestamp 1676037725
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_238
timestamp 1676037725
transform 1 0 23000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1676037725
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_267
timestamp 1676037725
transform 1 0 25668 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_292
timestamp 1676037725
transform 1 0 27968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_303
timestamp 1676037725
transform 1 0 28980 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_310
timestamp 1676037725
transform 1 0 29624 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_316
timestamp 1676037725
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_323
timestamp 1676037725
transform 1 0 30820 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1676037725
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_347
timestamp 1676037725
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1676037725
transform 1 0 33580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_366
timestamp 1676037725
transform 1 0 34776 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_379
timestamp 1676037725
transform 1 0 35972 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_397
timestamp 1676037725
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_406
timestamp 1676037725
transform 1 0 38456 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_415
timestamp 1676037725
transform 1 0 39284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_421
timestamp 1676037725
transform 1 0 39836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_425
timestamp 1676037725
transform 1 0 40204 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_440
timestamp 1676037725
transform 1 0 41584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1676037725
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_453
timestamp 1676037725
transform 1 0 42780 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_460
timestamp 1676037725
transform 1 0 43424 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1676037725
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_172
timestamp 1676037725
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_183
timestamp 1676037725
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1676037725
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_204
timestamp 1676037725
transform 1 0 19872 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_216
timestamp 1676037725
transform 1 0 20976 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_224
timestamp 1676037725
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_229
timestamp 1676037725
transform 1 0 22172 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1676037725
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_244
timestamp 1676037725
transform 1 0 23552 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_261
timestamp 1676037725
transform 1 0 25116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_267
timestamp 1676037725
transform 1 0 25668 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_292
timestamp 1676037725
transform 1 0 27968 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1676037725
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_324
timestamp 1676037725
transform 1 0 30912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_348
timestamp 1676037725
transform 1 0 33120 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1676037725
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_373
timestamp 1676037725
transform 1 0 35420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_383
timestamp 1676037725
transform 1 0 36340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_393
timestamp 1676037725
transform 1 0 37260 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_407
timestamp 1676037725
transform 1 0 38548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1676037725
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_430
timestamp 1676037725
transform 1 0 40664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_446
timestamp 1676037725
transform 1 0 42136 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_461
timestamp 1676037725
transform 1 0 43516 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_131
timestamp 1676037725
transform 1 0 13156 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_140
timestamp 1676037725
transform 1 0 13984 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_148
timestamp 1676037725
transform 1 0 14720 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1676037725
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_157
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1676037725
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_175
timestamp 1676037725
transform 1 0 17204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 1676037725
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_195
timestamp 1676037725
transform 1 0 19044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_215
timestamp 1676037725
transform 1 0 20884 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_231
timestamp 1676037725
transform 1 0 22356 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_235
timestamp 1676037725
transform 1 0 22724 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_256
timestamp 1676037725
transform 1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_267
timestamp 1676037725
transform 1 0 25668 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1676037725
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_299
timestamp 1676037725
transform 1 0 28612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_310
timestamp 1676037725
transform 1 0 29624 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_319
timestamp 1676037725
transform 1 0 30452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_328
timestamp 1676037725
transform 1 0 31280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_344
timestamp 1676037725
transform 1 0 32752 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_354
timestamp 1676037725
transform 1 0 33672 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_358
timestamp 1676037725
transform 1 0 34040 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_367
timestamp 1676037725
transform 1 0 34868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_377
timestamp 1676037725
transform 1 0 35788 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1676037725
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_401
timestamp 1676037725
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_407
timestamp 1676037725
transform 1 0 38548 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_411
timestamp 1676037725
transform 1 0 38916 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_420
timestamp 1676037725
transform 1 0 39744 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_426
timestamp 1676037725
transform 1 0 40296 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_430
timestamp 1676037725
transform 1 0 40664 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_443
timestamp 1676037725
transform 1 0 41860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_456
timestamp 1676037725
transform 1 0 43056 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_113
timestamp 1676037725
transform 1 0 11500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_131
timestamp 1676037725
transform 1 0 13156 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_146
timestamp 1676037725
transform 1 0 14536 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_154
timestamp 1676037725
transform 1 0 15272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1676037725
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_171
timestamp 1676037725
transform 1 0 16836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_178
timestamp 1676037725
transform 1 0 17480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1676037725
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_190
timestamp 1676037725
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_201
timestamp 1676037725
transform 1 0 19596 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_210
timestamp 1676037725
transform 1 0 20424 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_222
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1676037725
transform 1 0 25208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_268
timestamp 1676037725
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_288
timestamp 1676037725
transform 1 0 27600 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_294
timestamp 1676037725
transform 1 0 28152 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_300
timestamp 1676037725
transform 1 0 28704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1676037725
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_327
timestamp 1676037725
transform 1 0 31188 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_337
timestamp 1676037725
transform 1 0 32108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_346
timestamp 1676037725
transform 1 0 32936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_353
timestamp 1676037725
transform 1 0 33580 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1676037725
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_371
timestamp 1676037725
transform 1 0 35236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_379
timestamp 1676037725
transform 1 0 35972 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_386
timestamp 1676037725
transform 1 0 36616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_397
timestamp 1676037725
transform 1 0 37628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_404
timestamp 1676037725
transform 1 0 38272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_408
timestamp 1676037725
transform 1 0 38640 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1676037725
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_430
timestamp 1676037725
transform 1 0 40664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_434
timestamp 1676037725
transform 1 0 41032 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_441
timestamp 1676037725
transform 1 0 41676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_450
timestamp 1676037725
transform 1 0 42504 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_459
timestamp 1676037725
transform 1 0 43332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_122
timestamp 1676037725
transform 1 0 12328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_132
timestamp 1676037725
transform 1 0 13248 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_157
timestamp 1676037725
transform 1 0 15548 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1676037725
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_191
timestamp 1676037725
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1676037725
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_211
timestamp 1676037725
transform 1 0 20516 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1676037725
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_239
timestamp 1676037725
transform 1 0 23092 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1676037725
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_271
timestamp 1676037725
transform 1 0 26036 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1676037725
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_291
timestamp 1676037725
transform 1 0 27876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_302
timestamp 1676037725
transform 1 0 28888 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_308
timestamp 1676037725
transform 1 0 29440 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_312
timestamp 1676037725
transform 1 0 29808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_318
timestamp 1676037725
transform 1 0 30360 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_324
timestamp 1676037725
transform 1 0 30912 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1676037725
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1676037725
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_346
timestamp 1676037725
transform 1 0 32936 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_354
timestamp 1676037725
transform 1 0 33672 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_364
timestamp 1676037725
transform 1 0 34592 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_372
timestamp 1676037725
transform 1 0 35328 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_378
timestamp 1676037725
transform 1 0 35880 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_386
timestamp 1676037725
transform 1 0 36616 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1676037725
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_403
timestamp 1676037725
transform 1 0 38180 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_416
timestamp 1676037725
transform 1 0 39376 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_423
timestamp 1676037725
transform 1 0 40020 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_436
timestamp 1676037725
transform 1 0 41216 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1676037725
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_457
timestamp 1676037725
transform 1 0 43148 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_145
timestamp 1676037725
transform 1 0 14444 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_173
timestamp 1676037725
transform 1 0 17020 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_178
timestamp 1676037725
transform 1 0 17480 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_186
timestamp 1676037725
transform 1 0 18216 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_206
timestamp 1676037725
transform 1 0 20056 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_212
timestamp 1676037725
transform 1 0 20608 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1676037725
transform 1 0 20884 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_222
timestamp 1676037725
transform 1 0 21528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_232
timestamp 1676037725
transform 1 0 22448 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_241
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1676037725
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_273
timestamp 1676037725
transform 1 0 26220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_279
timestamp 1676037725
transform 1 0 26772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_300
timestamp 1676037725
transform 1 0 28704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1676037725
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_317
timestamp 1676037725
transform 1 0 30268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_323
timestamp 1676037725
transform 1 0 30820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_331
timestamp 1676037725
transform 1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_337
timestamp 1676037725
transform 1 0 32108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_349
timestamp 1676037725
transform 1 0 33212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1676037725
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_376
timestamp 1676037725
transform 1 0 35696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_385
timestamp 1676037725
transform 1 0 36524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_397
timestamp 1676037725
transform 1 0 37628 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_406
timestamp 1676037725
transform 1 0 38456 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_414
timestamp 1676037725
transform 1 0 39192 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 1676037725
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_426
timestamp 1676037725
transform 1 0 40296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_439
timestamp 1676037725
transform 1 0 41492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_446
timestamp 1676037725
transform 1 0 42136 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_460
timestamp 1676037725
transform 1 0 43424 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_117
timestamp 1676037725
transform 1 0 11868 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_122
timestamp 1676037725
transform 1 0 12328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_135
timestamp 1676037725
transform 1 0 13524 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_144
timestamp 1676037725
transform 1 0 14352 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_150
timestamp 1676037725
transform 1 0 14904 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1676037725
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_176
timestamp 1676037725
transform 1 0 17296 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_192
timestamp 1676037725
transform 1 0 18768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_198
timestamp 1676037725
transform 1 0 19320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_214
timestamp 1676037725
transform 1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1676037725
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_244
timestamp 1676037725
transform 1 0 23552 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_257
timestamp 1676037725
transform 1 0 24748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_263
timestamp 1676037725
transform 1 0 25300 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1676037725
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_306
timestamp 1676037725
transform 1 0 29256 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_312
timestamp 1676037725
transform 1 0 29808 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_320
timestamp 1676037725
transform 1 0 30544 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_328
timestamp 1676037725
transform 1 0 31280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1676037725
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_346
timestamp 1676037725
transform 1 0 32936 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_352
timestamp 1676037725
transform 1 0 33488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1676037725
transform 1 0 34408 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_371
timestamp 1676037725
transform 1 0 35236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_382
timestamp 1676037725
transform 1 0 36248 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1676037725
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_401
timestamp 1676037725
transform 1 0 37996 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_410
timestamp 1676037725
transform 1 0 38824 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_430
timestamp 1676037725
transform 1 0 40664 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_438
timestamp 1676037725
transform 1 0 41400 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_446
timestamp 1676037725
transform 1 0 42136 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_457
timestamp 1676037725
transform 1 0 43148 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_126
timestamp 1676037725
transform 1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1676037725
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1676037725
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_150
timestamp 1676037725
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_156
timestamp 1676037725
transform 1 0 15456 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_169
timestamp 1676037725
transform 1 0 16652 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_175
timestamp 1676037725
transform 1 0 17204 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_188
timestamp 1676037725
transform 1 0 18400 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1676037725
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_215
timestamp 1676037725
transform 1 0 20884 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_223
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_230
timestamp 1676037725
transform 1 0 22264 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1676037725
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_263
timestamp 1676037725
transform 1 0 25300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp 1676037725
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_285
timestamp 1676037725
transform 1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_291
timestamp 1676037725
transform 1 0 27876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_299
timestamp 1676037725
transform 1 0 28612 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_313
timestamp 1676037725
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_318
timestamp 1676037725
transform 1 0 30360 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_324
timestamp 1676037725
transform 1 0 30912 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_329
timestamp 1676037725
transform 1 0 31372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_340
timestamp 1676037725
transform 1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_348
timestamp 1676037725
transform 1 0 33120 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_354
timestamp 1676037725
transform 1 0 33672 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1676037725
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_372
timestamp 1676037725
transform 1 0 35328 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_386
timestamp 1676037725
transform 1 0 36616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_392
timestamp 1676037725
transform 1 0 37168 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_396
timestamp 1676037725
transform 1 0 37536 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_405
timestamp 1676037725
transform 1 0 38364 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1676037725
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_431
timestamp 1676037725
transform 1 0 40756 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_437
timestamp 1676037725
transform 1 0 41308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_458
timestamp 1676037725
transform 1 0 43240 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_133
timestamp 1676037725
transform 1 0 13340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_143
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_153
timestamp 1676037725
transform 1 0 15180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_177
timestamp 1676037725
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_185
timestamp 1676037725
transform 1 0 18124 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_199
timestamp 1676037725
transform 1 0 19412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_215
timestamp 1676037725
transform 1 0 20884 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1676037725
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_242
timestamp 1676037725
transform 1 0 23368 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1676037725
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_285
timestamp 1676037725
transform 1 0 27324 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_297
timestamp 1676037725
transform 1 0 28428 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_301
timestamp 1676037725
transform 1 0 28796 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_310
timestamp 1676037725
transform 1 0 29624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_327
timestamp 1676037725
transform 1 0 31188 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1676037725
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_347
timestamp 1676037725
transform 1 0 33028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_351
timestamp 1676037725
transform 1 0 33396 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_356
timestamp 1676037725
transform 1 0 33856 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_362
timestamp 1676037725
transform 1 0 34408 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_366
timestamp 1676037725
transform 1 0 34776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_383
timestamp 1676037725
transform 1 0 36340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1676037725
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1676037725
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_420
timestamp 1676037725
transform 1 0 39744 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_434
timestamp 1676037725
transform 1 0 41032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_454
timestamp 1676037725
transform 1 0 42872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_460
timestamp 1676037725
transform 1 0 43424 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_126
timestamp 1676037725
transform 1 0 12696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_134
timestamp 1676037725
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_149
timestamp 1676037725
transform 1 0 14812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_162
timestamp 1676037725
transform 1 0 16008 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_171
timestamp 1676037725
transform 1 0 16836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 1676037725
transform 1 0 17940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_187
timestamp 1676037725
transform 1 0 18308 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1676037725
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_203
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_213
timestamp 1676037725
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_226
timestamp 1676037725
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_237
timestamp 1676037725
transform 1 0 22908 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1676037725
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_257
timestamp 1676037725
transform 1 0 24748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1676037725
transform 1 0 26036 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_275
timestamp 1676037725
transform 1 0 26404 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_283
timestamp 1676037725
transform 1 0 27140 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_292
timestamp 1676037725
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_296
timestamp 1676037725
transform 1 0 28336 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1676037725
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_315
timestamp 1676037725
transform 1 0 30084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_323
timestamp 1676037725
transform 1 0 30820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_329
timestamp 1676037725
transform 1 0 31372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_340
timestamp 1676037725
transform 1 0 32384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_348
timestamp 1676037725
transform 1 0 33120 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_354
timestamp 1676037725
transform 1 0 33672 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1676037725
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_371
timestamp 1676037725
transform 1 0 35236 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_381
timestamp 1676037725
transform 1 0 36156 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_390
timestamp 1676037725
transform 1 0 36984 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_399
timestamp 1676037725
transform 1 0 37812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_405
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1676037725
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_426
timestamp 1676037725
transform 1 0 40296 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_460
timestamp 1676037725
transform 1 0 43424 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_119
timestamp 1676037725
transform 1 0 12052 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_122
timestamp 1676037725
transform 1 0 12328 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_132
timestamp 1676037725
transform 1 0 13248 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_142
timestamp 1676037725
transform 1 0 14168 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_150
timestamp 1676037725
transform 1 0 14904 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1676037725
transform 1 0 15180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1676037725
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1676037725
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_178
timestamp 1676037725
transform 1 0 17480 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_185
timestamp 1676037725
transform 1 0 18124 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_202
timestamp 1676037725
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_213
timestamp 1676037725
transform 1 0 20700 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1676037725
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_229
timestamp 1676037725
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_234
timestamp 1676037725
transform 1 0 22632 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_248
timestamp 1676037725
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_255
timestamp 1676037725
transform 1 0 24564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_266
timestamp 1676037725
transform 1 0 25576 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_272
timestamp 1676037725
transform 1 0 26128 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1676037725
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_285
timestamp 1676037725
transform 1 0 27324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_289
timestamp 1676037725
transform 1 0 27692 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_298
timestamp 1676037725
transform 1 0 28520 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_304
timestamp 1676037725
transform 1 0 29072 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_316
timestamp 1676037725
transform 1 0 30176 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_322
timestamp 1676037725
transform 1 0 30728 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_327
timestamp 1676037725
transform 1 0 31188 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_345
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_364
timestamp 1676037725
transform 1 0 34592 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_381
timestamp 1676037725
transform 1 0 36156 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1676037725
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_404
timestamp 1676037725
transform 1 0 38272 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_412
timestamp 1676037725
transform 1 0 39008 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_418
timestamp 1676037725
transform 1 0 39560 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_424
timestamp 1676037725
transform 1 0 40112 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_435
timestamp 1676037725
transform 1 0 41124 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_446
timestamp 1676037725
transform 1 0 42136 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_454
timestamp 1676037725
transform 1 0 42872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_460
timestamp 1676037725
transform 1 0 43424 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_127
timestamp 1676037725
transform 1 0 12788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_149
timestamp 1676037725
transform 1 0 14812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_156
timestamp 1676037725
transform 1 0 15456 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_173
timestamp 1676037725
transform 1 0 17020 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_188
timestamp 1676037725
transform 1 0 18400 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_203
timestamp 1676037725
transform 1 0 19780 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_206
timestamp 1676037725
transform 1 0 20056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_216
timestamp 1676037725
transform 1 0 20976 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_222
timestamp 1676037725
transform 1 0 21528 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_230
timestamp 1676037725
transform 1 0 22264 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_238
timestamp 1676037725
transform 1 0 23000 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1676037725
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1676037725
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_273
timestamp 1676037725
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_283
timestamp 1676037725
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1676037725
transform 1 0 28244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_299
timestamp 1676037725
transform 1 0 28612 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1676037725
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_314
timestamp 1676037725
transform 1 0 29992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_320
timestamp 1676037725
transform 1 0 30544 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_328
timestamp 1676037725
transform 1 0 31280 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_337
timestamp 1676037725
transform 1 0 32108 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_353
timestamp 1676037725
transform 1 0 33580 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1676037725
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_369
timestamp 1676037725
transform 1 0 35052 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_381
timestamp 1676037725
transform 1 0 36156 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_396
timestamp 1676037725
transform 1 0 37536 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_407
timestamp 1676037725
transform 1 0 38548 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_417
timestamp 1676037725
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_439
timestamp 1676037725
transform 1 0 41492 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_459
timestamp 1676037725
transform 1 0 43332 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_133
timestamp 1676037725
transform 1 0 13340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_141
timestamp 1676037725
transform 1 0 14076 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_151
timestamp 1676037725
transform 1 0 14996 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_159
timestamp 1676037725
transform 1 0 15732 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_178
timestamp 1676037725
transform 1 0 17480 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_201
timestamp 1676037725
transform 1 0 19596 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1676037725
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_235
timestamp 1676037725
transform 1 0 22724 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_252
timestamp 1676037725
transform 1 0 24288 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1676037725
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1676037725
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_308
timestamp 1676037725
transform 1 0 29440 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1676037725
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_324
timestamp 1676037725
transform 1 0 30912 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_328
timestamp 1676037725
transform 1 0 31280 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1676037725
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_350
timestamp 1676037725
transform 1 0 33304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_365
timestamp 1676037725
transform 1 0 34684 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_380
timestamp 1676037725
transform 1 0 36064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1676037725
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_402
timestamp 1676037725
transform 1 0 38088 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_422
timestamp 1676037725
transform 1 0 39928 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_428
timestamp 1676037725
transform 1 0 40480 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_434
timestamp 1676037725
transform 1 0 41032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_440
timestamp 1676037725
transform 1 0 41584 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1676037725
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_454
timestamp 1676037725
transform 1 0 42872 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_460
timestamp 1676037725
transform 1 0 43424 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_148
timestamp 1676037725
transform 1 0 14720 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_157
timestamp 1676037725
transform 1 0 15548 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_172
timestamp 1676037725
transform 1 0 16928 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_178
timestamp 1676037725
transform 1 0 17480 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_188
timestamp 1676037725
transform 1 0 18400 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_203
timestamp 1676037725
transform 1 0 19780 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_222
timestamp 1676037725
transform 1 0 21528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_234
timestamp 1676037725
transform 1 0 22632 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1676037725
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_269
timestamp 1676037725
transform 1 0 25852 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_275
timestamp 1676037725
transform 1 0 26404 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_284
timestamp 1676037725
transform 1 0 27232 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_292
timestamp 1676037725
transform 1 0 27968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1676037725
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_328
timestamp 1676037725
transform 1 0 31280 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_336
timestamp 1676037725
transform 1 0 32016 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_344
timestamp 1676037725
transform 1 0 32752 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1676037725
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_384
timestamp 1676037725
transform 1 0 36432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_390
timestamp 1676037725
transform 1 0 36984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_399
timestamp 1676037725
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_406
timestamp 1676037725
transform 1 0 38456 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_412
timestamp 1676037725
transform 1 0 39008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_418
timestamp 1676037725
transform 1 0 39560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_427
timestamp 1676037725
transform 1 0 40388 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_435
timestamp 1676037725
transform 1 0 41124 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_455
timestamp 1676037725
transform 1 0 42964 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_461
timestamp 1676037725
transform 1 0 43516 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1676037725
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_147
timestamp 1676037725
transform 1 0 14628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_154
timestamp 1676037725
transform 1 0 15272 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_160
timestamp 1676037725
transform 1 0 15824 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1676037725
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_177
timestamp 1676037725
transform 1 0 17388 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_184
timestamp 1676037725
transform 1 0 18032 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_207
timestamp 1676037725
transform 1 0 20148 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_213
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_216
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_244
timestamp 1676037725
transform 1 0 23552 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_256
timestamp 1676037725
transform 1 0 24656 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_272
timestamp 1676037725
transform 1 0 26128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_291
timestamp 1676037725
transform 1 0 27876 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_297
timestamp 1676037725
transform 1 0 28428 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_306
timestamp 1676037725
transform 1 0 29256 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_318
timestamp 1676037725
transform 1 0 30360 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_324
timestamp 1676037725
transform 1 0 30912 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1676037725
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_348
timestamp 1676037725
transform 1 0 33120 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_356
timestamp 1676037725
transform 1 0 33856 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_363
timestamp 1676037725
transform 1 0 34500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_382
timestamp 1676037725
transform 1 0 36248 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1676037725
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1676037725
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_409
timestamp 1676037725
transform 1 0 38732 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_415
timestamp 1676037725
transform 1 0 39284 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_424
timestamp 1676037725
transform 1 0 40112 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_436
timestamp 1676037725
transform 1 0 41216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_445
timestamp 1676037725
transform 1 0 42044 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_454
timestamp 1676037725
transform 1 0 42872 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_460
timestamp 1676037725
transform 1 0 43424 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1676037725
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_102
timestamp 1676037725
transform 1 0 10488 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_114
timestamp 1676037725
transform 1 0 11592 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_126
timestamp 1676037725
transform 1 0 12696 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_160
timestamp 1676037725
transform 1 0 15824 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_183
timestamp 1676037725
transform 1 0 17940 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_191
timestamp 1676037725
transform 1 0 18676 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_208
timestamp 1676037725
transform 1 0 20240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_212
timestamp 1676037725
transform 1 0 20608 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1676037725
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_239
timestamp 1676037725
transform 1 0 23092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_267
timestamp 1676037725
transform 1 0 25668 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_278
timestamp 1676037725
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_299
timestamp 1676037725
transform 1 0 28612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1676037725
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_323
timestamp 1676037725
transform 1 0 30820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_334
timestamp 1676037725
transform 1 0 31832 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_346
timestamp 1676037725
transform 1 0 32936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_371
timestamp 1676037725
transform 1 0 35236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_379
timestamp 1676037725
transform 1 0 35972 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1676037725
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_407
timestamp 1676037725
transform 1 0 38548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1676037725
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_431
timestamp 1676037725
transform 1 0 40756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_440
timestamp 1676037725
transform 1 0 41584 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_460
timestamp 1676037725
transform 1 0 43424 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_142
timestamp 1676037725
transform 1 0 14168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_148
timestamp 1676037725
transform 1 0 14720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_154
timestamp 1676037725
transform 1 0 15272 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_160
timestamp 1676037725
transform 1 0 15824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1676037725
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_188
timestamp 1676037725
transform 1 0 18400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_208
timestamp 1676037725
transform 1 0 20240 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_216
timestamp 1676037725
transform 1 0 20976 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_236
timestamp 1676037725
transform 1 0 22816 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_244
timestamp 1676037725
transform 1 0 23552 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1676037725
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_263
timestamp 1676037725
transform 1 0 25300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_267
timestamp 1676037725
transform 1 0 25668 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1676037725
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_290
timestamp 1676037725
transform 1 0 27784 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_294
timestamp 1676037725
transform 1 0 28152 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_309
timestamp 1676037725
transform 1 0 29532 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_320
timestamp 1676037725
transform 1 0 30544 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_326
timestamp 1676037725
transform 1 0 31096 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1676037725
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_348
timestamp 1676037725
transform 1 0 33120 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_362
timestamp 1676037725
transform 1 0 34408 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_376
timestamp 1676037725
transform 1 0 35696 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_382
timestamp 1676037725
transform 1 0 36248 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1676037725
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_397
timestamp 1676037725
transform 1 0 37628 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_420
timestamp 1676037725
transform 1 0 39744 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_432
timestamp 1676037725
transform 1 0 40848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_439
timestamp 1676037725
transform 1 0 41492 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_446
timestamp 1676037725
transform 1 0 42136 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_453
timestamp 1676037725
transform 1 0 42780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_460
timestamp 1676037725
transform 1 0 43424 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1676037725
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_152
timestamp 1676037725
transform 1 0 15088 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_158
timestamp 1676037725
transform 1 0 15640 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1676037725
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_170
timestamp 1676037725
transform 1 0 16744 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_176
timestamp 1676037725
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_182
timestamp 1676037725
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_188
timestamp 1676037725
transform 1 0 18400 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_202
timestamp 1676037725
transform 1 0 19688 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1676037725
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_234
timestamp 1676037725
transform 1 0 22632 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_269
timestamp 1676037725
transform 1 0 25852 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_284
timestamp 1676037725
transform 1 0 27232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_302
timestamp 1676037725
transform 1 0 28888 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_329
timestamp 1676037725
transform 1 0 31372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_341
timestamp 1676037725
transform 1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_347
timestamp 1676037725
transform 1 0 33028 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1676037725
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_375
timestamp 1676037725
transform 1 0 35604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_390
timestamp 1676037725
transform 1 0 36984 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_411
timestamp 1676037725
transform 1 0 38916 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1676037725
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_431
timestamp 1676037725
transform 1 0 40756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_439
timestamp 1676037725
transform 1 0 41492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_459
timestamp 1676037725
transform 1 0 43332 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_154
timestamp 1676037725
transform 1 0 15272 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_160
timestamp 1676037725
transform 1 0 15824 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_173
timestamp 1676037725
transform 1 0 17020 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_176
timestamp 1676037725
transform 1 0 17296 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_182
timestamp 1676037725
transform 1 0 17848 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_189
timestamp 1676037725
transform 1 0 18492 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_202
timestamp 1676037725
transform 1 0 19688 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1676037725
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_235
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1676037725
transform 1 0 23460 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_258
timestamp 1676037725
transform 1 0 24840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_270
timestamp 1676037725
transform 1 0 25944 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1676037725
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_292
timestamp 1676037725
transform 1 0 27968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_304
timestamp 1676037725
transform 1 0 29072 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_315
timestamp 1676037725
transform 1 0 30084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_323
timestamp 1676037725
transform 1 0 30820 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1676037725
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_346
timestamp 1676037725
transform 1 0 32936 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_352
timestamp 1676037725
transform 1 0 33488 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_364
timestamp 1676037725
transform 1 0 34592 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_378
timestamp 1676037725
transform 1 0 35880 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1676037725
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_397
timestamp 1676037725
transform 1 0 37628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_401
timestamp 1676037725
transform 1 0 37996 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_419
timestamp 1676037725
transform 1 0 39652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_431
timestamp 1676037725
transform 1 0 40756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_440
timestamp 1676037725
transform 1 0 41584 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_446
timestamp 1676037725
transform 1 0 42136 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_453
timestamp 1676037725
transform 1 0 42780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_459
timestamp 1676037725
transform 1 0 43332 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_168
timestamp 1676037725
transform 1 0 16560 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_174
timestamp 1676037725
transform 1 0 17112 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1676037725
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_208
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_212
timestamp 1676037725
transform 1 0 20608 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_239
timestamp 1676037725
transform 1 0 23092 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1676037725
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_263
timestamp 1676037725
transform 1 0 25300 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_269
timestamp 1676037725
transform 1 0 25852 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_281
timestamp 1676037725
transform 1 0 26956 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_287
timestamp 1676037725
transform 1 0 27508 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_291
timestamp 1676037725
transform 1 0 27876 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_300
timestamp 1676037725
transform 1 0 28704 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1676037725
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_316
timestamp 1676037725
transform 1 0 30176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_322
timestamp 1676037725
transform 1 0 30728 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_326
timestamp 1676037725
transform 1 0 31096 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_334
timestamp 1676037725
transform 1 0 31832 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_342
timestamp 1676037725
transform 1 0 32568 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_374
timestamp 1676037725
transform 1 0 35512 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_380
timestamp 1676037725
transform 1 0 36064 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_384
timestamp 1676037725
transform 1 0 36432 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_402
timestamp 1676037725
transform 1 0 38088 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_408
timestamp 1676037725
transform 1 0 38640 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_414
timestamp 1676037725
transform 1 0 39192 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_427
timestamp 1676037725
transform 1 0 40388 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_440
timestamp 1676037725
transform 1 0 41584 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_460
timestamp 1676037725
transform 1 0 43424 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_173
timestamp 1676037725
transform 1 0 17020 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_179
timestamp 1676037725
transform 1 0 17572 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_185
timestamp 1676037725
transform 1 0 18124 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_215
timestamp 1676037725
transform 1 0 20884 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_219
timestamp 1676037725
transform 1 0 21252 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1676037725
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_235
timestamp 1676037725
transform 1 0 22724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_241
timestamp 1676037725
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_254
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_262
timestamp 1676037725
transform 1 0 25208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_268
timestamp 1676037725
transform 1 0 25760 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1676037725
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_299
timestamp 1676037725
transform 1 0 28612 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_307
timestamp 1676037725
transform 1 0 29348 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_313
timestamp 1676037725
transform 1 0 29900 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_326
timestamp 1676037725
transform 1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1676037725
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_341
timestamp 1676037725
transform 1 0 32476 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_362
timestamp 1676037725
transform 1 0 34408 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_383
timestamp 1676037725
transform 1 0 36340 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1676037725
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_411
timestamp 1676037725
transform 1 0 38916 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_428
timestamp 1676037725
transform 1 0 40480 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_437
timestamp 1676037725
transform 1 0 41308 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_443
timestamp 1676037725
transform 1 0 41860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_453
timestamp 1676037725
transform 1 0 42780 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_459
timestamp 1676037725
transform 1 0 43332 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_182
timestamp 1676037725
transform 1 0 17848 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_188
timestamp 1676037725
transform 1 0 18400 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_202
timestamp 1676037725
transform 1 0 19688 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_212
timestamp 1676037725
transform 1 0 20608 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_232
timestamp 1676037725
transform 1 0 22448 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_238
timestamp 1676037725
transform 1 0 23000 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_246
timestamp 1676037725
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_257
timestamp 1676037725
transform 1 0 24748 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_263
timestamp 1676037725
transform 1 0 25300 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_269
timestamp 1676037725
transform 1 0 25852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_280
timestamp 1676037725
transform 1 0 26864 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_300
timestamp 1676037725
transform 1 0 28704 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1676037725
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_313
timestamp 1676037725
transform 1 0 29900 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_339
timestamp 1676037725
transform 1 0 32292 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_352
timestamp 1676037725
transform 1 0 33488 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_358
timestamp 1676037725
transform 1 0 34040 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_374
timestamp 1676037725
transform 1 0 35512 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_383
timestamp 1676037725
transform 1 0 36340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_391
timestamp 1676037725
transform 1 0 37076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_397
timestamp 1676037725
transform 1 0 37628 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_403
timestamp 1676037725
transform 1 0 38180 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1676037725
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_439
timestamp 1676037725
transform 1 0 41492 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_459
timestamp 1676037725
transform 1 0 43332 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_195
timestamp 1676037725
transform 1 0 19044 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_202
timestamp 1676037725
transform 1 0 19688 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_231
timestamp 1676037725
transform 1 0 22356 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_242
timestamp 1676037725
transform 1 0 23368 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_248
timestamp 1676037725
transform 1 0 23920 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_259
timestamp 1676037725
transform 1 0 24932 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_268
timestamp 1676037725
transform 1 0 25760 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_274
timestamp 1676037725
transform 1 0 26312 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_285
timestamp 1676037725
transform 1 0 27324 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_291
timestamp 1676037725
transform 1 0 27876 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_313
timestamp 1676037725
transform 1 0 29900 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_319
timestamp 1676037725
transform 1 0 30452 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_327
timestamp 1676037725
transform 1 0 31188 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1676037725
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_341
timestamp 1676037725
transform 1 0 32476 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_354
timestamp 1676037725
transform 1 0 33672 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_367
timestamp 1676037725
transform 1 0 34868 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_371
timestamp 1676037725
transform 1 0 35236 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_388
timestamp 1676037725
transform 1 0 36800 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_397
timestamp 1676037725
transform 1 0 37628 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_403
timestamp 1676037725
transform 1 0 38180 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_409
timestamp 1676037725
transform 1 0 38732 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_415
timestamp 1676037725
transform 1 0 39284 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_421
timestamp 1676037725
transform 1 0 39836 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_427
timestamp 1676037725
transform 1 0 40388 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_433
timestamp 1676037725
transform 1 0 40940 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_439
timestamp 1676037725
transform 1 0 41492 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_445
timestamp 1676037725
transform 1 0 42044 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_453
timestamp 1676037725
transform 1 0 42780 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_457
timestamp 1676037725
transform 1 0 43148 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_460
timestamp 1676037725
transform 1 0 43424 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1676037725
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_203
timestamp 1676037725
transform 1 0 19780 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_206
timestamp 1676037725
transform 1 0 20056 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_217
timestamp 1676037725
transform 1 0 21068 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_223
timestamp 1676037725
transform 1 0 21620 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_227
timestamp 1676037725
transform 1 0 21988 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_230
timestamp 1676037725
transform 1 0 22264 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_259
timestamp 1676037725
transform 1 0 24932 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_276
timestamp 1676037725
transform 1 0 26496 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_282
timestamp 1676037725
transform 1 0 27048 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_288
timestamp 1676037725
transform 1 0 27600 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_291
timestamp 1676037725
transform 1 0 27876 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_299
timestamp 1676037725
transform 1 0 28612 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_305
timestamp 1676037725
transform 1 0 29164 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_313
timestamp 1676037725
transform 1 0 29900 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_319
timestamp 1676037725
transform 1 0 30452 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_325
timestamp 1676037725
transform 1 0 31004 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_329
timestamp 1676037725
transform 1 0 31372 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_339
timestamp 1676037725
transform 1 0 32292 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_359
timestamp 1676037725
transform 1 0 34132 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_369
timestamp 1676037725
transform 1 0 35052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_390
timestamp 1676037725
transform 1 0 36984 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_403
timestamp 1676037725
transform 1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1676037725
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_439
timestamp 1676037725
transform 1 0 41492 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_451
timestamp 1676037725
transform 1 0 42596 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_461
timestamp 1676037725
transform 1 0 43516 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_203
timestamp 1676037725
transform 1 0 19780 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_209
timestamp 1676037725
transform 1 0 20332 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1676037725
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_229
timestamp 1676037725
transform 1 0 22172 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_232
timestamp 1676037725
transform 1 0 22448 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_245
timestamp 1676037725
transform 1 0 23644 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_251
timestamp 1676037725
transform 1 0 24196 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_259
timestamp 1676037725
transform 1 0 24932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_272
timestamp 1676037725
transform 1 0 26128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1676037725
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_292
timestamp 1676037725
transform 1 0 27968 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_311
timestamp 1676037725
transform 1 0 29716 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_330
timestamp 1676037725
transform 1 0 31464 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_355
timestamp 1676037725
transform 1 0 33764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_370
timestamp 1676037725
transform 1 0 35144 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 1676037725
transform 1 0 36984 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_411
timestamp 1676037725
transform 1 0 38916 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_431
timestamp 1676037725
transform 1 0 40756 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_438
timestamp 1676037725
transform 1 0 41400 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1676037725
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_453
timestamp 1676037725
transform 1 0 42780 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_459
timestamp 1676037725
transform 1 0 43332 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_229
timestamp 1676037725
transform 1 0 22172 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_246
timestamp 1676037725
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_276
timestamp 1676037725
transform 1 0 26496 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_296
timestamp 1676037725
transform 1 0 28336 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1676037725
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_327
timestamp 1676037725
transform 1 0 31188 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_347
timestamp 1676037725
transform 1 0 33028 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_383
timestamp 1676037725
transform 1 0 36340 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_390
timestamp 1676037725
transform 1 0 36984 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_394
timestamp 1676037725
transform 1 0 37352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_398
timestamp 1676037725
transform 1 0 37720 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_404
timestamp 1676037725
transform 1 0 38272 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_411
timestamp 1676037725
transform 1 0 38916 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_417
timestamp 1676037725
transform 1 0 39468 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_432
timestamp 1676037725
transform 1 0 40848 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_438
timestamp 1676037725
transform 1 0 41400 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_447
timestamp 1676037725
transform 1 0 42228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_453
timestamp 1676037725
transform 1 0 42780 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_459
timestamp 1676037725
transform 1 0 43332 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_29
timestamp 1676037725
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_41
timestamp 1676037725
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1676037725
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_85
timestamp 1676037725
transform 1 0 8924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_97
timestamp 1676037725
transform 1 0 10028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_109
timestamp 1676037725
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_141
timestamp 1676037725
transform 1 0 14076 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_146
timestamp 1676037725
transform 1 0 14536 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_154
timestamp 1676037725
transform 1 0 15272 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_159
timestamp 1676037725
transform 1 0 15732 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_197
timestamp 1676037725
transform 1 0 19228 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_203
timestamp 1676037725
transform 1 0 19780 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_206
timestamp 1676037725
transform 1 0 20056 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_213
timestamp 1676037725
transform 1 0 20700 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_219
timestamp 1676037725
transform 1 0 21252 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_229
timestamp 1676037725
transform 1 0 22172 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_236
timestamp 1676037725
transform 1 0 22816 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_244
timestamp 1676037725
transform 1 0 23552 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_250
timestamp 1676037725
transform 1 0 24104 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_253
timestamp 1676037725
transform 1 0 24380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_258
timestamp 1676037725
transform 1 0 24840 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_265
timestamp 1676037725
transform 1 0 25484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_269
timestamp 1676037725
transform 1 0 25852 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_272
timestamp 1676037725
transform 1 0 26128 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1676037725
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_286
timestamp 1676037725
transform 1 0 27416 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_292
timestamp 1676037725
transform 1 0 27968 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_298
timestamp 1676037725
transform 1 0 28520 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_306
timestamp 1676037725
transform 1 0 29256 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_309
timestamp 1676037725
transform 1 0 29532 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_313
timestamp 1676037725
transform 1 0 29900 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_324
timestamp 1676037725
transform 1 0 30912 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_328
timestamp 1676037725
transform 1 0 31280 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_331
timestamp 1676037725
transform 1 0 31556 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_342
timestamp 1676037725
transform 1 0 32568 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_350
timestamp 1676037725
transform 1 0 33304 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_356
timestamp 1676037725
transform 1 0 33856 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_362
timestamp 1676037725
transform 1 0 34408 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_365
timestamp 1676037725
transform 1 0 34684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_370
timestamp 1676037725
transform 1 0 35144 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_376
timestamp 1676037725
transform 1 0 35696 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_382
timestamp 1676037725
transform 1 0 36248 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1676037725
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_397
timestamp 1676037725
transform 1 0 37628 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_403
timestamp 1676037725
transform 1 0 38180 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_409
timestamp 1676037725
transform 1 0 38732 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_415
timestamp 1676037725
transform 1 0 39284 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_419
timestamp 1676037725
transform 1 0 39652 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_421
timestamp 1676037725
transform 1 0 39836 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_425
timestamp 1676037725
transform 1 0 40204 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_431
timestamp 1676037725
transform 1 0 40756 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_437
timestamp 1676037725
transform 1 0 41308 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_443
timestamp 1676037725
transform 1 0 41860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_453
timestamp 1676037725
transform 1 0 42780 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_460
timestamp 1676037725
transform 1 0 43424 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 43884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 43884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 43884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 43884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 43884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 43884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 43884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 43884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 43884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 43884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 43884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 43884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 43884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 43884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 43884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 43884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 43884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 43884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 43884 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 43884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 43884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 43884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 43884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 43884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 43884 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 43884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 43884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 43884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 43884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 43884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 43884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 43884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 43884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 43884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 43884 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 43884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 43884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 43884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 43884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 43884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 43884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 43884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 43884 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 43884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 43884 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 43884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 43884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 43884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 43884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 43884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 43884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 43884 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 43884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 43884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 43884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 43884 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 43884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 43884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 43884 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 34592 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 36156 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42596 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 40848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0980_
timestamp 1676037725
transform -1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 1676037725
transform 1 0 40480 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0982_
timestamp 1676037725
transform -1 0 40388 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1676037725
transform -1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 43148 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0985_
timestamp 1676037725
transform -1 0 42136 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 41492 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 40572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1676037725
transform 1 0 40756 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0989_
timestamp 1676037725
transform 1 0 41860 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 1676037725
transform -1 0 39560 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 43332 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0993_
timestamp 1676037725
transform 1 0 34868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0994_
timestamp 1676037725
transform -1 0 43148 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0995_
timestamp 1676037725
transform -1 0 42596 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 38824 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0997_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0998_
timestamp 1676037725
transform 1 0 40940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0999_
timestamp 1676037725
transform -1 0 40572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_4  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31556 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1002_
timestamp 1676037725
transform -1 0 43148 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1003_
timestamp 1676037725
transform -1 0 42136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 42412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1676037725
transform -1 0 41676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1007_
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1676037725
transform -1 0 34408 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1676037725
transform -1 0 32752 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32384 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1012_
timestamp 1676037725
transform 1 0 33304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 42964 0 1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_1  _1014_
timestamp 1676037725
transform 1 0 33120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1015_
timestamp 1676037725
transform 1 0 33120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1676037725
transform 1 0 28428 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1017_
timestamp 1676037725
transform 1 0 28704 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1018_
timestamp 1676037725
transform 1 0 33856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1019_
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1676037725
transform -1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1676037725
transform -1 0 35880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1022_
timestamp 1676037725
transform -1 0 41676 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp 1676037725
transform -1 0 36984 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1024_
timestamp 1676037725
transform -1 0 42136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1025_
timestamp 1676037725
transform -1 0 40296 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1026_
timestamp 1676037725
transform -1 0 40020 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42964 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1028_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36616 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1029_
timestamp 1676037725
transform 1 0 36984 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1676037725
transform -1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1031_
timestamp 1676037725
transform -1 0 42504 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1033_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1034_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36708 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1676037725
transform -1 0 42228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1036_
timestamp 1676037725
transform -1 0 41216 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1037_
timestamp 1676037725
transform -1 0 32936 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _1038_
timestamp 1676037725
transform -1 0 41952 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1039_
timestamp 1676037725
transform -1 0 33948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1040_
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1041_
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1676037725
transform 1 0 30820 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1043_
timestamp 1676037725
transform 1 0 31556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_4  _1044_
timestamp 1676037725
transform -1 0 42136 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1045_
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_4  _1046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1047_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25116 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1048_
timestamp 1676037725
transform -1 0 25116 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1676037725
transform 1 0 14904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _1050_
timestamp 1676037725
transform -1 0 41860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1051_
timestamp 1676037725
transform -1 0 34592 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37996 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1053_
timestamp 1676037725
transform -1 0 36708 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42320 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 43148 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1056_
timestamp 1676037725
transform -1 0 39284 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 1676037725
transform -1 0 38456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1676037725
transform -1 0 37812 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 41584 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1061_
timestamp 1676037725
transform -1 0 35328 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _1062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 36984 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1676037725
transform -1 0 31740 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1064_
timestamp 1676037725
transform 1 0 31188 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1065_
timestamp 1676037725
transform -1 0 37996 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1066_
timestamp 1676037725
transform -1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31648 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1069_
timestamp 1676037725
transform 1 0 32292 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_4  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32108 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__a22o_1  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26404 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1072_
timestamp 1676037725
transform 1 0 15824 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1676037725
transform 1 0 15364 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1676037725
transform -1 0 16928 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 1676037725
transform -1 0 16376 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1676037725
transform -1 0 14812 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1077_
timestamp 1676037725
transform -1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1078_
timestamp 1676037725
transform -1 0 22356 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1079_
timestamp 1676037725
transform 1 0 40388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1080_
timestamp 1676037725
transform 1 0 42780 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1081_
timestamp 1676037725
transform -1 0 43056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41676 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1676037725
transform 1 0 42780 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31740 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1086_
timestamp 1676037725
transform -1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1087_
timestamp 1676037725
transform 1 0 29992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1088_
timestamp 1676037725
transform -1 0 31372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 36248 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1090_
timestamp 1676037725
transform -1 0 36524 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32936 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1092_
timestamp 1676037725
transform -1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34224 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1094_
timestamp 1676037725
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1096_
timestamp 1676037725
transform 1 0 36432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34776 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_2  _1098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33488 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1099_
timestamp 1676037725
transform -1 0 42044 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1676037725
transform -1 0 40388 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1101_
timestamp 1676037725
transform 1 0 33580 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 1676037725
transform -1 0 32568 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32660 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1104_
timestamp 1676037725
transform -1 0 29624 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1105_
timestamp 1676037725
transform -1 0 34500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _1106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34224 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_1  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33856 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 43332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1109_
timestamp 1676037725
transform -1 0 39008 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1676037725
transform 1 0 33856 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34776 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_4  _1112_
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33580 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21344 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1116_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_2  _1117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _1118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _1119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1676037725
transform -1 0 24840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1121_
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _1122_
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16192 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1126_
timestamp 1676037725
transform -1 0 30268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30176 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1128_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1130_
timestamp 1676037725
transform 1 0 24932 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1676037725
transform -1 0 23092 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1676037725
transform -1 0 21528 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1676037725
transform -1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1134_
timestamp 1676037725
transform -1 0 20976 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1676037725
transform 1 0 19872 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1136_
timestamp 1676037725
transform -1 0 14720 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1137_
timestamp 1676037725
transform -1 0 15824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1138_
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1676037725
transform -1 0 28428 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1140_
timestamp 1676037725
transform 1 0 28888 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1141_
timestamp 1676037725
transform 1 0 28704 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1142_
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1143_
timestamp 1676037725
transform 1 0 20056 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1144_
timestamp 1676037725
transform -1 0 14168 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1676037725
transform -1 0 15640 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1146_
timestamp 1676037725
transform -1 0 16008 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1147_
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1148_
timestamp 1676037725
transform -1 0 38548 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1149_
timestamp 1676037725
transform -1 0 30820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1150_
timestamp 1676037725
transform 1 0 23368 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1151_
timestamp 1676037725
transform -1 0 25392 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1152_
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1153_
timestamp 1676037725
transform -1 0 22632 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1154_
timestamp 1676037725
transform -1 0 22816 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1155_
timestamp 1676037725
transform -1 0 22908 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1156_
timestamp 1676037725
transform 1 0 21068 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1157_
timestamp 1676037725
transform 1 0 14996 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1160_
timestamp 1676037725
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1161_
timestamp 1676037725
transform -1 0 16008 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1162_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1163_
timestamp 1676037725
transform -1 0 35512 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1164_
timestamp 1676037725
transform -1 0 31188 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1165_
timestamp 1676037725
transform 1 0 23000 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1166_
timestamp 1676037725
transform -1 0 25668 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1167_
timestamp 1676037725
transform -1 0 24380 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1168_
timestamp 1676037725
transform -1 0 23276 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1169_
timestamp 1676037725
transform -1 0 21528 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1170_
timestamp 1676037725
transform -1 0 21528 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1171_
timestamp 1676037725
transform 1 0 21896 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1172_
timestamp 1676037725
transform -1 0 23828 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1173_
timestamp 1676037725
transform -1 0 22264 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1175_
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _1176_
timestamp 1676037725
transform -1 0 12328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1676037725
transform -1 0 14352 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1676037725
transform 1 0 12696 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_4  _1179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1676037725
transform 1 0 17848 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1181_
timestamp 1676037725
transform -1 0 23184 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1182_
timestamp 1676037725
transform -1 0 22356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 1676037725
transform 1 0 23552 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1184_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1185_
timestamp 1676037725
transform -1 0 24196 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 1676037725
transform -1 0 32384 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1676037725
transform -1 0 31188 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1188_
timestamp 1676037725
transform 1 0 23460 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1189_
timestamp 1676037725
transform -1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1191_
timestamp 1676037725
transform -1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1676037725
transform -1 0 23552 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1194_
timestamp 1676037725
transform 1 0 22356 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1196_
timestamp 1676037725
transform -1 0 30544 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1197_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1198_
timestamp 1676037725
transform 1 0 21804 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1199_
timestamp 1676037725
transform -1 0 19872 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1676037725
transform -1 0 29992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1676037725
transform -1 0 31004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1203_
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1204_
timestamp 1676037725
transform -1 0 29256 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1206_
timestamp 1676037725
transform -1 0 30452 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1207_
timestamp 1676037725
transform -1 0 35236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1208_
timestamp 1676037725
transform -1 0 34776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1676037725
transform 1 0 34868 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1210_
timestamp 1676037725
transform 1 0 33764 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1211_
timestamp 1676037725
transform -1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1212_
timestamp 1676037725
transform -1 0 33212 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1676037725
transform 1 0 29716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1214_
timestamp 1676037725
transform -1 0 29624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1215_
timestamp 1676037725
transform 1 0 17204 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1216_
timestamp 1676037725
transform 1 0 17848 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1217_
timestamp 1676037725
transform 1 0 17296 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1218_
timestamp 1676037725
transform -1 0 17204 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1219_
timestamp 1676037725
transform -1 0 25208 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 1676037725
transform 1 0 16008 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 1676037725
transform -1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1222_
timestamp 1676037725
transform -1 0 20976 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1223_
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1224_
timestamp 1676037725
transform -1 0 20976 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1676037725
transform 1 0 19688 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1226_
timestamp 1676037725
transform -1 0 21344 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1227_
timestamp 1676037725
transform -1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1228_
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1229_
timestamp 1676037725
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1676037725
transform -1 0 22816 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1231_
timestamp 1676037725
transform -1 0 33028 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1232_
timestamp 1676037725
transform -1 0 31280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1233_
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1234_
timestamp 1676037725
transform -1 0 18952 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1235_
timestamp 1676037725
transform 1 0 15640 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1236_
timestamp 1676037725
transform 1 0 15732 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1237_
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1238_
timestamp 1676037725
transform -1 0 24748 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1676037725
transform -1 0 24104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1241_
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1242_
timestamp 1676037725
transform -1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1243_
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1244_
timestamp 1676037725
transform 1 0 21896 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1245_
timestamp 1676037725
transform 1 0 15456 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1676037725
transform -1 0 13984 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1247_
timestamp 1676037725
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1248_
timestamp 1676037725
transform -1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1249_
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1250_
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1251_
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1252_
timestamp 1676037725
transform -1 0 15364 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1254_
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1676037725
transform -1 0 22448 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _1256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1257_
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1676037725
transform -1 0 13340 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1259_
timestamp 1676037725
transform 1 0 13064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13248 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1261_
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1676037725
transform -1 0 16192 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1264_
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 1676037725
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1266_
timestamp 1676037725
transform -1 0 38088 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1267_
timestamp 1676037725
transform 1 0 28612 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28060 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1269_
timestamp 1676037725
transform -1 0 26312 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1270_
timestamp 1676037725
transform 1 0 18400 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1271_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1272_
timestamp 1676037725
transform -1 0 19688 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1273_
timestamp 1676037725
transform 1 0 18676 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1274_
timestamp 1676037725
transform -1 0 18124 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1275_
timestamp 1676037725
transform -1 0 16376 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1276_
timestamp 1676037725
transform -1 0 16284 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1277_
timestamp 1676037725
transform 1 0 16376 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1278_
timestamp 1676037725
transform -1 0 16284 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1279_
timestamp 1676037725
transform -1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14720 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1281_
timestamp 1676037725
transform 1 0 15088 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16192 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1283_
timestamp 1676037725
transform 1 0 12420 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1284_
timestamp 1676037725
transform -1 0 27324 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1285_
timestamp 1676037725
transform 1 0 18584 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1286_
timestamp 1676037725
transform -1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1287_
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1289_
timestamp 1676037725
transform 1 0 17572 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1676037725
transform 1 0 17480 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1291_
timestamp 1676037725
transform 1 0 17112 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1676037725
transform 1 0 17848 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1676037725
transform -1 0 16376 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1294_
timestamp 1676037725
transform -1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1676037725
transform 1 0 16928 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1676037725
transform -1 0 18032 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1297_
timestamp 1676037725
transform 1 0 17756 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1298_
timestamp 1676037725
transform -1 0 18400 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1299_
timestamp 1676037725
transform -1 0 13800 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1300_
timestamp 1676037725
transform 1 0 13616 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1676037725
transform -1 0 15272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16928 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1303_
timestamp 1676037725
transform 1 0 16928 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1676037725
transform -1 0 25484 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1676037725
transform -1 0 23276 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1306_
timestamp 1676037725
transform -1 0 18860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1676037725
transform 1 0 17388 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1308_
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1676037725
transform 1 0 32752 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1310_
timestamp 1676037725
transform 1 0 34868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1311_
timestamp 1676037725
transform -1 0 40296 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1312_
timestamp 1676037725
transform -1 0 40664 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1313_
timestamp 1676037725
transform 1 0 41400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_
timestamp 1676037725
transform 1 0 40664 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1315_
timestamp 1676037725
transform 1 0 40020 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1676037725
transform -1 0 36984 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1317_
timestamp 1676037725
transform -1 0 35972 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1318_
timestamp 1676037725
transform 1 0 35880 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29900 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1321_
timestamp 1676037725
transform 1 0 38916 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1322_
timestamp 1676037725
transform -1 0 36156 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1323_
timestamp 1676037725
transform 1 0 29900 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1324_
timestamp 1676037725
transform 1 0 30452 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1325_
timestamp 1676037725
transform 1 0 39192 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1326_
timestamp 1676037725
transform -1 0 43056 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1327_
timestamp 1676037725
transform -1 0 38456 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1328_
timestamp 1676037725
transform 1 0 27232 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp 1676037725
transform -1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1676037725
transform -1 0 36616 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1331_
timestamp 1676037725
transform 1 0 37444 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1332_
timestamp 1676037725
transform 1 0 29440 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1676037725
transform -1 0 30176 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1676037725
transform -1 0 35328 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34868 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1336_
timestamp 1676037725
transform -1 0 24656 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1337_
timestamp 1676037725
transform -1 0 20608 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1338_
timestamp 1676037725
transform -1 0 20884 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1339_
timestamp 1676037725
transform -1 0 19688 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 1676037725
transform -1 0 38456 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp 1676037725
transform 1 0 36432 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1342_
timestamp 1676037725
transform -1 0 26680 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25484 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1344_
timestamp 1676037725
transform 1 0 20424 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1345_
timestamp 1676037725
transform -1 0 23736 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31832 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1347_
timestamp 1676037725
transform -1 0 25300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1348_
timestamp 1676037725
transform -1 0 24472 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1349_
timestamp 1676037725
transform 1 0 22724 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1350_
timestamp 1676037725
transform 1 0 25300 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1351_
timestamp 1676037725
transform -1 0 25944 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1352_
timestamp 1676037725
transform -1 0 25208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1353_
timestamp 1676037725
transform 1 0 24288 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1354_
timestamp 1676037725
transform 1 0 24840 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1355_
timestamp 1676037725
transform -1 0 26956 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1356_
timestamp 1676037725
transform 1 0 26312 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1357_
timestamp 1676037725
transform 1 0 26220 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1358_
timestamp 1676037725
transform 1 0 27232 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1359_
timestamp 1676037725
transform 1 0 27968 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1360_
timestamp 1676037725
transform 1 0 28980 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1361_
timestamp 1676037725
transform 1 0 28060 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1676037725
transform 1 0 28704 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1363_
timestamp 1676037725
transform 1 0 34868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1364_
timestamp 1676037725
transform -1 0 32476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1365_
timestamp 1676037725
transform -1 0 31188 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1366_
timestamp 1676037725
transform -1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1367_
timestamp 1676037725
transform 1 0 30636 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1676037725
transform 1 0 31556 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1369_
timestamp 1676037725
transform 1 0 34868 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1370_
timestamp 1676037725
transform 1 0 34868 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1371_
timestamp 1676037725
transform 1 0 35788 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1372_
timestamp 1676037725
transform 1 0 35972 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1373_
timestamp 1676037725
transform 1 0 33672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1374_
timestamp 1676037725
transform 1 0 34960 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1375_
timestamp 1676037725
transform 1 0 34868 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1376_
timestamp 1676037725
transform 1 0 33856 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1377_
timestamp 1676037725
transform 1 0 35144 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1378_
timestamp 1676037725
transform 1 0 35880 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1379_
timestamp 1676037725
transform 1 0 36708 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1676037725
transform -1 0 36984 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1381_
timestamp 1676037725
transform 1 0 33580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1382_
timestamp 1676037725
transform 1 0 40020 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1383_
timestamp 1676037725
transform 1 0 38916 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1676037725
transform 1 0 34868 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1385_
timestamp 1676037725
transform 1 0 40020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1386_
timestamp 1676037725
transform 1 0 40020 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1387_
timestamp 1676037725
transform -1 0 40388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1388_
timestamp 1676037725
transform 1 0 41032 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1389_
timestamp 1676037725
transform 1 0 36708 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1390_
timestamp 1676037725
transform 1 0 40020 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1391_
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1392_
timestamp 1676037725
transform 1 0 37812 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1676037725
transform 1 0 40112 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1394_
timestamp 1676037725
transform 1 0 41124 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1395_
timestamp 1676037725
transform -1 0 41492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1676037725
transform -1 0 42136 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1397_
timestamp 1676037725
transform 1 0 37076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1398_
timestamp 1676037725
transform 1 0 40480 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1399_
timestamp 1676037725
transform 1 0 41216 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1676037725
transform 1 0 41124 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1401_
timestamp 1676037725
transform 1 0 41584 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1402_
timestamp 1676037725
transform 1 0 42596 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1403_
timestamp 1676037725
transform 1 0 37444 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1404_
timestamp 1676037725
transform 1 0 39376 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1405_
timestamp 1676037725
transform 1 0 40480 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1406_
timestamp 1676037725
transform -1 0 13524 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1407_
timestamp 1676037725
transform -1 0 12696 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1408_
timestamp 1676037725
transform -1 0 12328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1409_
timestamp 1676037725
transform 1 0 12696 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1676037725
transform -1 0 13800 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1411_
timestamp 1676037725
transform -1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1414_
timestamp 1676037725
transform 1 0 41032 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1415_
timestamp 1676037725
transform -1 0 39376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1416_
timestamp 1676037725
transform 1 0 39284 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1417_
timestamp 1676037725
transform -1 0 38364 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1418_
timestamp 1676037725
transform -1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1419_
timestamp 1676037725
transform 1 0 40480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1420_
timestamp 1676037725
transform -1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1421_
timestamp 1676037725
transform -1 0 36708 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1422_
timestamp 1676037725
transform 1 0 42596 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1423_
timestamp 1676037725
transform -1 0 38732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1424_
timestamp 1676037725
transform 1 0 42596 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1425_
timestamp 1676037725
transform -1 0 38272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1426_
timestamp 1676037725
transform 1 0 36800 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1427_
timestamp 1676037725
transform -1 0 40572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1428_
timestamp 1676037725
transform -1 0 39100 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1429_
timestamp 1676037725
transform -1 0 36708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1430_
timestamp 1676037725
transform 1 0 36432 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1431_
timestamp 1676037725
transform 1 0 36340 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1432_
timestamp 1676037725
transform -1 0 39560 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1433_
timestamp 1676037725
transform 1 0 38916 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1434_
timestamp 1676037725
transform 1 0 39008 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1435_
timestamp 1676037725
transform -1 0 36984 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1437_
timestamp 1676037725
transform -1 0 35420 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1438_
timestamp 1676037725
transform -1 0 38732 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1440_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1441_
timestamp 1676037725
transform -1 0 39100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1442_
timestamp 1676037725
transform -1 0 38456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1443_
timestamp 1676037725
transform -1 0 39836 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1444_
timestamp 1676037725
transform -1 0 36984 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1445_
timestamp 1676037725
transform 1 0 36432 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1446_
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1447_
timestamp 1676037725
transform -1 0 34408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1448_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1449_
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1450_
timestamp 1676037725
transform -1 0 35328 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1452_
timestamp 1676037725
transform 1 0 38640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1453_
timestamp 1676037725
transform 1 0 35696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1454_
timestamp 1676037725
transform 1 0 40664 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1455_
timestamp 1676037725
transform 1 0 37076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1456_
timestamp 1676037725
transform 1 0 37444 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1457_
timestamp 1676037725
transform -1 0 37720 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1458_
timestamp 1676037725
transform 1 0 38088 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1459_
timestamp 1676037725
transform -1 0 40204 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1460_
timestamp 1676037725
transform 1 0 38732 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1461_
timestamp 1676037725
transform 1 0 37720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1462_
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1463_
timestamp 1676037725
transform -1 0 38456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1464_
timestamp 1676037725
transform 1 0 37628 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1676037725
transform -1 0 40296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1466_
timestamp 1676037725
transform -1 0 35236 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1676037725
transform -1 0 35880 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1468_
timestamp 1676037725
transform -1 0 36340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1469_
timestamp 1676037725
transform -1 0 35696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1470_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1471_
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1472_
timestamp 1676037725
transform 1 0 38916 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1473_
timestamp 1676037725
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1474_
timestamp 1676037725
transform -1 0 38732 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1475_
timestamp 1676037725
transform -1 0 37996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1476_
timestamp 1676037725
transform -1 0 37628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1477_
timestamp 1676037725
transform 1 0 37536 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1479_
timestamp 1676037725
transform 1 0 28336 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1480_
timestamp 1676037725
transform -1 0 33580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1481_
timestamp 1676037725
transform -1 0 34408 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1482_
timestamp 1676037725
transform -1 0 34684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1483_
timestamp 1676037725
transform -1 0 35604 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1676037725
transform 1 0 35972 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1485_
timestamp 1676037725
transform -1 0 39284 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 39284 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1487_
timestamp 1676037725
transform 1 0 37904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1488_
timestamp 1676037725
transform -1 0 37536 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1489_
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1490_
timestamp 1676037725
transform -1 0 38180 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1492_
timestamp 1676037725
transform 1 0 39100 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1676037725
transform -1 0 37536 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1494_
timestamp 1676037725
transform -1 0 38272 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1495_
timestamp 1676037725
transform -1 0 38732 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1676037725
transform 1 0 37904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1497_
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1498_
timestamp 1676037725
transform 1 0 34408 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1500_
timestamp 1676037725
transform -1 0 39284 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1501_
timestamp 1676037725
transform -1 0 38272 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1502_
timestamp 1676037725
transform -1 0 36892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1503_
timestamp 1676037725
transform -1 0 37904 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1504_
timestamp 1676037725
transform -1 0 36984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1505_
timestamp 1676037725
transform 1 0 36064 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1506_
timestamp 1676037725
transform -1 0 37076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1507_
timestamp 1676037725
transform 1 0 37444 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1508_
timestamp 1676037725
transform 1 0 38732 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1509_
timestamp 1676037725
transform 1 0 40020 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1676037725
transform 1 0 40020 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1513_
timestamp 1676037725
transform 1 0 38916 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1676037725
transform 1 0 35236 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1515_
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1516_
timestamp 1676037725
transform -1 0 38180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1517_
timestamp 1676037725
transform 1 0 37628 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1518_
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1676037725
transform 1 0 40664 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1676037725
transform -1 0 40112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1521_
timestamp 1676037725
transform -1 0 36984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1522_
timestamp 1676037725
transform 1 0 38640 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1523_
timestamp 1676037725
transform -1 0 39284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1524_
timestamp 1676037725
transform 1 0 38548 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1525_
timestamp 1676037725
transform 1 0 38824 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1526_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1676037725
transform -1 0 40296 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1528_
timestamp 1676037725
transform -1 0 38732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1529_
timestamp 1676037725
transform 1 0 36432 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1530_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1531_
timestamp 1676037725
transform 1 0 39192 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1532_
timestamp 1676037725
transform -1 0 41124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1676037725
transform 1 0 40020 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1534_
timestamp 1676037725
transform -1 0 40112 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1535_
timestamp 1676037725
transform -1 0 32660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 1676037725
transform 1 0 36616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1537_
timestamp 1676037725
transform 1 0 36800 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1538_
timestamp 1676037725
transform -1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1539_
timestamp 1676037725
transform -1 0 38732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1540_
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1676037725
transform 1 0 42596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1676037725
transform 1 0 39652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1543_
timestamp 1676037725
transform -1 0 39468 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1545_
timestamp 1676037725
transform 1 0 35604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1546_
timestamp 1676037725
transform 1 0 39192 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1547_
timestamp 1676037725
transform 1 0 39100 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1548_
timestamp 1676037725
transform 1 0 39008 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1676037725
transform -1 0 41124 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1551_
timestamp 1676037725
transform -1 0 38180 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1552_
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1553_
timestamp 1676037725
transform -1 0 31832 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _1554_
timestamp 1676037725
transform 1 0 40112 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_4  _1555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38548 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1556_
timestamp 1676037725
transform 1 0 37352 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 1676037725
transform -1 0 39560 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1558_
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 38272 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _1560_
timestamp 1676037725
transform 1 0 36708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1561_
timestamp 1676037725
transform -1 0 31280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1676037725
transform -1 0 24104 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1563_
timestamp 1676037725
transform 1 0 32752 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _1564_
timestamp 1676037725
transform -1 0 32108 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1565_
timestamp 1676037725
transform -1 0 32844 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _1566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23552 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__a2bb2o_1  _1567_
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 35904
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_1  _1569_
timestamp 1676037725
transform 1 0 23368 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1570_
timestamp 1676037725
transform 1 0 28060 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1571_
timestamp 1676037725
transform -1 0 24012 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1572_
timestamp 1676037725
transform -1 0 22724 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1573_
timestamp 1676037725
transform 1 0 21620 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1575_
timestamp 1676037725
transform -1 0 22724 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1576_
timestamp 1676037725
transform 1 0 21896 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1577_
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1578_
timestamp 1676037725
transform 1 0 20700 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1579_
timestamp 1676037725
transform -1 0 22816 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1580_
timestamp 1676037725
transform 1 0 21804 0 1 38080
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1581_
timestamp 1676037725
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1582_
timestamp 1676037725
transform -1 0 24104 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1583_
timestamp 1676037725
transform 1 0 23552 0 -1 38080
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1584_
timestamp 1676037725
transform 1 0 25760 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1585_
timestamp 1676037725
transform 1 0 27140 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1586_
timestamp 1676037725
transform 1 0 25944 0 1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1587_
timestamp 1676037725
transform 1 0 27232 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1588_
timestamp 1676037725
transform -1 0 28520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1589_
timestamp 1676037725
transform 1 0 27600 0 1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _1590_
timestamp 1676037725
transform 1 0 28336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1591_
timestamp 1676037725
transform -1 0 29256 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1592_
timestamp 1676037725
transform 1 0 28244 0 -1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_1  _1593_
timestamp 1676037725
transform 1 0 33304 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1594_
timestamp 1676037725
transform -1 0 33948 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1595_
timestamp 1676037725
transform -1 0 32936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1596_
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1597_
timestamp 1676037725
transform 1 0 32660 0 1 38080
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _1598_
timestamp 1676037725
transform 1 0 32476 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1599_
timestamp 1676037725
transform 1 0 32292 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31188 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1601_
timestamp 1676037725
transform 1 0 31188 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1602_
timestamp 1676037725
transform 1 0 32844 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1676037725
transform 1 0 34868 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1604_
timestamp 1676037725
transform 1 0 34776 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1676037725
transform 1 0 36248 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1606_
timestamp 1676037725
transform 1 0 36524 0 1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1676037725
transform 1 0 36340 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1608_
timestamp 1676037725
transform 1 0 37352 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1676037725
transform 1 0 36340 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1610_
timestamp 1676037725
transform -1 0 39652 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1676037725
transform -1 0 39560 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1612_
timestamp 1676037725
transform -1 0 39744 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1676037725
transform -1 0 27968 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32108 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1615_
timestamp 1676037725
transform -1 0 27784 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _1616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1617_
timestamp 1676037725
transform -1 0 25668 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1618_
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_4  _1619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _1620_
timestamp 1676037725
transform -1 0 25484 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1621_
timestamp 1676037725
transform -1 0 27232 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1676037725
transform -1 0 25576 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1624_
timestamp 1676037725
transform -1 0 33120 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1625_
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_4  _1626_
timestamp 1676037725
transform 1 0 24840 0 -1 34816
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1676037725
transform -1 0 27692 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1628_
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _1629_
timestamp 1676037725
transform -1 0 21528 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__o21a_1  _1630_
timestamp 1676037725
transform -1 0 34500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1631_
timestamp 1676037725
transform -1 0 33580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1632_
timestamp 1676037725
transform 1 0 33488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1633_
timestamp 1676037725
transform 1 0 33764 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1634_
timestamp 1676037725
transform -1 0 21528 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1636_
timestamp 1676037725
transform 1 0 30360 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1676037725
transform -1 0 30360 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1638_
timestamp 1676037725
transform -1 0 29440 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1639_
timestamp 1676037725
transform -1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1640_
timestamp 1676037725
transform 1 0 26496 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1641_
timestamp 1676037725
transform -1 0 28244 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26312 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1643_
timestamp 1676037725
transform -1 0 30360 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1644_
timestamp 1676037725
transform 1 0 28060 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1645_
timestamp 1676037725
transform 1 0 27324 0 -1 34816
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1646_
timestamp 1676037725
transform -1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1647_
timestamp 1676037725
transform -1 0 43056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1648_
timestamp 1676037725
transform -1 0 42872 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1650_
timestamp 1676037725
transform -1 0 42872 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1651_
timestamp 1676037725
transform -1 0 42872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1652_
timestamp 1676037725
transform -1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1653_
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1654_
timestamp 1676037725
transform -1 0 31188 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1655_
timestamp 1676037725
transform 1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1656_
timestamp 1676037725
transform -1 0 19964 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1657_
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1658_
timestamp 1676037725
transform 1 0 22448 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1676037725
transform -1 0 22724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1660_
timestamp 1676037725
transform -1 0 21896 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1661_
timestamp 1676037725
transform -1 0 22540 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1662_
timestamp 1676037725
transform -1 0 21528 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1663_
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1664_
timestamp 1676037725
transform -1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1665_
timestamp 1676037725
transform 1 0 22356 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1666_
timestamp 1676037725
transform -1 0 22632 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1676037725
transform -1 0 23460 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1676037725
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 1676037725
transform -1 0 21160 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1670_
timestamp 1676037725
transform -1 0 20240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1671_
timestamp 1676037725
transform -1 0 19872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1672_
timestamp 1676037725
transform 1 0 21344 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1673_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1675_
timestamp 1676037725
transform -1 0 18952 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1676_
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1677_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1678_
timestamp 1676037725
transform 1 0 20424 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1681_
timestamp 1676037725
transform -1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1682_
timestamp 1676037725
transform 1 0 20056 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1676037725
transform -1 0 12604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1685_
timestamp 1676037725
transform 1 0 22724 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1686_
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1687_
timestamp 1676037725
transform -1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1688_
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1689_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1690_
timestamp 1676037725
transform -1 0 25300 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1676037725
transform -1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1693_
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1694_
timestamp 1676037725
transform -1 0 23276 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1695_
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1696_
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1697_
timestamp 1676037725
transform 1 0 23644 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1698_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1676037725
transform 1 0 13432 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1700_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1701_
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1703_
timestamp 1676037725
transform -1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26496 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1707_
timestamp 1676037725
transform -1 0 19872 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1708_
timestamp 1676037725
transform -1 0 19688 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1676037725
transform -1 0 21528 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1676037725
transform -1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1676037725
transform -1 0 20516 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1715_
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1716_
timestamp 1676037725
transform -1 0 17388 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1676037725
transform 1 0 15548 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 1676037725
transform -1 0 18676 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1676037725
transform -1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 1676037725
transform 1 0 17664 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1676037725
transform 1 0 17480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1725_
timestamp 1676037725
transform 1 0 41032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1726_
timestamp 1676037725
transform -1 0 39468 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1727_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1728_
timestamp 1676037725
transform 1 0 35236 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1729_
timestamp 1676037725
transform -1 0 33212 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1730_
timestamp 1676037725
transform 1 0 35512 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1731_
timestamp 1676037725
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1732_
timestamp 1676037725
transform 1 0 35052 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1733_
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1734_
timestamp 1676037725
transform -1 0 38364 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1735_
timestamp 1676037725
transform -1 0 36984 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1736_
timestamp 1676037725
transform -1 0 35788 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1737_
timestamp 1676037725
transform 1 0 33396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1739_
timestamp 1676037725
transform 1 0 19412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1741_
timestamp 1676037725
transform 1 0 18216 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 1676037725
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1743_
timestamp 1676037725
transform 1 0 19412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1676037725
transform 1 0 20700 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1745_
timestamp 1676037725
transform 1 0 20424 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1676037725
transform 1 0 22540 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1676037725
transform 1 0 25300 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1676037725
transform 1 0 25208 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1676037725
transform 1 0 27140 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1676037725
transform 1 0 27140 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1676037725
transform -1 0 29164 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1676037725
transform -1 0 28980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1754_
timestamp 1676037725
transform -1 0 31096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 1676037725
transform 1 0 30360 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1756_
timestamp 1676037725
transform 1 0 28704 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 1676037725
transform -1 0 30360 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1759_
timestamp 1676037725
transform 1 0 31280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1760_
timestamp 1676037725
transform -1 0 31280 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1761_
timestamp 1676037725
transform 1 0 30912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1762_
timestamp 1676037725
transform -1 0 34040 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1763_
timestamp 1676037725
transform 1 0 29716 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1765_
timestamp 1676037725
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1766_
timestamp 1676037725
transform 1 0 26220 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1767_
timestamp 1676037725
transform 1 0 25760 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1768_
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1676037725
transform 1 0 27876 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1676037725
transform 1 0 26680 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1772_
timestamp 1676037725
transform -1 0 24012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1773_
timestamp 1676037725
transform 1 0 27232 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1774_
timestamp 1676037725
transform 1 0 27324 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1676037725
transform 1 0 25668 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1776_
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1676037725
transform 1 0 28336 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1778_
timestamp 1676037725
transform 1 0 27876 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1779_
timestamp 1676037725
transform 1 0 27324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1781_
timestamp 1676037725
transform -1 0 26680 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1782_
timestamp 1676037725
transform -1 0 29440 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1676037725
transform -1 0 27784 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1785_
timestamp 1676037725
transform -1 0 32108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1786_
timestamp 1676037725
transform -1 0 28704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1787_
timestamp 1676037725
transform 1 0 28152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 1676037725
transform 1 0 25300 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1789_
timestamp 1676037725
transform 1 0 24656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1790_
timestamp 1676037725
transform -1 0 32476 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1676037725
transform 1 0 31004 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1676037725
transform 1 0 30544 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1793_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1794_
timestamp 1676037725
transform 1 0 31188 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1676037725
transform 1 0 30084 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1796_
timestamp 1676037725
transform -1 0 30452 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1797_
timestamp 1676037725
transform -1 0 29808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1798_
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1799_
timestamp 1676037725
transform 1 0 18308 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1800_
timestamp 1676037725
transform 1 0 19320 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1801_
timestamp 1676037725
transform 1 0 19504 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1802_
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1803_
timestamp 1676037725
transform 1 0 27140 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1804_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 1676037725
transform 1 0 25944 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1806_
timestamp 1676037725
transform -1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1807_
timestamp 1676037725
transform 1 0 40756 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1808_
timestamp 1676037725
transform 1 0 41124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 1676037725
transform -1 0 39560 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1810_
timestamp 1676037725
transform 1 0 39192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 1676037725
transform 1 0 40664 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1812_
timestamp 1676037725
transform 1 0 40664 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1676037725
transform 1 0 42320 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1814_
timestamp 1676037725
transform -1 0 42136 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 1676037725
transform 1 0 42596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1816_
timestamp 1676037725
transform -1 0 42136 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 1676037725
transform -1 0 43056 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1818_
timestamp 1676037725
transform 1 0 42596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1676037725
transform 1 0 40756 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1820_
timestamp 1676037725
transform -1 0 39560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1821_
timestamp 1676037725
transform 1 0 42596 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1822_
timestamp 1676037725
transform 1 0 41308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1823_
timestamp 1676037725
transform 1 0 42596 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1824_
timestamp 1676037725
transform 1 0 42412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1825_
timestamp 1676037725
transform -1 0 40388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1826_
timestamp 1676037725
transform 1 0 40112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1827_
timestamp 1676037725
transform -1 0 41032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1828_
timestamp 1676037725
transform -1 0 39560 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1829_
timestamp 1676037725
transform -1 0 33672 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1830_
timestamp 1676037725
transform 1 0 33764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1831_
timestamp 1676037725
transform -1 0 35328 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1832_
timestamp 1676037725
transform 1 0 33580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1833_
timestamp 1676037725
transform -1 0 33212 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1834_
timestamp 1676037725
transform -1 0 32752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1835_
timestamp 1676037725
transform -1 0 35328 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1836_
timestamp 1676037725
transform -1 0 34408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1837_
timestamp 1676037725
transform -1 0 31832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1838_
timestamp 1676037725
transform -1 0 32752 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1839_
timestamp 1676037725
transform -1 0 33764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1840_
timestamp 1676037725
transform -1 0 35328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1841_
timestamp 1676037725
transform -1 0 34960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1842_
timestamp 1676037725
transform -1 0 34776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1843_
timestamp 1676037725
transform -1 0 34408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1844_
timestamp 1676037725
transform -1 0 32752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1845_
timestamp 1676037725
transform 1 0 26036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 1676037725
transform 1 0 25576 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1847_
timestamp 1676037725
transform 1 0 25392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1848_
timestamp 1676037725
transform -1 0 40572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1849_
timestamp 1676037725
transform 1 0 38916 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1850_
timestamp 1676037725
transform -1 0 31832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33120 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1852_
timestamp 1676037725
transform -1 0 33028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1853_
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1854_
timestamp 1676037725
transform 1 0 32568 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1855_
timestamp 1676037725
transform -1 0 31832 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1856_
timestamp 1676037725
transform 1 0 36984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1857_
timestamp 1676037725
transform -1 0 29992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1858_
timestamp 1676037725
transform -1 0 31188 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1859_
timestamp 1676037725
transform 1 0 30360 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1860_
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1861_
timestamp 1676037725
transform -1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1862_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1863_
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1864_
timestamp 1676037725
transform 1 0 32476 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1865_
timestamp 1676037725
transform 1 0 30728 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1866_
timestamp 1676037725
transform 1 0 30544 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1867_
timestamp 1676037725
transform -1 0 34040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1868_
timestamp 1676037725
transform 1 0 36248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1869_
timestamp 1676037725
transform -1 0 35052 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1870_
timestamp 1676037725
transform 1 0 32384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1871_
timestamp 1676037725
transform -1 0 36064 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1872_
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1873_
timestamp 1676037725
transform -1 0 35236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1874_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1875_
timestamp 1676037725
transform 1 0 33856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1876_
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1877_
timestamp 1676037725
transform 1 0 34408 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1878_
timestamp 1676037725
transform -1 0 34408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1879_
timestamp 1676037725
transform -1 0 31832 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1880_
timestamp 1676037725
transform 1 0 30084 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1881_
timestamp 1676037725
transform 1 0 28980 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1882_
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1883_
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1884_
timestamp 1676037725
transform 1 0 29808 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1885_
timestamp 1676037725
transform 1 0 29072 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 35512 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1887_
timestamp 1676037725
transform 1 0 28980 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1888_
timestamp 1676037725
transform -1 0 28152 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1889_
timestamp 1676037725
transform -1 0 30820 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 1676037725
transform -1 0 29256 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1891_
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1892_
timestamp 1676037725
transform -1 0 26036 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1893_
timestamp 1676037725
transform -1 0 33764 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1894_
timestamp 1676037725
transform 1 0 28520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1895_
timestamp 1676037725
transform -1 0 28152 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1896_
timestamp 1676037725
transform -1 0 33396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1897_
timestamp 1676037725
transform 1 0 24840 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1898_
timestamp 1676037725
transform -1 0 24472 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1899_
timestamp 1676037725
transform -1 0 30360 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1900_
timestamp 1676037725
transform -1 0 28152 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1901_
timestamp 1676037725
transform -1 0 26956 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1902_
timestamp 1676037725
transform -1 0 29256 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1903_
timestamp 1676037725
transform 1 0 30084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1904_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _1905_
timestamp 1676037725
transform -1 0 34684 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1906_
timestamp 1676037725
transform 1 0 31464 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1907_
timestamp 1676037725
transform -1 0 29992 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1908_
timestamp 1676037725
transform -1 0 31096 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1909_
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1910_
timestamp 1676037725
transform 1 0 25300 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1911_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1912_
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1913_
timestamp 1676037725
transform 1 0 39928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1914_
timestamp 1676037725
transform -1 0 28060 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1915_
timestamp 1676037725
transform 1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1916_
timestamp 1676037725
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1917_
timestamp 1676037725
transform -1 0 26680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1918_
timestamp 1676037725
transform 1 0 26772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1919_
timestamp 1676037725
transform -1 0 32844 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1920_
timestamp 1676037725
transform -1 0 32568 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1921_
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1922_
timestamp 1676037725
transform -1 0 32016 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1923_
timestamp 1676037725
transform 1 0 31188 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1924_
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1925_
timestamp 1676037725
transform -1 0 29624 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1926_
timestamp 1676037725
transform 1 0 28612 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1927_
timestamp 1676037725
transform -1 0 30452 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1928_
timestamp 1676037725
transform 1 0 33672 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1929_
timestamp 1676037725
transform -1 0 31004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1930_
timestamp 1676037725
transform -1 0 42136 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1931_
timestamp 1676037725
transform 1 0 38640 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1932_
timestamp 1676037725
transform -1 0 32292 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 1676037725
transform -1 0 32568 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1934_
timestamp 1676037725
transform 1 0 30636 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1935_
timestamp 1676037725
transform -1 0 30912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1936_
timestamp 1676037725
transform -1 0 33672 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1937_
timestamp 1676037725
transform 1 0 34040 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1938_
timestamp 1676037725
transform -1 0 35144 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1939_
timestamp 1676037725
transform -1 0 35144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1940_
timestamp 1676037725
transform -1 0 36984 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1941_
timestamp 1676037725
transform 1 0 36708 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1942_
timestamp 1676037725
transform 1 0 37352 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1943_
timestamp 1676037725
transform -1 0 37720 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1944_
timestamp 1676037725
transform 1 0 38548 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1945_
timestamp 1676037725
transform -1 0 38916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1946_
timestamp 1676037725
transform -1 0 40848 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1947_
timestamp 1676037725
transform -1 0 41400 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1948_
timestamp 1676037725
transform 1 0 20056 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1949_
timestamp 1676037725
transform -1 0 20424 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1950_
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1951_
timestamp 1676037725
transform -1 0 21528 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1952_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1953_
timestamp 1676037725
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1954_
timestamp 1676037725
transform -1 0 19596 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1955_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1956_
timestamp 1676037725
transform 1 0 14260 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1957_
timestamp 1676037725
transform -1 0 13892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1958_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1959_
timestamp 1676037725
transform -1 0 13156 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1960_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1961_
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1962_
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1963_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1964_
timestamp 1676037725
transform 1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1965_
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1966_
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1967_
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1968_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1969_
timestamp 1676037725
transform -1 0 19780 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1970_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1971_
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1972_
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1973_
timestamp 1676037725
transform -1 0 19688 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1974_
timestamp 1676037725
transform 1 0 16192 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1975_
timestamp 1676037725
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1976_
timestamp 1676037725
transform 1 0 15548 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1977_
timestamp 1676037725
transform -1 0 15456 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1978_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1979_
timestamp 1676037725
transform -1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1980_
timestamp 1676037725
transform -1 0 18676 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1981_
timestamp 1676037725
transform 1 0 18584 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1982_
timestamp 1676037725
transform 1 0 17020 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1983_
timestamp 1676037725
transform -1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40204 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1985_
timestamp 1676037725
transform 1 0 41492 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40296 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41400 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1988_
timestamp 1676037725
transform -1 0 43240 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41308 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1676037725
transform -1 0 24012 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1676037725
transform 1 0 13340 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1994_
timestamp 1676037725
transform 1 0 13340 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1995_
timestamp 1676037725
transform 1 0 13248 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1996_
timestamp 1676037725
transform 1 0 13248 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1997_
timestamp 1676037725
transform 1 0 13432 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1998_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1999_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2000_
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2001_
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2002_
timestamp 1676037725
transform 1 0 15272 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2003_
timestamp 1676037725
transform -1 0 18860 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2004_
timestamp 1676037725
transform 1 0 17204 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2005_
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _2006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 -1 34816
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2007_
timestamp 1676037725
transform 1 0 18400 0 -1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _2008_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _2010_
timestamp 1676037725
transform 1 0 14628 0 -1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2011_
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2012_
timestamp 1676037725
transform 1 0 13800 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _2013_
timestamp 1676037725
transform 1 0 14260 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2014_
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _2015_
timestamp 1676037725
transform 1 0 16192 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _2016_
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2017_
timestamp 1676037725
transform 1 0 16836 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2018_
timestamp 1676037725
transform 1 0 29900 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2019_
timestamp 1676037725
transform 1 0 20056 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2020_
timestamp 1676037725
transform 1 0 20976 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1676037725
transform -1 0 24104 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1676037725
transform 1 0 25024 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2023_
timestamp 1676037725
transform 1 0 27140 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2024_
timestamp 1676037725
transform 1 0 28428 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2025_
timestamp 1676037725
transform -1 0 31740 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2026_
timestamp 1676037725
transform -1 0 36800 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2027_
timestamp 1676037725
transform -1 0 38916 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2028_
timestamp 1676037725
transform 1 0 40020 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2029_
timestamp 1676037725
transform 1 0 41860 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2030_
timestamp 1676037725
transform 1 0 41952 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2031_
timestamp 1676037725
transform 1 0 41860 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2032_
timestamp 1676037725
transform 1 0 41952 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2033_
timestamp 1676037725
transform 1 0 41492 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2034_
timestamp 1676037725
transform 1 0 18768 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2035_
timestamp 1676037725
transform 1 0 17480 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2036_
timestamp 1676037725
transform 1 0 18492 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2037_
timestamp 1676037725
transform 1 0 19964 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2038_
timestamp 1676037725
transform 1 0 22264 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2039_
timestamp 1676037725
transform 1 0 25024 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2040_
timestamp 1676037725
transform 1 0 26864 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2041_
timestamp 1676037725
transform 1 0 29716 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2042_
timestamp 1676037725
transform -1 0 29256 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2043_
timestamp 1676037725
transform -1 0 23828 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2044_
timestamp 1676037725
transform 1 0 26128 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2045_
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2046_
timestamp 1676037725
transform 1 0 27140 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2047_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2048_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2049_
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2050_
timestamp 1676037725
transform 1 0 38732 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2051_
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2052_
timestamp 1676037725
transform 1 0 41952 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2053_
timestamp 1676037725
transform 1 0 41860 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2054_
timestamp 1676037725
transform 1 0 41952 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2055_
timestamp 1676037725
transform 1 0 40020 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2056_
timestamp 1676037725
transform 1 0 40664 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2057_
timestamp 1676037725
transform 1 0 41952 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2058_
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2059_
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2060_
timestamp 1676037725
transform -1 0 39928 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2061_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2062_
timestamp 1676037725
transform 1 0 30360 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2063_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2064_
timestamp 1676037725
transform -1 0 33672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2065_
timestamp 1676037725
transform 1 0 33580 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2066_
timestamp 1676037725
transform 1 0 35144 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2067_
timestamp 1676037725
transform 1 0 29532 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2068_
timestamp 1676037725
transform 1 0 27784 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2069_
timestamp 1676037725
transform -1 0 29900 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2070_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2071_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2072_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2073_
timestamp 1676037725
transform -1 0 28612 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2074_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2075_
timestamp 1676037725
transform 1 0 28520 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2076_
timestamp 1676037725
transform -1 0 26036 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2077_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2078_
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2079_
timestamp 1676037725
transform -1 0 26496 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2080_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2081_
timestamp 1676037725
transform 1 0 25852 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2082_
timestamp 1676037725
transform -1 0 33120 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2083_
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2084_
timestamp 1676037725
transform -1 0 28612 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2085_
timestamp 1676037725
transform 1 0 26680 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2086_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2087_
timestamp 1676037725
transform 1 0 29624 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2088_
timestamp 1676037725
transform 1 0 33764 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2089_
timestamp 1676037725
transform -1 0 31556 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2090_
timestamp 1676037725
transform 1 0 27324 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2091_
timestamp 1676037725
transform 1 0 25208 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2092_
timestamp 1676037725
transform 1 0 24840 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2093_
timestamp 1676037725
transform -1 0 43332 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2094_
timestamp 1676037725
transform 1 0 40020 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2095_
timestamp 1676037725
transform 1 0 32292 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2096_
timestamp 1676037725
transform 1 0 31556 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2097_
timestamp 1676037725
transform -1 0 34132 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2098_
timestamp 1676037725
transform -1 0 36340 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2099_
timestamp 1676037725
transform 1 0 35512 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2100_
timestamp 1676037725
transform 1 0 37444 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2101_
timestamp 1676037725
transform 1 0 39284 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2102_
timestamp 1676037725
transform -1 0 41492 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2103_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2104_
timestamp 1676037725
transform 1 0 20792 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2105_
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2106_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2107_
timestamp 1676037725
transform 1 0 13524 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2108_
timestamp 1676037725
transform 1 0 13432 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2109_
timestamp 1676037725
transform 1 0 13432 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2110_
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2111_
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2112_
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2113_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2114_
timestamp 1676037725
transform 1 0 15824 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2115_
timestamp 1676037725
transform 1 0 15548 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2116_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2117_
timestamp 1676037725
transform -1 0 18860 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2118_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30176 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21528 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform 1 0 23092 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform -1 0 21344 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform -1 0 29072 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform -1 0 30820 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform 1 0 32384 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform 1 0 33028 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform -1 0 24012 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform -1 0 24288 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform -1 0 26128 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 35144 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform 1 0 35052 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform -1 0 34684 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1676037725
transform -1 0 43424 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1676037725
transform -1 0 43424 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1676037725
transform -1 0 43424 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1676037725
transform -1 0 43424 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1676037725
transform -1 0 42136 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1676037725
transform -1 0 43424 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform -1 0 43424 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1676037725
transform -1 0 43424 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1676037725
transform 1 0 42504 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 43148 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1676037725
transform -1 0 43424 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14536 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_13
timestamp 1676037725
transform -1 0 15732 0 -1 42432
box -38 -48 314 592
<< labels >>
flabel metal3 s 44200 38844 45000 39084 0 FreeSans 960 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 44200 2124 45000 2364 0 FreeSans 960 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 44200 5796 45000 6036 0 FreeSans 960 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 44200 9468 45000 9708 0 FreeSans 960 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 44200 13140 45000 13380 0 FreeSans 960 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 44200 16812 45000 17052 0 FreeSans 960 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 44200 20484 45000 20724 0 FreeSans 960 0 0 0 io_in[5]
port 6 nsew signal input
flabel metal3 s 44200 24156 45000 24396 0 FreeSans 960 0 0 0 io_in[6]
port 7 nsew signal input
flabel metal3 s 44200 27828 45000 28068 0 FreeSans 960 0 0 0 io_in[7]
port 8 nsew signal input
flabel metal3 s 44200 31500 45000 31740 0 FreeSans 960 0 0 0 io_in[8]
port 9 nsew signal input
flabel metal3 s 44200 35172 45000 35412 0 FreeSans 960 0 0 0 io_in[9]
port 10 nsew signal input
flabel metal2 s 43506 44200 43618 45000 0 FreeSans 448 90 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 1278 44200 1390 45000 0 FreeSans 448 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 16918 44200 17030 45000 0 FreeSans 448 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 18482 44200 18594 45000 0 FreeSans 448 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 20046 44200 20158 45000 0 FreeSans 448 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 21610 44200 21722 45000 0 FreeSans 448 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 23174 44200 23286 45000 0 FreeSans 448 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 24738 44200 24850 45000 0 FreeSans 448 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 26302 44200 26414 45000 0 FreeSans 448 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 27866 44200 27978 45000 0 FreeSans 448 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 29430 44200 29542 45000 0 FreeSans 448 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 30994 44200 31106 45000 0 FreeSans 448 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 2842 44200 2954 45000 0 FreeSans 448 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 32558 44200 32670 45000 0 FreeSans 448 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 34122 44200 34234 45000 0 FreeSans 448 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 35686 44200 35798 45000 0 FreeSans 448 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 37250 44200 37362 45000 0 FreeSans 448 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 38814 44200 38926 45000 0 FreeSans 448 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 40378 44200 40490 45000 0 FreeSans 448 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 41942 44200 42054 45000 0 FreeSans 448 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 4406 44200 4518 45000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 5970 44200 6082 45000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 7534 44200 7646 45000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 9098 44200 9210 45000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 10662 44200 10774 45000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 12226 44200 12338 45000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 13790 44200 13902 45000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 15354 44200 15466 45000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal3 s 44200 42516 45000 42756 0 FreeSans 960 0 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 42480 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 42480 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 42480 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
rlabel metal1 22494 41888 22494 41888 0 vccd1
rlabel metal1 22494 42432 22494 42432 0 vssd1
rlabel viali 33810 36754 33810 36754 0 MOS6502.ABH\[0\]
rlabel metal1 32752 41446 32752 41446 0 MOS6502.ABH\[1\]
rlabel viali 33718 37230 33718 37230 0 MOS6502.ABH\[2\]
rlabel metal1 34822 41446 34822 41446 0 MOS6502.ABH\[3\]
rlabel metal1 37168 40494 37168 40494 0 MOS6502.ABH\[4\]
rlabel via1 38024 36142 38024 36142 0 MOS6502.ABH\[5\]
rlabel metal1 43056 41446 43056 41446 0 MOS6502.ABH\[6\]
rlabel metal1 40250 40698 40250 40698 0 MOS6502.ABH\[7\]
rlabel metal2 20194 36346 20194 36346 0 MOS6502.ABL\[0\]
rlabel metal1 19090 38182 19090 38182 0 MOS6502.ABL\[1\]
rlabel metal1 19918 38828 19918 38828 0 MOS6502.ABL\[2\]
rlabel metal1 21344 41174 21344 41174 0 MOS6502.ABL\[3\]
rlabel metal1 23920 41446 23920 41446 0 MOS6502.ABL\[4\]
rlabel metal1 26588 41446 26588 41446 0 MOS6502.ABL\[5\]
rlabel metal1 27922 41242 27922 41242 0 MOS6502.ABL\[6\]
rlabel metal1 31050 41446 31050 41446 0 MOS6502.ABL\[7\]
rlabel metal1 33442 41990 33442 41990 0 MOS6502.ADD\[0\]
rlabel metal1 38686 42126 38686 42126 0 MOS6502.ADD\[1\]
rlabel metal1 34086 42126 34086 42126 0 MOS6502.ADD\[2\]
rlabel metal1 40342 41990 40342 41990 0 MOS6502.ADD\[3\]
rlabel metal1 17204 36006 17204 36006 0 MOS6502.ADD\[4\]
rlabel metal2 37582 42024 37582 42024 0 MOS6502.ADD\[5\]
rlabel metal2 17802 36890 17802 36890 0 MOS6502.ADD\[6\]
rlabel metal2 20010 36176 20010 36176 0 MOS6502.ADD\[7\]
rlabel metal1 18216 30634 18216 30634 0 MOS6502.AI\[7\]
rlabel metal2 18630 26010 18630 26010 0 MOS6502.ALU.AI7
rlabel metal2 18538 26316 18538 26316 0 MOS6502.ALU.BI7
rlabel metal1 19826 34578 19826 34578 0 MOS6502.ALU.CO
rlabel metal1 20454 26282 20454 26282 0 MOS6502.ALU.HC
rlabel metal1 21564 27438 21564 27438 0 MOS6502.ALU.temp\[0\]
rlabel metal1 14812 28186 14812 28186 0 MOS6502.ALU.temp\[1\]
rlabel metal1 13892 27846 13892 27846 0 MOS6502.ALU.temp\[2\]
rlabel metal1 13938 29818 13938 29818 0 MOS6502.ALU.temp\[3\]
rlabel metal2 12650 34578 12650 34578 0 MOS6502.ALU.temp\[4\]
rlabel metal2 16238 35972 16238 35972 0 MOS6502.ALU.temp\[5\]
rlabel metal1 16330 35802 16330 35802 0 MOS6502.ALU.temp\[6\]
rlabel metal1 18354 35666 18354 35666 0 MOS6502.ALU.temp\[7\]
rlabel metal1 17199 27030 17199 27030 0 MOS6502.ALU.temp_BI\[7\]
rlabel metal1 13386 31858 13386 31858 0 MOS6502.ALU.temp_HC
rlabel metal1 21298 16218 21298 16218 0 MOS6502.AXYS\[0\]\[0\]
rlabel metal2 21666 20196 21666 20196 0 MOS6502.AXYS\[0\]\[1\]
rlabel metal1 19964 18394 19964 18394 0 MOS6502.AXYS\[0\]\[2\]
rlabel metal1 16928 20774 16928 20774 0 MOS6502.AXYS\[0\]\[3\]
rlabel metal1 17296 22134 17296 22134 0 MOS6502.AXYS\[0\]\[4\]
rlabel metal1 18492 17306 18492 17306 0 MOS6502.AXYS\[0\]\[5\]
rlabel metal1 18630 21998 18630 21998 0 MOS6502.AXYS\[0\]\[6\]
rlabel metal1 18170 15130 18170 15130 0 MOS6502.AXYS\[0\]\[7\]
rlabel metal2 23414 16762 23414 16762 0 MOS6502.AXYS\[1\]\[0\]
rlabel metal1 22954 20910 22954 20910 0 MOS6502.AXYS\[1\]\[1\]
rlabel metal2 20562 17442 20562 17442 0 MOS6502.AXYS\[1\]\[2\]
rlabel metal1 17894 20332 17894 20332 0 MOS6502.AXYS\[1\]\[3\]
rlabel metal1 16882 25126 16882 25126 0 MOS6502.AXYS\[1\]\[4\]
rlabel metal1 17802 16218 17802 16218 0 MOS6502.AXYS\[1\]\[5\]
rlabel via1 18630 24106 18630 24106 0 MOS6502.AXYS\[1\]\[6\]
rlabel metal1 16928 15674 16928 15674 0 MOS6502.AXYS\[1\]\[7\]
rlabel metal1 23736 13498 23736 13498 0 MOS6502.AXYS\[2\]\[0\]
rlabel metal1 22954 15470 22954 15470 0 MOS6502.AXYS\[2\]\[1\]
rlabel metal2 20838 16422 20838 16422 0 MOS6502.AXYS\[2\]\[2\]
rlabel metal1 15180 19482 15180 19482 0 MOS6502.AXYS\[2\]\[3\]
rlabel metal2 14766 21760 14766 21760 0 MOS6502.AXYS\[2\]\[4\]
rlabel metal2 14674 16864 14674 16864 0 MOS6502.AXYS\[2\]\[5\]
rlabel metal1 14582 21998 14582 21998 0 MOS6502.AXYS\[2\]\[6\]
rlabel metal2 14858 16694 14858 16694 0 MOS6502.AXYS\[2\]\[7\]
rlabel metal1 21758 13192 21758 13192 0 MOS6502.AXYS\[3\]\[0\]
rlabel metal1 22586 16218 22586 16218 0 MOS6502.AXYS\[3\]\[1\]
rlabel metal1 19596 15130 19596 15130 0 MOS6502.AXYS\[3\]\[2\]
rlabel metal1 15180 20026 15180 20026 0 MOS6502.AXYS\[3\]\[3\]
rlabel metal2 14674 23902 14674 23902 0 MOS6502.AXYS\[3\]\[4\]
rlabel metal1 14904 17306 14904 17306 0 MOS6502.AXYS\[3\]\[5\]
rlabel metal1 14674 23698 14674 23698 0 MOS6502.AXYS\[3\]\[6\]
rlabel metal1 15594 14382 15594 14382 0 MOS6502.AXYS\[3\]\[7\]
rlabel metal1 27922 36754 27922 36754 0 MOS6502.C
rlabel metal1 25622 21658 25622 21658 0 MOS6502.D
rlabel viali 31602 33489 31602 33489 0 MOS6502.I
rlabel metal1 39974 11730 39974 11730 0 MOS6502.IRHOLD\[0\]
rlabel metal2 41170 11526 41170 11526 0 MOS6502.IRHOLD\[1\]
rlabel metal2 43102 11968 43102 11968 0 MOS6502.IRHOLD\[2\]
rlabel metal1 43194 13498 43194 13498 0 MOS6502.IRHOLD\[3\]
rlabel metal1 42734 16626 42734 16626 0 MOS6502.IRHOLD\[4\]
rlabel metal2 41078 13056 41078 13056 0 MOS6502.IRHOLD\[5\]
rlabel metal2 40986 15878 40986 15878 0 MOS6502.IRHOLD\[6\]
rlabel metal1 43240 17850 43240 17850 0 MOS6502.IRHOLD\[7\]
rlabel metal1 40848 12750 40848 12750 0 MOS6502.IRHOLD_valid
rlabel metal2 28106 15708 28106 15708 0 MOS6502.IR\[5\]
rlabel metal1 32936 16150 32936 16150 0 MOS6502.IR\[6\]
rlabel metal2 34178 17085 34178 17085 0 MOS6502.IR\[7\]
rlabel metal1 28474 29274 28474 29274 0 MOS6502.N
rlabel metal2 41906 33558 41906 33558 0 MOS6502.NMI_1
rlabel metal2 41078 33864 41078 33864 0 MOS6502.NMI_edge
rlabel metal1 30636 37978 30636 37978 0 MOS6502.PC\[0\]
rlabel metal1 32890 35666 32890 35666 0 MOS6502.PC\[10\]
rlabel metal1 19366 38930 19366 38930 0 MOS6502.PC\[11\]
rlabel metal2 37122 36108 37122 36108 0 MOS6502.PC\[12\]
rlabel metal2 38134 36465 38134 36465 0 MOS6502.PC\[13\]
rlabel via2 16974 38811 16974 38811 0 MOS6502.PC\[14\]
rlabel via1 39514 35666 39514 35666 0 MOS6502.PC\[15\]
rlabel metal1 21942 40154 21942 40154 0 MOS6502.PC\[1\]
rlabel metal1 22678 39270 22678 39270 0 MOS6502.PC\[2\]
rlabel metal1 22724 40358 22724 40358 0 MOS6502.PC\[3\]
rlabel metal1 33166 34000 33166 34000 0 MOS6502.PC\[4\]
rlabel metal1 28520 38726 28520 38726 0 MOS6502.PC\[5\]
rlabel metal2 26818 32538 26818 32538 0 MOS6502.PC\[6\]
rlabel metal1 29946 34986 29946 34986 0 MOS6502.PC\[7\]
rlabel metal1 33718 38352 33718 38352 0 MOS6502.PC\[8\]
rlabel metal1 37398 38726 37398 38726 0 MOS6502.PC\[9\]
rlabel metal1 26450 32878 26450 32878 0 MOS6502.V
rlabel metal1 25576 32878 25576 32878 0 MOS6502.Z
rlabel metal1 24518 21862 24518 21862 0 MOS6502.adc_bcd
rlabel metal2 28566 17544 28566 17544 0 MOS6502.adc_sbc
rlabel metal1 22916 25126 22916 25126 0 MOS6502.adj_bcd
rlabel metal1 27968 30226 27968 30226 0 MOS6502.backwards
rlabel metal1 28520 11866 28520 11866 0 MOS6502.bit_ins
rlabel metal1 30866 18054 30866 18054 0 MOS6502.clc
rlabel metal1 28244 18870 28244 18870 0 MOS6502.cld
rlabel metal1 32660 20026 32660 20026 0 MOS6502.cli
rlabel metal1 27508 14586 27508 14586 0 MOS6502.clv
rlabel metal1 27600 15062 27600 15062 0 MOS6502.compare
rlabel metal1 28658 28050 28658 28050 0 MOS6502.cond_code\[0\]
rlabel via2 26634 16235 26634 16235 0 MOS6502.cond_code\[1\]
rlabel metal1 26404 19482 26404 19482 0 MOS6502.cond_code\[2\]
rlabel metal1 32936 17646 32936 17646 0 MOS6502.dst_reg\[0\]
rlabel metal1 32706 21420 32706 21420 0 MOS6502.dst_reg\[1\]
rlabel metal1 29900 25126 29900 25126 0 MOS6502.inc
rlabel metal1 34914 20570 34914 20570 0 MOS6502.index_y
rlabel via1 34454 27965 34454 27965 0 MOS6502.load_only
rlabel metal2 31142 20162 31142 20162 0 MOS6502.load_reg
rlabel via2 24610 16779 24610 16779 0 MOS6502.op\[0\]
rlabel metal1 25668 17850 25668 17850 0 MOS6502.op\[1\]
rlabel metal2 26082 15215 26082 15215 0 MOS6502.op\[2\]
rlabel metal1 27738 17680 27738 17680 0 MOS6502.op\[3\]
rlabel metal2 33994 19057 33994 19057 0 MOS6502.php
rlabel metal1 31188 21522 31188 21522 0 MOS6502.plp
rlabel metal2 36846 34850 36846 34850 0 MOS6502.res
rlabel metal1 30038 21964 30038 21964 0 MOS6502.rotate
rlabel metal1 31188 18938 31188 18938 0 MOS6502.sec
rlabel metal2 28014 19618 28014 19618 0 MOS6502.sed
rlabel metal2 32614 19516 32614 19516 0 MOS6502.sei
rlabel metal1 28842 23698 28842 23698 0 MOS6502.shift
rlabel metal2 25254 14144 25254 14144 0 MOS6502.shift_right
rlabel metal1 31924 21998 31924 21998 0 MOS6502.src_reg\[0\]
rlabel via2 32246 11339 32246 11339 0 MOS6502.src_reg\[1\]
rlabel metal1 40296 25942 40296 25942 0 MOS6502.state\[0\]
rlabel metal1 42642 26758 42642 26758 0 MOS6502.state\[1\]
rlabel metal1 41860 23290 41860 23290 0 MOS6502.state\[2\]
rlabel metal1 40940 25398 40940 25398 0 MOS6502.state\[3\]
rlabel metal1 42918 28492 42918 28492 0 MOS6502.state\[4\]
rlabel metal1 39422 32334 39422 32334 0 MOS6502.state\[5\]
rlabel metal1 36800 21318 36800 21318 0 MOS6502.store
rlabel metal1 35282 21080 35282 21080 0 MOS6502.write_back
rlabel via1 23510 23086 23510 23086 0 _0000_
rlabel metal1 17572 34510 17572 34510 0 _0001_
rlabel metal1 30120 37230 30120 37230 0 _0002_
rlabel metal1 40240 39406 40240 39406 0 _0003_
rlabel metal2 41170 39202 41170 39202 0 _0004_
rlabel metal1 42172 38318 42172 38318 0 _0005_
rlabel metal2 41998 37026 41998 37026 0 _0006_
rlabel metal2 42642 35938 42642 35938 0 _0007_
rlabel metal1 41239 34918 41239 34918 0 _0008_
rlabel metal1 20184 40018 20184 40018 0 _0009_
rlabel metal1 21196 39406 21196 39406 0 _0010_
rlabel metal1 23460 39950 23460 39950 0 _0011_
rlabel metal2 24886 40188 24886 40188 0 _0012_
rlabel metal1 27124 38998 27124 38998 0 _0013_
rlabel metal1 28704 39610 28704 39610 0 _0014_
rlabel metal1 31520 39406 31520 39406 0 _0015_
rlabel metal2 35466 39780 35466 39780 0 _0016_
rlabel metal1 37724 38998 37724 38998 0 _0017_
rlabel metal2 40526 20196 40526 20196 0 _0018_
rlabel metal1 40526 19754 40526 19754 0 _0019_
rlabel metal2 40710 21726 40710 21726 0 _0020_
rlabel metal1 41446 22406 41446 22406 0 _0021_
rlabel metal2 42918 32028 42918 32028 0 _0022_
rlabel metal2 41630 33150 41630 33150 0 _0023_
rlabel metal2 41906 19992 41906 19992 0 _0024_
rlabel metal2 42918 20026 42918 20026 0 _0025_
rlabel metal1 42281 21590 42281 21590 0 _0026_
rlabel metal1 42090 22406 42090 22406 0 _0027_
rlabel metal1 42596 33286 42596 33286 0 _0028_
rlabel metal2 42734 33694 42734 33694 0 _0029_
rlabel metal1 22627 13226 22627 13226 0 _0030_
rlabel via1 23694 15062 23694 15062 0 _0031_
rlabel metal1 19304 14314 19304 14314 0 _0032_
rlabel metal1 13416 19414 13416 19414 0 _0033_
rlabel metal2 12558 21658 12558 21658 0 _0034_
rlabel metal1 13278 16150 13278 16150 0 _0035_
rlabel via1 13565 22610 13565 22610 0 _0036_
rlabel metal1 14025 14994 14025 14994 0 _0037_
rlabel metal1 21482 17068 21482 17068 0 _0038_
rlabel metal2 22310 21726 22310 21726 0 _0039_
rlabel metal2 20930 16966 20930 16966 0 _0040_
rlabel metal1 17608 19822 17608 19822 0 _0041_
rlabel via1 15589 25262 15589 25262 0 _0042_
rlabel via1 18542 16150 18542 16150 0 _0043_
rlabel via1 17521 24854 17521 24854 0 _0044_
rlabel metal1 15543 15470 15543 15470 0 _0045_
rlabel metal1 19269 36754 19269 36754 0 _0046_
rlabel metal2 18262 38114 18262 38114 0 _0047_
rlabel metal1 18855 38998 18855 38998 0 _0048_
rlabel metal1 20373 41514 20373 41514 0 _0049_
rlabel via1 22581 41582 22581 41582 0 _0050_
rlabel viali 25341 41582 25341 41582 0 _0051_
rlabel via1 27181 41582 27181 41582 0 _0052_
rlabel metal1 29470 41514 29470 41514 0 _0053_
rlabel metal1 28892 24854 28892 24854 0 _0054_
rlabel metal2 25530 27812 25530 27812 0 _0055_
rlabel metal1 27032 29206 27032 29206 0 _0056_
rlabel metal1 24784 20910 24784 20910 0 _0057_
rlabel metal1 29936 29614 29936 29614 0 _0058_
rlabel metal1 25238 23766 25238 23766 0 _0059_
rlabel metal1 39146 10234 39146 10234 0 _0060_
rlabel metal2 40710 10642 40710 10642 0 _0061_
rlabel metal2 42090 12002 42090 12002 0 _0062_
rlabel metal1 42136 12954 42136 12954 0 _0063_
rlabel metal2 42642 15266 42642 15266 0 _0064_
rlabel metal1 39912 13226 39912 13226 0 _0065_
rlabel metal1 41308 15130 41308 15130 0 _0066_
rlabel via1 42269 17646 42269 17646 0 _0067_
rlabel metal1 40935 18326 40935 18326 0 _0068_
rlabel via1 25433 11798 25433 11798 0 _0069_
rlabel metal1 39008 34170 39008 34170 0 _0070_
rlabel metal1 32184 17238 32184 17238 0 _0071_
rlabel metal1 30298 10710 30298 10710 0 _0072_
rlabel metal2 30590 10642 30590 10642 0 _0073_
rlabel metal1 32798 10778 32798 10778 0 _0074_
rlabel metal2 33902 20230 33902 20230 0 _0075_
rlabel metal1 34898 11050 34898 11050 0 _0076_
rlabel metal2 30130 15878 30130 15878 0 _0077_
rlabel metal2 28382 10914 28382 10914 0 _0078_
rlabel via1 29582 12818 29582 12818 0 _0079_
rlabel metal1 27508 16762 27508 16762 0 _0080_
rlabel metal1 29608 23018 29608 23018 0 _0081_
rlabel metal2 25438 21250 25438 21250 0 _0082_
rlabel metal1 27926 13974 27926 13974 0 _0083_
rlabel via1 24881 13226 24881 13226 0 _0084_
rlabel metal2 29762 21862 29762 21862 0 _0085_
rlabel metal1 26327 16490 26327 16490 0 _0086_
rlabel metal1 25116 17034 25116 17034 0 _0087_
rlabel metal1 25024 14586 25024 14586 0 _0088_
rlabel metal2 27462 18054 27462 18054 0 _0089_
rlabel metal1 27416 12614 27416 12614 0 _0090_
rlabel metal2 26818 13906 26818 13906 0 _0091_
rlabel via1 32802 18734 32802 18734 0 _0092_
rlabel metal1 31832 19482 31832 19482 0 _0093_
rlabel via1 28294 19414 28294 19414 0 _0094_
rlabel metal1 27503 18734 27503 18734 0 _0095_
rlabel metal1 29608 18666 29608 18666 0 _0096_
rlabel metal1 29900 17850 29900 17850 0 _0097_
rlabel metal1 34178 18938 34178 18938 0 _0098_
rlabel metal2 30406 20434 30406 20434 0 _0099_
rlabel metal2 38962 33762 38962 33762 0 _0100_
rlabel metal1 32568 41990 32568 41990 0 _0101_
rlabel metal1 31362 41582 31362 41582 0 _0102_
rlabel metal1 34040 40154 34040 40154 0 _0103_
rlabel metal2 35466 41786 35466 41786 0 _0104_
rlabel metal1 36524 41446 36524 41446 0 _0105_
rlabel metal1 37720 41446 37720 41446 0 _0106_
rlabel metal1 39146 41718 39146 41718 0 _0107_
rlabel metal1 41272 40494 41272 40494 0 _0108_
rlabel metal1 21781 12954 21781 12954 0 _0109_
rlabel metal1 20730 15402 20730 15402 0 _0110_
rlabel metal1 19504 13498 19504 13498 0 _0111_
rlabel metal1 14198 19754 14198 19754 0 _0112_
rlabel metal1 13468 24786 13468 24786 0 _0113_
rlabel metal2 13570 16966 13570 16966 0 _0114_
rlabel metal2 14306 25670 14306 25670 0 _0115_
rlabel metal1 14582 13498 14582 13498 0 _0116_
rlabel metal1 20184 14994 20184 14994 0 _0117_
rlabel metal1 20741 19754 20741 19754 0 _0118_
rlabel metal1 19550 16218 19550 16218 0 _0119_
rlabel via1 16141 20910 16141 20910 0 _0120_
rlabel metal2 15410 21522 15410 21522 0 _0121_
rlabel via1 17153 17170 17153 17170 0 _0122_
rlabel via1 18542 22610 18542 22610 0 _0123_
rlabel via1 17153 14994 17153 14994 0 _0124_
rlabel metal1 21298 25262 21298 25262 0 _0125_
rlabel metal1 21758 25874 21758 25874 0 _0126_
rlabel metal1 20792 24582 20792 24582 0 _0127_
rlabel metal2 22402 24174 22402 24174 0 _0128_
rlabel metal1 20654 24140 20654 24140 0 _0129_
rlabel metal2 22586 23868 22586 23868 0 _0130_
rlabel metal2 22678 19261 22678 19261 0 _0131_
rlabel metal2 23414 15878 23414 15878 0 _0132_
rlabel metal2 20746 24106 20746 24106 0 _0133_
rlabel metal1 20930 24242 20930 24242 0 _0134_
rlabel metal2 20654 24004 20654 24004 0 _0135_
rlabel metal1 21068 23698 21068 23698 0 _0136_
rlabel metal1 19918 19482 19918 19482 0 _0137_
rlabel metal2 20286 14212 20286 14212 0 _0138_
rlabel metal1 20792 23086 20792 23086 0 _0139_
rlabel metal1 20562 23188 20562 23188 0 _0140_
rlabel metal1 20930 21658 20930 21658 0 _0141_
rlabel metal2 18262 21182 18262 21182 0 _0142_
rlabel metal2 13018 20230 13018 20230 0 _0143_
rlabel metal1 13616 21998 13616 21998 0 _0144_
rlabel metal1 12880 21862 12880 21862 0 _0145_
rlabel metal1 23414 25874 23414 25874 0 _0146_
rlabel metal1 23092 26418 23092 26418 0 _0147_
rlabel metal1 24380 25330 24380 25330 0 _0148_
rlabel metal1 24564 24174 24564 24174 0 _0149_
rlabel metal1 25208 23154 25208 23154 0 _0150_
rlabel metal1 17618 16660 17618 16660 0 _0151_
rlabel metal1 12834 17204 12834 17204 0 _0152_
rlabel metal1 24012 25194 24012 25194 0 _0153_
rlabel metal2 24058 24412 24058 24412 0 _0154_
rlabel metal2 23874 24548 23874 24548 0 _0155_
rlabel metal1 24380 24786 24380 24786 0 _0156_
rlabel metal2 18170 23936 18170 23936 0 _0157_
rlabel metal2 14306 22644 14306 22644 0 _0158_
rlabel metal1 24978 25942 24978 25942 0 _0159_
rlabel metal2 24610 26044 24610 26044 0 _0160_
rlabel metal2 25714 26044 25714 26044 0 _0161_
rlabel metal1 25484 25806 25484 25806 0 _0162_
rlabel metal2 16974 16320 16974 16320 0 _0163_
rlabel metal2 15318 15266 15318 15266 0 _0164_
rlabel metal2 19458 20230 19458 20230 0 _0165_
rlabel metal1 17112 15538 17112 15538 0 _0166_
rlabel metal1 21298 17068 21298 17068 0 _0167_
rlabel metal2 22126 21556 22126 21556 0 _0168_
rlabel metal1 20884 16558 20884 16558 0 _0169_
rlabel metal1 17480 21114 17480 21114 0 _0170_
rlabel metal1 15732 24922 15732 24922 0 _0171_
rlabel metal2 18630 16116 18630 16116 0 _0172_
rlabel metal2 17710 24820 17710 24820 0 _0173_
rlabel metal2 15594 16388 15594 16388 0 _0174_
rlabel metal1 38548 31858 38548 31858 0 _0175_
rlabel metal1 38732 31994 38732 31994 0 _0176_
rlabel metal2 35374 28968 35374 28968 0 _0177_
rlabel metal2 35926 28866 35926 28866 0 _0178_
rlabel metal1 28934 28628 28934 28628 0 _0179_
rlabel metal2 35926 28356 35926 28356 0 _0180_
rlabel metal2 35190 27132 35190 27132 0 _0181_
rlabel metal1 35650 27098 35650 27098 0 _0182_
rlabel metal1 36294 28628 36294 28628 0 _0183_
rlabel metal2 37674 32368 37674 32368 0 _0184_
rlabel metal1 36156 33082 36156 33082 0 _0185_
rlabel metal1 39698 40562 39698 40562 0 _0186_
rlabel metal1 23690 41990 23690 41990 0 _0187_
rlabel metal1 19412 36346 19412 36346 0 _0188_
rlabel metal1 18676 37842 18676 37842 0 _0189_
rlabel metal2 19458 38964 19458 38964 0 _0190_
rlabel metal1 20700 42194 20700 42194 0 _0191_
rlabel metal1 22816 41242 22816 41242 0 _0192_
rlabel metal1 25392 41242 25392 41242 0 _0193_
rlabel metal1 27278 41242 27278 41242 0 _0194_
rlabel metal1 28934 41582 28934 41582 0 _0195_
rlabel metal2 30774 22406 30774 22406 0 _0196_
rlabel metal2 30406 23222 30406 23222 0 _0197_
rlabel metal1 29762 23698 29762 23698 0 _0198_
rlabel metal2 30314 23936 30314 23936 0 _0199_
rlabel metal1 29348 24038 29348 24038 0 _0200_
rlabel metal1 32614 24752 32614 24752 0 _0201_
rlabel metal2 30774 24208 30774 24208 0 _0202_
rlabel metal1 30452 24378 30452 24378 0 _0203_
rlabel metal2 32706 25840 32706 25840 0 _0204_
rlabel metal1 29440 24242 29440 24242 0 _0205_
rlabel metal1 28566 24378 28566 24378 0 _0206_
rlabel metal1 27324 26962 27324 26962 0 _0207_
rlabel metal1 26312 26486 26312 26486 0 _0208_
rlabel metal2 27094 26554 27094 26554 0 _0209_
rlabel metal1 27186 26452 27186 26452 0 _0210_
rlabel metal1 27462 25466 27462 25466 0 _0211_
rlabel metal1 26450 26554 26450 26554 0 _0212_
rlabel metal1 27232 20502 27232 20502 0 _0213_
rlabel metal1 27646 20570 27646 20570 0 _0214_
rlabel metal1 26818 26010 26818 26010 0 _0215_
rlabel metal2 25714 27268 25714 27268 0 _0216_
rlabel metal1 28014 28186 28014 28186 0 _0217_
rlabel metal1 27876 26758 27876 26758 0 _0218_
rlabel metal2 27370 27812 27370 27812 0 _0219_
rlabel metal1 26818 28186 26818 28186 0 _0220_
rlabel metal1 28244 20774 28244 20774 0 _0221_
rlabel metal1 27692 21114 27692 21114 0 _0222_
rlabel metal1 26496 21658 26496 21658 0 _0223_
rlabel metal1 35466 19924 35466 19924 0 _0224_
rlabel metal1 28290 20570 28290 20570 0 _0225_
rlabel metal2 28198 21250 28198 21250 0 _0226_
rlabel metal1 25116 21522 25116 21522 0 _0227_
rlabel metal2 31510 25636 31510 25636 0 _0228_
rlabel metal2 31050 26112 31050 26112 0 _0229_
rlabel metal2 30590 27472 30590 27472 0 _0230_
rlabel metal2 32338 25092 32338 25092 0 _0231_
rlabel metal1 31004 25466 31004 25466 0 _0232_
rlabel metal1 30222 28730 30222 28730 0 _0233_
rlabel metal2 30038 29750 30038 29750 0 _0234_
rlabel metal1 26910 24208 26910 24208 0 _0235_
rlabel metal1 19136 25806 19136 25806 0 _0236_
rlabel metal2 19826 26588 19826 26588 0 _0237_
rlabel metal1 21666 24310 21666 24310 0 _0238_
rlabel metal2 27370 23562 27370 23562 0 _0239_
rlabel metal1 26818 22950 26818 22950 0 _0240_
rlabel metal1 26910 23154 26910 23154 0 _0241_
rlabel metal2 25990 23494 25990 23494 0 _0242_
rlabel metal2 41170 18122 41170 18122 0 _0243_
rlabel metal1 42918 11118 42918 11118 0 _0244_
rlabel metal2 39422 10506 39422 10506 0 _0245_
rlabel metal2 40894 10234 40894 10234 0 _0246_
rlabel metal2 42366 11526 42366 11526 0 _0247_
rlabel metal1 42274 12818 42274 12818 0 _0248_
rlabel metal2 42826 15708 42826 15708 0 _0249_
rlabel metal1 39330 13328 39330 13328 0 _0250_
rlabel metal1 41584 14994 41584 14994 0 _0251_
rlabel metal2 42642 18564 42642 18564 0 _0252_
rlabel metal2 40158 18292 40158 18292 0 _0253_
rlabel metal1 40480 18938 40480 18938 0 _0254_
rlabel metal2 35006 11798 35006 11798 0 _0255_
rlabel metal2 31786 13464 31786 13464 0 _0256_
rlabel metal2 32798 11900 32798 11900 0 _0257_
rlabel metal1 34822 12886 34822 12886 0 _0258_
rlabel metal1 33534 12954 33534 12954 0 _0259_
rlabel metal1 32430 11866 32430 11866 0 _0260_
rlabel metal2 31602 14144 31602 14144 0 _0261_
rlabel metal2 34546 14756 34546 14756 0 _0262_
rlabel metal2 34178 13770 34178 13770 0 _0263_
rlabel metal2 32292 12716 32292 12716 0 _0264_
rlabel metal2 32522 13260 32522 13260 0 _0265_
rlabel metal1 32752 12750 32752 12750 0 _0266_
rlabel metal1 34500 12274 34500 12274 0 _0267_
rlabel metal1 28842 15130 28842 15130 0 _0268_
rlabel metal1 34316 12614 34316 12614 0 _0269_
rlabel metal1 33166 12138 33166 12138 0 _0270_
rlabel metal2 32062 11934 32062 11934 0 _0271_
rlabel metal1 32706 10608 32706 10608 0 _0272_
rlabel metal2 25622 11764 25622 11764 0 _0273_
rlabel metal1 40020 16762 40020 16762 0 _0274_
rlabel metal1 31464 13362 31464 13362 0 _0275_
rlabel metal2 32982 13056 32982 13056 0 _0276_
rlabel metal1 32246 12614 32246 12614 0 _0277_
rlabel metal1 31832 13498 31832 13498 0 _0278_
rlabel metal2 32154 17340 32154 17340 0 _0279_
rlabel metal1 34868 11322 34868 11322 0 _0280_
rlabel metal1 30268 12342 30268 12342 0 _0281_
rlabel metal1 31050 12614 31050 12614 0 _0282_
rlabel metal2 30866 11968 30866 11968 0 _0283_
rlabel metal1 29762 10608 29762 10608 0 _0284_
rlabel metal2 32798 15708 32798 15708 0 _0285_
rlabel metal1 32706 15572 32706 15572 0 _0286_
rlabel metal2 31878 13124 31878 13124 0 _0287_
rlabel metal2 30774 11594 30774 11594 0 _0288_
rlabel metal1 34316 11798 34316 11798 0 _0289_
rlabel metal2 34776 11730 34776 11730 0 _0290_
rlabel metal1 32798 10540 32798 10540 0 _0291_
rlabel metal1 35006 14960 35006 14960 0 _0292_
rlabel via1 34717 15062 34717 15062 0 _0293_
rlabel metal1 35328 15130 35328 15130 0 _0294_
rlabel metal1 34500 19822 34500 19822 0 _0295_
rlabel metal1 35190 10778 35190 10778 0 _0296_
rlabel metal1 34316 10778 34316 10778 0 _0297_
rlabel metal1 31004 15538 31004 15538 0 _0298_
rlabel metal1 28796 10642 28796 10642 0 _0299_
rlabel metal2 29394 19584 29394 19584 0 _0300_
rlabel metal1 29486 13498 29486 13498 0 _0301_
rlabel metal2 35328 23460 35328 23460 0 _0302_
rlabel metal1 28842 16966 28842 16966 0 _0303_
rlabel metal1 30176 21930 30176 21930 0 _0304_
rlabel metal1 28198 17850 28198 17850 0 _0305_
rlabel metal1 28750 14960 28750 14960 0 _0306_
rlabel metal1 28336 14994 28336 14994 0 _0307_
rlabel metal1 25346 14008 25346 14008 0 _0308_
rlabel metal1 24564 13906 24564 13906 0 _0309_
rlabel metal2 27646 16388 27646 16388 0 _0310_
rlabel metal2 29210 14790 29210 14790 0 _0311_
rlabel metal2 30130 14212 30130 14212 0 _0312_
rlabel metal2 29762 14688 29762 14688 0 _0313_
rlabel metal2 28750 14433 28750 14433 0 _0314_
rlabel metal2 31510 14620 31510 14620 0 _0315_
rlabel metal1 25760 15538 25760 15538 0 _0316_
rlabel metal1 28612 18666 28612 18666 0 _0317_
rlabel metal2 25254 14858 25254 14858 0 _0318_
rlabel metal1 28198 16762 28198 16762 0 _0319_
rlabel metal2 39974 17391 39974 17391 0 _0320_
rlabel metal1 27278 12818 27278 12818 0 _0321_
rlabel metal1 26772 13362 26772 13362 0 _0322_
rlabel metal1 32476 20434 32476 20434 0 _0323_
rlabel metal2 32338 19414 32338 19414 0 _0324_
rlabel metal2 30406 17204 30406 17204 0 _0325_
rlabel metal1 40158 33320 40158 33320 0 _0326_
rlabel metal1 32292 40698 32292 40698 0 _0327_
rlabel metal2 30682 41718 30682 41718 0 _0328_
rlabel metal1 34270 40052 34270 40052 0 _0329_
rlabel metal1 34868 42194 34868 42194 0 _0330_
rlabel metal2 36938 41140 36938 41140 0 _0331_
rlabel metal1 37444 40698 37444 40698 0 _0332_
rlabel metal1 38640 40698 38640 40698 0 _0333_
rlabel metal1 40986 41446 40986 41446 0 _0334_
rlabel metal2 20470 20706 20470 20706 0 _0335_
rlabel metal1 15042 20366 15042 20366 0 _0336_
rlabel metal2 21298 12988 21298 12988 0 _0337_
rlabel metal1 21114 15470 21114 15470 0 _0338_
rlabel metal1 19550 13294 19550 13294 0 _0339_
rlabel metal1 13984 20434 13984 20434 0 _0340_
rlabel metal1 13616 24378 13616 24378 0 _0341_
rlabel metal1 14030 16558 14030 16558 0 _0342_
rlabel metal1 14306 23834 14306 23834 0 _0343_
rlabel metal2 14858 13770 14858 13770 0 _0344_
rlabel metal1 18446 21522 18446 21522 0 _0345_
rlabel metal2 17710 15538 17710 15538 0 _0346_
rlabel metal1 19550 15504 19550 15504 0 _0347_
rlabel metal1 21206 18938 21206 18938 0 _0348_
rlabel metal1 19412 16082 19412 16082 0 _0349_
rlabel metal1 16284 20026 16284 20026 0 _0350_
rlabel metal1 15410 22406 15410 22406 0 _0351_
rlabel metal1 17112 16422 17112 16422 0 _0352_
rlabel metal2 18630 22610 18630 22610 0 _0353_
rlabel metal1 17020 14586 17020 14586 0 _0354_
rlabel metal1 35374 33422 35374 33422 0 _0355_
rlabel metal2 39238 15521 39238 15521 0 _0356_
rlabel metal1 39514 14348 39514 14348 0 _0357_
rlabel metal1 40302 17170 40302 17170 0 _0358_
rlabel metal1 39744 16014 39744 16014 0 _0359_
rlabel metal2 38778 13124 38778 13124 0 _0360_
rlabel metal1 38226 13940 38226 13940 0 _0361_
rlabel metal1 40434 13906 40434 13906 0 _0362_
rlabel via1 39790 14450 39790 14450 0 _0363_
rlabel metal2 41998 30906 41998 30906 0 _0364_
rlabel metal1 38824 26894 38824 26894 0 _0365_
rlabel metal1 40434 27472 40434 27472 0 _0366_
rlabel metal1 37812 29070 37812 29070 0 _0367_
rlabel metal1 41032 24786 41032 24786 0 _0368_
rlabel metal1 41285 29070 41285 29070 0 _0369_
rlabel metal1 37444 29138 37444 29138 0 _0370_
rlabel metal1 35098 31280 35098 31280 0 _0371_
rlabel via2 34546 30243 34546 30243 0 _0372_
rlabel metal1 38226 28628 38226 28628 0 _0373_
rlabel metal1 42596 27438 42596 27438 0 _0374_
rlabel metal2 41354 25772 41354 25772 0 _0375_
rlabel metal2 38410 29308 38410 29308 0 _0376_
rlabel metal1 32338 30294 32338 30294 0 _0377_
rlabel metal1 36754 25806 36754 25806 0 _0378_
rlabel metal2 41354 29682 41354 29682 0 _0379_
rlabel metal2 40158 34782 40158 34782 0 _0380_
rlabel metal1 32568 31994 32568 31994 0 _0381_
rlabel metal1 42366 30226 42366 30226 0 _0382_
rlabel metal2 35742 31297 35742 31297 0 _0383_
rlabel metal1 41630 23290 41630 23290 0 _0384_
rlabel metal1 34730 23698 34730 23698 0 _0385_
rlabel metal1 33396 27506 33396 27506 0 _0386_
rlabel metal2 32522 28628 32522 28628 0 _0387_
rlabel metal2 40526 26826 40526 26826 0 _0388_
rlabel metal1 34500 27574 34500 27574 0 _0389_
rlabel metal1 32522 31790 32522 31790 0 _0390_
rlabel metal1 31809 31994 31809 31994 0 _0391_
rlabel metal2 39054 29784 39054 29784 0 _0392_
rlabel metal1 37812 26282 37812 26282 0 _0393_
rlabel metal1 32982 26384 32982 26384 0 _0394_
rlabel metal1 38870 39814 38870 39814 0 _0395_
rlabel metal2 28842 33490 28842 33490 0 _0396_
rlabel metal1 21114 34510 21114 34510 0 _0397_
rlabel via1 35653 27438 35653 27438 0 _0398_
rlabel metal1 42826 22746 42826 22746 0 _0399_
rlabel metal2 40710 24276 40710 24276 0 _0400_
rlabel metal2 35558 28288 35558 28288 0 _0401_
rlabel metal1 39698 30226 39698 30226 0 _0402_
rlabel metal1 34822 30294 34822 30294 0 _0403_
rlabel metal1 37766 32470 37766 32470 0 _0404_
rlabel metal1 40066 30226 40066 30226 0 _0405_
rlabel metal1 37766 30702 37766 30702 0 _0406_
rlabel metal1 41170 30192 41170 30192 0 _0407_
rlabel metal1 36846 29274 36846 29274 0 _0408_
rlabel metal1 36800 24174 36800 24174 0 _0409_
rlabel metal1 41262 20808 41262 20808 0 _0410_
rlabel metal1 39422 29172 39422 29172 0 _0411_
rlabel metal1 37260 29750 37260 29750 0 _0412_
rlabel metal1 37076 33966 37076 33966 0 _0413_
rlabel metal3 40756 31756 40756 31756 0 _0414_
rlabel metal1 31878 29512 31878 29512 0 _0415_
rlabel metal1 35236 25262 35236 25262 0 _0416_
rlabel metal1 34224 24582 34224 24582 0 _0417_
rlabel metal2 31418 27268 31418 27268 0 _0418_
rlabel metal2 33718 35360 33718 35360 0 _0419_
rlabel metal2 31234 29410 31234 29410 0 _0420_
rlabel metal1 29785 27030 29785 27030 0 _0421_
rlabel metal1 40940 28390 40940 28390 0 _0422_
rlabel metal1 28290 30668 28290 30668 0 _0423_
rlabel metal1 15916 32334 15916 32334 0 _0424_
rlabel metal1 24840 27098 24840 27098 0 _0425_
rlabel metal1 19274 27438 19274 27438 0 _0426_
rlabel metal2 15226 31994 15226 31994 0 _0427_
rlabel metal2 40986 30192 40986 30192 0 _0428_
rlabel metal2 33994 29308 33994 29308 0 _0429_
rlabel metal1 36800 30634 36800 30634 0 _0430_
rlabel metal2 36386 27132 36386 27132 0 _0431_
rlabel metal2 39192 25262 39192 25262 0 _0432_
rlabel metal2 43102 25483 43102 25483 0 _0433_
rlabel metal1 38732 26350 38732 26350 0 _0434_
rlabel metal1 37858 25194 37858 25194 0 _0435_
rlabel metal2 36478 25670 36478 25670 0 _0436_
rlabel metal1 36662 26316 36662 26316 0 _0437_
rlabel metal1 40710 32810 40710 32810 0 _0438_
rlabel metal1 36432 20366 36432 20366 0 _0439_
rlabel metal1 36110 28594 36110 28594 0 _0440_
rlabel metal2 31234 28220 31234 28220 0 _0441_
rlabel metal1 31050 27846 31050 27846 0 _0442_
rlabel metal1 37352 27574 37352 27574 0 _0443_
rlabel metal2 37766 25160 37766 25160 0 _0444_
rlabel metal1 32292 23630 32292 23630 0 _0445_
rlabel metal1 32614 27438 32614 27438 0 _0446_
rlabel metal2 32982 28356 32982 28356 0 _0447_
rlabel metal1 32614 28628 32614 28628 0 _0448_
rlabel metal1 17342 31858 17342 31858 0 _0449_
rlabel metal1 15226 31994 15226 31994 0 _0450_
rlabel metal1 16008 29682 16008 29682 0 _0451_
rlabel metal1 15962 29104 15962 29104 0 _0452_
rlabel metal1 15042 31824 15042 31824 0 _0453_
rlabel metal1 13846 33320 13846 33320 0 _0454_
rlabel metal2 20378 29036 20378 29036 0 _0455_
rlabel metal2 18262 34510 18262 34510 0 _0456_
rlabel metal2 41722 27200 41722 27200 0 _0457_
rlabel metal2 42918 24038 42918 24038 0 _0458_
rlabel metal1 42826 25670 42826 25670 0 _0459_
rlabel metal2 42826 24718 42826 24718 0 _0460_
rlabel metal1 36018 32368 36018 32368 0 _0461_
rlabel metal1 25162 30158 25162 30158 0 _0462_
rlabel metal1 22862 30192 22862 30192 0 _0463_
rlabel metal1 20378 32300 20378 32300 0 _0464_
rlabel metal2 34270 31926 34270 31926 0 _0465_
rlabel metal1 27232 32878 27232 32878 0 _0466_
rlabel metal2 36294 27982 36294 27982 0 _0467_
rlabel metal1 34638 30634 34638 30634 0 _0468_
rlabel metal2 32338 30906 32338 30906 0 _0469_
rlabel metal1 28842 31280 28842 31280 0 _0470_
rlabel metal1 30774 28016 30774 28016 0 _0471_
rlabel metal1 32384 27370 32384 27370 0 _0472_
rlabel metal1 34178 29172 34178 29172 0 _0473_
rlabel metal2 40986 32776 40986 32776 0 _0474_
rlabel metal2 32338 27676 32338 27676 0 _0475_
rlabel metal1 33902 21522 33902 21522 0 _0476_
rlabel metal2 40342 24735 40342 24735 0 _0477_
rlabel metal2 39514 24140 39514 24140 0 _0478_
rlabel metal1 33166 21386 33166 21386 0 _0479_
rlabel metal1 32338 27098 32338 27098 0 _0480_
rlabel metal2 31694 28322 31694 28322 0 _0481_
rlabel metal1 23874 32946 23874 32946 0 _0482_
rlabel metal2 34362 24038 34362 24038 0 _0483_
rlabel metal2 32982 21454 32982 21454 0 _0484_
rlabel metal2 34638 26044 34638 26044 0 _0485_
rlabel metal1 34684 25942 34684 25942 0 _0486_
rlabel metal1 38778 22032 38778 22032 0 _0487_
rlabel metal2 34086 26095 34086 26095 0 _0488_
rlabel metal1 33074 22746 33074 22746 0 _0489_
rlabel metal1 21114 17816 21114 17816 0 _0490_
rlabel metal2 33074 21114 33074 21114 0 _0491_
rlabel metal1 21114 20978 21114 20978 0 _0492_
rlabel metal1 20516 20502 20516 20502 0 _0493_
rlabel metal2 32890 21964 32890 21964 0 _0494_
rlabel metal1 23506 20468 23506 20468 0 _0495_
rlabel metal1 19274 20298 19274 20298 0 _0496_
rlabel metal1 18032 20366 18032 20366 0 _0497_
rlabel metal2 22954 17918 22954 17918 0 _0498_
rlabel metal1 15594 19380 15594 19380 0 _0499_
rlabel metal1 18170 18802 18170 18802 0 _0500_
rlabel metal1 15640 17306 15640 17306 0 _0501_
rlabel metal1 16146 18224 16146 18224 0 _0502_
rlabel metal2 17894 18751 17894 18751 0 _0503_
rlabel metal1 30176 32266 30176 32266 0 _0504_
rlabel metal1 29624 32878 29624 32878 0 _0505_
rlabel metal1 21620 32810 21620 32810 0 _0506_
rlabel metal2 20194 33014 20194 33014 0 _0507_
rlabel metal1 21298 30260 21298 30260 0 _0508_
rlabel metal1 20516 32878 20516 32878 0 _0509_
rlabel metal1 20976 31790 20976 31790 0 _0510_
rlabel metal1 20562 31858 20562 31858 0 _0511_
rlabel metal2 20470 33388 20470 33388 0 _0512_
rlabel metal1 20102 33082 20102 33082 0 _0513_
rlabel metal1 15134 23120 15134 23120 0 _0514_
rlabel metal1 16744 23290 16744 23290 0 _0515_
rlabel metal2 34362 32810 34362 32810 0 _0516_
rlabel metal1 28934 32368 28934 32368 0 _0517_
rlabel metal2 28750 31994 28750 31994 0 _0518_
rlabel metal2 19642 33184 19642 33184 0 _0519_
rlabel metal1 20884 33422 20884 33422 0 _0520_
rlabel metal1 14122 33422 14122 33422 0 _0521_
rlabel metal1 13478 33898 13478 33898 0 _0522_
rlabel metal1 15272 21658 15272 21658 0 _0523_
rlabel metal2 16330 23290 16330 23290 0 _0524_
rlabel metal1 18676 34918 18676 34918 0 _0525_
rlabel metal2 37950 33609 37950 33609 0 _0526_
rlabel metal2 23598 33303 23598 33303 0 _0527_
rlabel metal1 23000 33490 23000 33490 0 _0528_
rlabel metal1 20516 32402 20516 32402 0 _0529_
rlabel metal1 22310 32878 22310 32878 0 _0530_
rlabel metal2 22678 33116 22678 33116 0 _0531_
rlabel metal1 22540 32538 22540 32538 0 _0532_
rlabel metal1 21942 32742 21942 32742 0 _0533_
rlabel metal2 13938 32640 13938 32640 0 _0534_
rlabel metal2 15410 32334 15410 32334 0 _0535_
rlabel metal2 14122 32572 14122 32572 0 _0536_
rlabel metal1 13708 32470 13708 32470 0 _0537_
rlabel metal2 15318 19788 15318 19788 0 _0538_
rlabel metal2 15962 19958 15962 19958 0 _0539_
rlabel metal1 17204 20570 17204 20570 0 _0540_
rlabel metal1 34914 32300 34914 32300 0 _0541_
rlabel metal1 30774 32198 30774 32198 0 _0542_
rlabel metal1 21482 31348 21482 31348 0 _0543_
rlabel metal1 23092 30702 23092 30702 0 _0544_
rlabel metal1 18814 30668 18814 30668 0 _0545_
rlabel metal1 22724 30838 22724 30838 0 _0546_
rlabel metal1 21574 31790 21574 31790 0 _0547_
rlabel metal2 21666 30906 21666 30906 0 _0548_
rlabel metal2 21942 31076 21942 31076 0 _0549_
rlabel metal1 21850 31824 21850 31824 0 _0550_
rlabel metal2 22310 31484 22310 31484 0 _0551_
rlabel metal1 13386 31212 13386 31212 0 _0552_
rlabel metal1 12282 31348 12282 31348 0 _0553_
rlabel metal1 12604 31450 12604 31450 0 _0554_
rlabel metal1 13570 31314 13570 31314 0 _0555_
rlabel metal1 12098 30260 12098 30260 0 _0556_
rlabel metal2 20470 30498 20470 30498 0 _0557_
rlabel metal2 17894 29818 17894 29818 0 _0558_
rlabel metal1 22540 17578 22540 17578 0 _0559_
rlabel metal1 23046 19346 23046 19346 0 _0560_
rlabel metal2 23598 18870 23598 18870 0 _0561_
rlabel metal2 23690 19584 23690 19584 0 _0562_
rlabel metal2 24334 34544 24334 34544 0 _0563_
rlabel metal2 31786 33286 31786 33286 0 _0564_
rlabel metal1 23782 32878 23782 32878 0 _0565_
rlabel metal2 18354 33524 18354 33524 0 _0566_
rlabel metal1 19826 30294 19826 30294 0 _0567_
rlabel via1 19568 30226 19568 30226 0 _0568_
rlabel metal2 18170 29818 18170 29818 0 _0569_
rlabel metal1 22724 28458 22724 28458 0 _0570_
rlabel metal2 22494 20026 22494 20026 0 _0571_
rlabel metal1 22494 18394 22494 18394 0 _0572_
rlabel metal1 22172 20026 22172 20026 0 _0573_
rlabel metal2 29946 30906 29946 30906 0 _0574_
rlabel metal1 21850 28560 21850 28560 0 _0575_
rlabel metal1 20930 28628 20930 28628 0 _0576_
rlabel metal2 19366 29138 19366 29138 0 _0577_
rlabel metal2 18446 28798 18446 28798 0 _0578_
rlabel metal1 29716 26554 29716 26554 0 _0579_
rlabel metal1 30038 25296 30038 25296 0 _0580_
rlabel metal2 29210 27268 29210 27268 0 _0581_
rlabel metal2 29394 27846 29394 27846 0 _0582_
rlabel metal2 30406 27200 30406 27200 0 _0583_
rlabel metal1 30360 25466 30360 25466 0 _0584_
rlabel metal1 35420 23698 35420 23698 0 _0585_
rlabel metal1 34822 23766 34822 23766 0 _0586_
rlabel metal1 34822 31926 34822 31926 0 _0587_
rlabel metal1 33442 30906 33442 30906 0 _0588_
rlabel metal2 32844 30124 32844 30124 0 _0589_
rlabel metal2 30222 29104 30222 29104 0 _0590_
rlabel metal2 29578 27846 29578 27846 0 _0591_
rlabel metal1 17618 28084 17618 28084 0 _0592_
rlabel metal1 17434 28594 17434 28594 0 _0593_
rlabel metal1 17894 28594 17894 28594 0 _0594_
rlabel metal2 15226 28220 15226 28220 0 _0595_
rlabel metal2 16422 29376 16422 29376 0 _0596_
rlabel metal1 20240 28526 20240 28526 0 _0597_
rlabel metal2 15870 29308 15870 29308 0 _0598_
rlabel metal1 19274 29274 19274 29274 0 _0599_
rlabel metal1 20562 27982 20562 27982 0 _0600_
rlabel metal2 20102 29444 20102 29444 0 _0601_
rlabel metal1 20240 28730 20240 28730 0 _0602_
rlabel metal2 16146 29342 16146 29342 0 _0603_
rlabel metal2 20930 17629 20930 17629 0 _0604_
rlabel metal2 21206 18734 21206 18734 0 _0605_
rlabel metal1 20332 17714 20332 17714 0 _0606_
rlabel metal1 20056 17850 20056 17850 0 _0607_
rlabel via2 22770 19499 22770 19499 0 _0608_
rlabel metal2 32430 31790 32430 31790 0 _0609_
rlabel metal2 24978 31450 24978 31450 0 _0610_
rlabel metal2 22034 29852 22034 29852 0 _0611_
rlabel metal1 16560 29138 16560 29138 0 _0612_
rlabel metal1 15410 29138 15410 29138 0 _0613_
rlabel metal1 15502 28730 15502 28730 0 _0614_
rlabel metal1 13156 29614 13156 29614 0 _0615_
rlabel metal1 16146 30804 16146 30804 0 _0616_
rlabel metal2 21206 29818 21206 29818 0 _0617_
rlabel metal1 23644 29682 23644 29682 0 _0618_
rlabel metal1 22218 29546 22218 29546 0 _0619_
rlabel metal1 21804 29614 21804 29614 0 _0620_
rlabel metal1 22540 29274 22540 29274 0 _0621_
rlabel metal1 12190 29716 12190 29716 0 _0622_
rlabel metal2 13938 29886 13938 29886 0 _0623_
rlabel metal1 13938 29274 13938 29274 0 _0624_
rlabel metal1 14490 29580 14490 29580 0 _0625_
rlabel metal2 13018 29546 13018 29546 0 _0626_
rlabel metal1 12834 29818 12834 29818 0 _0627_
rlabel metal2 13294 32368 13294 32368 0 _0628_
rlabel metal2 15134 28186 15134 28186 0 _0629_
rlabel metal1 13294 28934 13294 28934 0 _0630_
rlabel metal1 16284 34986 16284 34986 0 _0631_
rlabel metal1 12512 31790 12512 31790 0 _0632_
rlabel metal1 13524 32402 13524 32402 0 _0633_
rlabel metal1 13202 32198 13202 32198 0 _0634_
rlabel metal2 13294 34034 13294 34034 0 _0635_
rlabel metal2 13570 33796 13570 33796 0 _0636_
rlabel metal2 14490 34374 14490 34374 0 _0637_
rlabel metal2 15502 17850 15502 17850 0 _0638_
rlabel metal1 16606 17612 16606 17612 0 _0639_
rlabel via2 17250 17629 17250 17629 0 _0640_
rlabel metal1 28934 30294 28934 30294 0 _0641_
rlabel metal1 37398 34374 37398 34374 0 _0642_
rlabel metal1 28336 31246 28336 31246 0 _0643_
rlabel metal2 18722 32606 18722 32606 0 _0644_
rlabel metal2 20010 32300 20010 32300 0 _0645_
rlabel metal1 19274 31926 19274 31926 0 _0646_
rlabel metal2 19182 32844 19182 32844 0 _0647_
rlabel metal1 18400 32470 18400 32470 0 _0648_
rlabel metal2 16514 32674 16514 32674 0 _0649_
rlabel metal2 16422 33388 16422 33388 0 _0650_
rlabel metal2 15778 33660 15778 33660 0 _0651_
rlabel metal1 16100 33626 16100 33626 0 _0652_
rlabel metal1 15180 34578 15180 34578 0 _0653_
rlabel metal1 15870 34544 15870 34544 0 _0654_
rlabel metal1 15318 34986 15318 34986 0 _0655_
rlabel metal2 15502 35462 15502 35462 0 _0656_
rlabel metal1 18676 31858 18676 31858 0 _0657_
rlabel metal2 18722 31076 18722 31076 0 _0658_
rlabel metal1 20194 31314 20194 31314 0 _0659_
rlabel metal1 19044 31110 19044 31110 0 _0660_
rlabel metal1 17572 33422 17572 33422 0 _0661_
rlabel metal1 17388 32878 17388 32878 0 _0662_
rlabel metal2 18078 34510 18078 34510 0 _0663_
rlabel metal1 17664 33490 17664 33490 0 _0664_
rlabel metal1 16790 33898 16790 33898 0 _0665_
rlabel metal2 17986 34510 17986 34510 0 _0666_
rlabel via1 16882 35054 16882 35054 0 _0667_
rlabel metal1 17572 35666 17572 35666 0 _0668_
rlabel metal1 17572 34170 17572 34170 0 _0669_
rlabel metal2 17434 34748 17434 34748 0 _0670_
rlabel metal1 13800 34170 13800 34170 0 _0671_
rlabel metal2 14030 35190 14030 35190 0 _0672_
rlabel metal2 17158 34748 17158 34748 0 _0673_
rlabel metal1 24794 22746 24794 22746 0 _0674_
rlabel metal2 18262 28220 18262 28220 0 _0675_
rlabel metal1 17848 27982 17848 27982 0 _0676_
rlabel metal1 38318 41446 38318 41446 0 _0677_
rlabel metal1 38824 41990 38824 41990 0 _0678_
rlabel metal1 39698 32810 39698 32810 0 _0679_
rlabel metal1 39882 31790 39882 31790 0 _0680_
rlabel metal1 40342 32436 40342 32436 0 _0681_
rlabel metal2 40710 32266 40710 32266 0 _0682_
rlabel metal1 40181 35666 40181 35666 0 _0683_
rlabel via2 35926 36125 35926 36125 0 _0684_
rlabel metal2 35006 35836 35006 35836 0 _0685_
rlabel metal1 31004 36142 31004 36142 0 _0686_
rlabel metal1 30360 36074 30360 36074 0 _0687_
rlabel metal1 39054 28424 39054 28424 0 _0688_
rlabel metal1 40204 15878 40204 15878 0 _0689_
rlabel metal1 35834 34986 35834 34986 0 _0690_
rlabel metal2 30498 37366 30498 37366 0 _0691_
rlabel metal1 29670 37774 29670 37774 0 _0692_
rlabel metal1 37950 32436 37950 32436 0 _0693_
rlabel metal1 40250 29716 40250 29716 0 _0694_
rlabel metal1 37076 31858 37076 31858 0 _0695_
rlabel metal1 36846 31348 36846 31348 0 _0696_
rlabel metal2 36754 30328 36754 30328 0 _0697_
rlabel metal1 36846 31994 36846 31994 0 _0698_
rlabel metal2 37490 32623 37490 32623 0 _0699_
rlabel metal2 29762 39032 29762 39032 0 _0700_
rlabel metal1 34408 33014 34408 33014 0 _0701_
rlabel via2 34914 35173 34914 35173 0 _0702_
rlabel metal2 20838 39270 20838 39270 0 _0703_
rlabel metal1 20378 39610 20378 39610 0 _0704_
rlabel metal1 20194 39066 20194 39066 0 _0705_
rlabel metal2 38318 34306 38318 34306 0 _0706_
rlabel metal2 36478 34527 36478 34527 0 _0707_
rlabel metal2 26082 36754 26082 36754 0 _0708_
rlabel metal1 25024 37162 25024 37162 0 _0709_
rlabel metal1 22954 40086 22954 40086 0 _0710_
rlabel metal1 30866 39984 30866 39984 0 _0711_
rlabel metal1 24518 38522 24518 38522 0 _0712_
rlabel metal1 24334 38794 24334 38794 0 _0713_
rlabel metal2 25070 39610 25070 39610 0 _0714_
rlabel metal1 25208 37706 25208 37706 0 _0715_
rlabel metal1 24748 39406 24748 39406 0 _0716_
rlabel metal1 25852 39406 25852 39406 0 _0717_
rlabel metal2 26358 38046 26358 38046 0 _0718_
rlabel metal1 26910 39338 26910 39338 0 _0719_
rlabel metal1 28612 39406 28612 39406 0 _0720_
rlabel metal2 28658 38726 28658 38726 0 _0721_
rlabel metal2 28382 39134 28382 39134 0 _0722_
rlabel metal2 30682 39678 30682 39678 0 _0723_
rlabel metal1 32522 37230 32522 37230 0 _0724_
rlabel metal1 31832 37094 31832 37094 0 _0725_
rlabel metal2 30866 39372 30866 39372 0 _0726_
rlabel metal2 31786 39542 31786 39542 0 _0727_
rlabel metal2 31050 39542 31050 39542 0 _0728_
rlabel metal2 35650 30532 35650 30532 0 _0729_
rlabel metal1 35604 35666 35604 35666 0 _0730_
rlabel metal1 35558 36822 35558 36822 0 _0731_
rlabel metal1 33902 37264 33902 37264 0 _0732_
rlabel metal1 34684 36754 34684 36754 0 _0733_
rlabel metal1 35512 36890 35512 36890 0 _0734_
rlabel metal1 35052 37842 35052 37842 0 _0735_
rlabel via1 36118 39270 36118 39270 0 _0736_
rlabel metal1 36524 38930 36524 38930 0 _0737_
rlabel metal2 36938 39236 36938 39236 0 _0738_
rlabel metal2 34270 37145 34270 37145 0 _0739_
rlabel metal1 40158 38726 40158 38726 0 _0740_
rlabel metal1 39422 37230 39422 37230 0 _0741_
rlabel metal1 40526 38250 40526 38250 0 _0742_
rlabel metal1 41262 38896 41262 38896 0 _0743_
rlabel metal2 41078 38726 41078 38726 0 _0744_
rlabel metal1 40066 36176 40066 36176 0 _0745_
rlabel metal2 41170 36788 41170 36788 0 _0746_
rlabel metal1 39330 36278 39330 36278 0 _0747_
rlabel metal2 40802 37026 40802 37026 0 _0748_
rlabel metal1 41492 36754 41492 36754 0 _0749_
rlabel metal1 42090 36788 42090 36788 0 _0750_
rlabel metal1 39146 35258 39146 35258 0 _0751_
rlabel metal1 41216 36142 41216 36142 0 _0752_
rlabel metal2 41354 36074 41354 36074 0 _0753_
rlabel metal2 41814 35836 41814 35836 0 _0754_
rlabel metal1 42412 35666 42412 35666 0 _0755_
rlabel metal1 38778 35666 38778 35666 0 _0756_
rlabel metal2 40618 35292 40618 35292 0 _0757_
rlabel metal1 12880 31994 12880 31994 0 _0758_
rlabel metal1 12466 30158 12466 30158 0 _0759_
rlabel metal2 13570 29818 13570 29818 0 _0760_
rlabel metal2 35926 23052 35926 23052 0 _0761_
rlabel metal1 37076 22406 37076 22406 0 _0762_
rlabel metal1 40802 14994 40802 14994 0 _0763_
rlabel metal1 34730 12614 34730 12614 0 _0764_
rlabel metal1 38134 11152 38134 11152 0 _0765_
rlabel metal1 37996 10710 37996 10710 0 _0766_
rlabel metal2 37306 14076 37306 14076 0 _0767_
rlabel metal2 39422 12036 39422 12036 0 _0768_
rlabel metal1 37490 12104 37490 12104 0 _0769_
rlabel metal2 35006 16422 35006 16422 0 _0770_
rlabel metal1 38916 14382 38916 14382 0 _0771_
rlabel metal1 38318 15062 38318 15062 0 _0772_
rlabel metal1 39054 12852 39054 12852 0 _0773_
rlabel metal2 36846 13634 36846 13634 0 _0774_
rlabel metal1 37398 14382 37398 14382 0 _0775_
rlabel metal2 39054 14382 39054 14382 0 _0776_
rlabel metal1 38732 17238 38732 17238 0 _0777_
rlabel metal2 32338 16320 32338 16320 0 _0778_
rlabel metal1 36892 15130 36892 15130 0 _0779_
rlabel metal2 36662 19822 36662 19822 0 _0780_
rlabel metal2 39468 31314 39468 31314 0 _0781_
rlabel metal2 39698 29580 39698 29580 0 _0782_
rlabel metal3 38157 21964 38157 21964 0 _0783_
rlabel metal1 36156 22066 36156 22066 0 _0784_
rlabel metal1 36432 20978 36432 20978 0 _0785_
rlabel metal1 36110 23290 36110 23290 0 _0786_
rlabel metal1 37260 13294 37260 13294 0 _0787_
rlabel metal2 37490 14450 37490 14450 0 _0788_
rlabel metal2 37766 17578 37766 17578 0 _0789_
rlabel metal2 37766 15572 37766 15572 0 _0790_
rlabel metal1 38088 16966 38088 16966 0 _0791_
rlabel metal1 33166 14416 33166 14416 0 _0792_
rlabel metal1 36524 18938 36524 18938 0 _0793_
rlabel metal1 36616 20026 36616 20026 0 _0794_
rlabel metal1 37950 20434 37950 20434 0 _0795_
rlabel metal1 34730 17850 34730 17850 0 _0796_
rlabel metal2 38502 16354 38502 16354 0 _0797_
rlabel metal1 31786 14484 31786 14484 0 _0798_
rlabel metal1 34868 17510 34868 17510 0 _0799_
rlabel metal1 38364 24174 38364 24174 0 _0800_
rlabel metal1 39330 17510 39330 17510 0 _0801_
rlabel metal2 36662 25024 36662 25024 0 _0802_
rlabel metal1 34914 28424 34914 28424 0 _0803_
rlabel metal1 37812 24378 37812 24378 0 _0804_
rlabel metal2 37674 27642 37674 27642 0 _0805_
rlabel metal1 38088 24174 38088 24174 0 _0806_
rlabel metal1 38778 19822 38778 19822 0 _0807_
rlabel metal2 39422 27438 39422 27438 0 _0808_
rlabel metal1 38456 23154 38456 23154 0 _0809_
rlabel metal2 37720 19482 37720 19482 0 _0810_
rlabel metal1 38088 19482 38088 19482 0 _0811_
rlabel metal1 37720 22950 37720 22950 0 _0812_
rlabel metal1 40066 19856 40066 19856 0 _0813_
rlabel metal1 37904 20910 37904 20910 0 _0814_
rlabel metal1 36294 12784 36294 12784 0 _0815_
rlabel metal2 35650 18530 35650 18530 0 _0816_
rlabel metal1 35144 20230 35144 20230 0 _0817_
rlabel metal2 35374 18428 35374 18428 0 _0818_
rlabel metal1 37536 21114 37536 21114 0 _0819_
rlabel metal1 37766 21012 37766 21012 0 _0820_
rlabel metal1 36018 19448 36018 19448 0 _0821_
rlabel metal2 38410 16422 38410 16422 0 _0822_
rlabel metal2 37582 18513 37582 18513 0 _0823_
rlabel metal2 37582 19890 37582 19890 0 _0824_
rlabel via1 38502 20978 38502 20978 0 _0825_
rlabel metal1 28198 27982 28198 27982 0 _0826_
rlabel metal1 33902 28492 33902 28492 0 _0827_
rlabel metal1 34132 28526 34132 28526 0 _0828_
rlabel metal1 36570 22202 36570 22202 0 _0829_
rlabel metal2 34546 17884 34546 17884 0 _0830_
rlabel metal1 34914 16966 34914 16966 0 _0831_
rlabel metal1 36708 17170 36708 17170 0 _0832_
rlabel metal1 38824 20910 38824 20910 0 _0833_
rlabel metal1 39146 20774 39146 20774 0 _0834_
rlabel metal2 37858 18836 37858 18836 0 _0835_
rlabel metal1 36938 16422 36938 16422 0 _0836_
rlabel metal1 37490 19822 37490 19822 0 _0837_
rlabel metal1 38364 20026 38364 20026 0 _0838_
rlabel metal1 38732 16014 38732 16014 0 _0839_
rlabel metal1 35374 13974 35374 13974 0 _0840_
rlabel metal2 38226 15878 38226 15878 0 _0841_
rlabel metal1 38732 18666 38732 18666 0 _0842_
rlabel metal1 36202 13260 36202 13260 0 _0843_
rlabel metal1 35788 18122 35788 18122 0 _0844_
rlabel metal1 35420 17306 35420 17306 0 _0845_
rlabel metal1 37674 18598 37674 18598 0 _0846_
rlabel metal1 37628 18394 37628 18394 0 _0847_
rlabel metal2 39054 18496 39054 18496 0 _0848_
rlabel metal1 37260 17306 37260 17306 0 _0849_
rlabel metal1 37168 11730 37168 11730 0 _0850_
rlabel metal1 28750 14416 28750 14416 0 _0851_
rlabel metal1 36432 14586 36432 14586 0 _0852_
rlabel metal1 37260 17646 37260 17646 0 _0853_
rlabel metal1 38686 17782 38686 17782 0 _0854_
rlabel via2 39330 18955 39330 18955 0 _0855_
rlabel metal1 39468 29682 39468 29682 0 _0856_
rlabel metal1 35006 29274 35006 29274 0 _0857_
rlabel metal1 39652 21522 39652 21522 0 _0858_
rlabel metal2 36846 28118 36846 28118 0 _0859_
rlabel metal1 40066 22032 40066 22032 0 _0860_
rlabel metal1 35742 21114 35742 21114 0 _0861_
rlabel metal1 37858 21964 37858 21964 0 _0862_
rlabel metal1 37582 21998 37582 21998 0 _0863_
rlabel metal1 38272 21522 38272 21522 0 _0864_
rlabel metal1 38824 21658 38824 21658 0 _0865_
rlabel metal2 40066 20162 40066 20162 0 _0866_
rlabel metal1 37812 20298 37812 20298 0 _0867_
rlabel metal1 39284 17306 39284 17306 0 _0868_
rlabel metal1 39330 22746 39330 22746 0 _0869_
rlabel metal1 38962 20434 38962 20434 0 _0870_
rlabel metal1 39744 20570 39744 20570 0 _0871_
rlabel metal1 40480 21114 40480 21114 0 _0872_
rlabel metal2 39698 21590 39698 21590 0 _0873_
rlabel metal1 36110 28050 36110 28050 0 _0874_
rlabel metal1 37214 21590 37214 21590 0 _0875_
rlabel metal1 39514 21420 39514 21420 0 _0876_
rlabel metal1 40388 21658 40388 21658 0 _0877_
rlabel metal2 40066 26690 40066 26690 0 _0878_
rlabel metal2 40250 25024 40250 25024 0 _0879_
rlabel metal2 32430 22542 32430 22542 0 _0880_
rlabel metal2 36846 22882 36846 22882 0 _0881_
rlabel metal1 40158 23188 40158 23188 0 _0882_
rlabel metal2 31786 15878 31786 15878 0 _0883_
rlabel metal1 39238 19210 39238 19210 0 _0884_
rlabel metal1 43056 32402 43056 32402 0 _0885_
rlabel metal1 39652 18394 39652 18394 0 _0886_
rlabel metal2 40204 21012 40204 21012 0 _0887_
rlabel metal1 35650 25228 35650 25228 0 _0888_
rlabel via3 37421 32300 37421 32300 0 _0889_
rlabel metal1 39284 23290 39284 23290 0 _0890_
rlabel metal2 39054 24174 39054 24174 0 _0891_
rlabel metal2 39698 24004 39698 24004 0 _0892_
rlabel metal3 40641 33252 40641 33252 0 _0893_
rlabel metal2 39330 35530 39330 35530 0 _0894_
rlabel metal2 31786 35190 31786 35190 0 _0895_
rlabel metal1 29762 36040 29762 36040 0 _0896_
rlabel metal1 39882 32402 39882 32402 0 _0897_
rlabel metal1 38318 33422 38318 33422 0 _0898_
rlabel metal1 37858 33354 37858 33354 0 _0899_
rlabel metal2 38502 32096 38502 32096 0 _0900_
rlabel metal1 37904 33490 37904 33490 0 _0901_
rlabel metal1 21528 36686 21528 36686 0 _0902_
rlabel metal1 34684 27846 34684 27846 0 _0903_
rlabel metal1 30498 37944 30498 37944 0 _0904_
rlabel metal1 23506 36244 23506 36244 0 _0905_
rlabel metal1 27508 36074 27508 36074 0 _0906_
rlabel metal1 28566 33490 28566 33490 0 _0907_
rlabel metal1 23828 35666 23828 35666 0 _0908_
rlabel metal1 23736 38318 23736 38318 0 _0909_
rlabel metal1 23230 35802 23230 35802 0 _0910_
rlabel metal1 24610 35258 24610 35258 0 _0911_
rlabel metal1 27002 37196 27002 37196 0 _0912_
rlabel metal1 19182 40018 19182 40018 0 _0913_
rlabel metal2 21942 37468 21942 37468 0 _0914_
rlabel metal2 22218 35700 22218 35700 0 _0915_
rlabel metal2 21022 38284 21022 38284 0 _0916_
rlabel metal1 21436 35258 21436 35258 0 _0917_
rlabel metal1 21758 38318 21758 38318 0 _0918_
rlabel metal1 22632 36890 22632 36890 0 _0919_
rlabel metal1 24058 37366 24058 37366 0 _0920_
rlabel metal1 24150 34170 24150 34170 0 _0921_
rlabel metal2 26450 37060 26450 37060 0 _0922_
rlabel metal1 27048 35462 27048 35462 0 _0923_
rlabel metal1 28014 37298 28014 37298 0 _0924_
rlabel metal1 28382 33626 28382 33626 0 _0925_
rlabel metal1 28934 36686 28934 36686 0 _0926_
rlabel metal1 29164 35802 29164 35802 0 _0927_
rlabel metal1 33396 35258 33396 35258 0 _0928_
rlabel metal1 32798 36040 32798 36040 0 _0929_
rlabel metal2 32706 36550 32706 36550 0 _0930_
rlabel metal2 33350 38794 33350 38794 0 _0931_
rlabel metal1 32982 36890 32982 36890 0 _0932_
rlabel metal2 32338 38182 32338 38182 0 _0933_
rlabel metal2 31786 38386 31786 38386 0 _0934_
rlabel metal1 35558 38522 35558 38522 0 _0935_
rlabel metal1 37122 37978 37122 37978 0 _0936_
rlabel metal1 37582 36890 37582 36890 0 _0937_
rlabel metal2 36938 37604 36938 37604 0 _0938_
rlabel metal2 38962 36482 38962 36482 0 _0939_
rlabel metal1 25530 35054 25530 35054 0 _0940_
rlabel metal1 30314 35700 30314 35700 0 _0941_
rlabel metal1 26082 35122 26082 35122 0 _0942_
rlabel metal1 33028 35734 33028 35734 0 _0943_
rlabel metal1 25346 35088 25346 35088 0 _0944_
rlabel metal1 24702 33626 24702 33626 0 _0945_
rlabel metal1 23644 32742 23644 32742 0 _0946_
rlabel metal1 23000 34578 23000 34578 0 _0947_
rlabel metal1 25346 33626 25346 33626 0 _0948_
rlabel metal2 32522 35105 32522 35105 0 _0949_
rlabel metal1 25300 34578 25300 34578 0 _0950_
rlabel metal1 25806 34000 25806 34000 0 _0951_
rlabel metal1 23598 34102 23598 34102 0 _0952_
rlabel metal1 33994 33966 33994 33966 0 _0953_
rlabel metal2 33534 33150 33534 33150 0 _0954_
rlabel metal1 33813 32538 33813 32538 0 _0955_
rlabel metal2 20654 33677 20654 33677 0 _0956_
rlabel metal1 29532 34170 29532 34170 0 _0957_
rlabel metal1 29302 34408 29302 34408 0 _0958_
rlabel metal2 29394 35020 29394 35020 0 _0959_
rlabel metal1 10166 36142 10166 36142 0 _0960_
rlabel metal2 27094 33524 27094 33524 0 _0961_
rlabel metal1 27278 34102 27278 34102 0 _0962_
rlabel metal1 28152 34578 28152 34578 0 _0963_
rlabel metal2 28014 34748 28014 34748 0 _0964_
rlabel metal2 21022 24786 21022 24786 0 _0965_
rlabel metal1 21850 13260 21850 13260 0 _0966_
rlabel metal2 30590 21046 30590 21046 0 _0967_
rlabel metal1 19864 21862 19864 21862 0 _0968_
rlabel metal1 19504 21862 19504 21862 0 _0969_
rlabel metal1 20930 13804 20930 13804 0 _0970_
rlabel metal2 22494 12954 22494 12954 0 _0971_
rlabel metal2 33074 25993 33074 25993 0 clk
rlabel metal1 21022 21998 21022 21998 0 clknet_0_clk
rlabel metal1 20102 18734 20102 18734 0 clknet_4_0_0_clk
rlabel metal1 21160 41582 21160 41582 0 clknet_4_10_0_clk
rlabel metal1 25024 41582 25024 41582 0 clknet_4_11_0_clk
rlabel metal2 17066 33014 17066 33014 0 clknet_4_12_0_clk
rlabel metal1 36524 41582 36524 41582 0 clknet_4_13_0_clk
rlabel metal1 40250 42058 40250 42058 0 clknet_4_14_0_clk
rlabel metal2 34086 37570 34086 37570 0 clknet_4_15_0_clk
rlabel metal1 22034 17204 22034 17204 0 clknet_4_1_0_clk
rlabel metal2 15870 20366 15870 20366 0 clknet_4_2_0_clk
rlabel metal2 22034 20638 22034 20638 0 clknet_4_3_0_clk
rlabel metal1 26818 18190 26818 18190 0 clknet_4_4_0_clk
rlabel metal1 28888 13838 28888 13838 0 clknet_4_5_0_clk
rlabel metal2 40342 21794 40342 21794 0 clknet_4_6_0_clk
rlabel metal1 40250 13294 40250 13294 0 clknet_4_7_0_clk
rlabel metal3 19228 31756 19228 31756 0 clknet_4_8_0_clk
rlabel metal1 24932 41990 24932 41990 0 clknet_4_9_0_clk
rlabel metal1 43700 2414 43700 2414 0 io_in[0]
rlabel via2 43378 5899 43378 5899 0 io_in[1]
rlabel metal1 43700 10030 43700 10030 0 io_in[2]
rlabel metal3 43524 13260 43524 13260 0 io_in[3]
rlabel metal1 42458 10778 42458 10778 0 io_in[4]
rlabel metal1 43332 20842 43332 20842 0 io_in[5]
rlabel metal1 43654 24174 43654 24174 0 io_in[6]
rlabel metal1 43424 39814 43424 39814 0 io_in[7]
rlabel metal2 18170 31059 18170 31059 0 io_in[8]
rlabel via2 14122 36635 14122 36635 0 io_in[9]
rlabel metal1 42872 41582 42872 41582 0 io_oeb
rlabel metal2 1334 40028 1334 40028 0 io_out[0]
rlabel metal1 19550 36210 19550 36210 0 io_out[10]
rlabel metal1 18952 37774 18952 37774 0 io_out[11]
rlabel metal2 20148 41684 20148 41684 0 io_out[12]
rlabel metal1 21528 41106 21528 41106 0 io_out[13]
rlabel metal2 23230 42827 23230 42827 0 io_out[14]
rlabel metal2 24840 44132 24840 44132 0 io_out[15]
rlabel metal2 27646 39134 27646 39134 0 io_out[16]
rlabel metal1 28612 41038 28612 41038 0 io_out[17]
rlabel metal1 30636 44098 30636 44098 0 io_out[18]
rlabel metal2 31050 42827 31050 42827 0 io_out[19]
rlabel metal2 2898 39688 2898 39688 0 io_out[1]
rlabel metal2 32660 42092 32660 42092 0 io_out[20]
rlabel metal1 34408 44098 34408 44098 0 io_out[21]
rlabel metal2 35742 44193 35742 44193 0 io_out[22]
rlabel metal1 37674 40426 37674 40426 0 io_out[23]
rlabel metal1 39284 40358 39284 40358 0 io_out[24]
rlabel metal1 40020 41446 40020 41446 0 io_out[25]
rlabel metal1 42044 41786 42044 41786 0 io_out[26]
rlabel metal2 4554 42092 4554 42092 0 io_out[2]
rlabel metal2 6026 39756 6026 39756 0 io_out[3]
rlabel metal2 7590 39365 7590 39365 0 io_out[4]
rlabel metal2 9706 38216 9706 38216 0 io_out[5]
rlabel metal2 10718 39093 10718 39093 0 io_out[6]
rlabel metal2 12282 39637 12282 39637 0 io_out[7]
rlabel metal1 43056 2482 43056 2482 0 net1
rlabel metal1 42090 33524 42090 33524 0 net10
rlabel metal1 42964 42126 42964 42126 0 net11
rlabel metal1 14076 42194 14076 42194 0 net12
rlabel metal1 15456 42194 15456 42194 0 net13
rlabel metal1 36432 41990 36432 41990 0 net2
rlabel metal2 43010 11526 43010 11526 0 net3
rlabel metal1 43102 9078 43102 9078 0 net4
rlabel metal1 42044 10438 42044 10438 0 net5
rlabel metal2 17250 37927 17250 37927 0 net6
rlabel metal1 42366 9894 42366 9894 0 net7
rlabel metal1 43470 10778 43470 10778 0 net8
rlabel metal2 35282 33337 35282 33337 0 net9
rlabel metal1 41308 42194 41308 42194 0 rst
<< properties >>
string FIXED_BBOX 0 0 45000 45000
<< end >>
