VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END io_in[8]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 1.910 8.880 344.080 337.920 ;
      LAYER met2 ;
        RECT 1.930 4.280 341.220 339.845 ;
        RECT 1.930 3.670 15.910 4.280 ;
        RECT 16.750 3.670 47.650 4.280 ;
        RECT 48.490 3.670 79.390 4.280 ;
        RECT 80.230 3.670 111.130 4.280 ;
        RECT 111.970 3.670 142.870 4.280 ;
        RECT 143.710 3.670 174.610 4.280 ;
        RECT 175.450 3.670 206.350 4.280 ;
        RECT 207.190 3.670 238.090 4.280 ;
        RECT 238.930 3.670 269.830 4.280 ;
        RECT 270.670 3.670 301.570 4.280 ;
        RECT 302.410 3.670 333.310 4.280 ;
        RECT 334.150 3.670 341.220 4.280 ;
      LAYER met3 ;
        RECT 4.400 338.960 331.135 339.825 ;
        RECT 1.905 328.120 331.135 338.960 ;
        RECT 4.400 326.720 331.135 328.120 ;
        RECT 1.905 315.880 331.135 326.720 ;
        RECT 4.400 314.480 331.135 315.880 ;
        RECT 1.905 303.640 331.135 314.480 ;
        RECT 4.400 302.240 331.135 303.640 ;
        RECT 1.905 291.400 331.135 302.240 ;
        RECT 4.400 290.000 331.135 291.400 ;
        RECT 1.905 279.160 331.135 290.000 ;
        RECT 4.400 277.760 331.135 279.160 ;
        RECT 1.905 266.920 331.135 277.760 ;
        RECT 4.400 265.520 331.135 266.920 ;
        RECT 1.905 254.680 331.135 265.520 ;
        RECT 4.400 253.280 331.135 254.680 ;
        RECT 1.905 242.440 331.135 253.280 ;
        RECT 4.400 241.040 331.135 242.440 ;
        RECT 1.905 230.200 331.135 241.040 ;
        RECT 4.400 228.800 331.135 230.200 ;
        RECT 1.905 217.960 331.135 228.800 ;
        RECT 4.400 216.560 331.135 217.960 ;
        RECT 1.905 205.720 331.135 216.560 ;
        RECT 4.400 204.320 331.135 205.720 ;
        RECT 1.905 193.480 331.135 204.320 ;
        RECT 4.400 192.080 331.135 193.480 ;
        RECT 1.905 181.240 331.135 192.080 ;
        RECT 4.400 179.840 331.135 181.240 ;
        RECT 1.905 169.000 331.135 179.840 ;
        RECT 4.400 167.600 331.135 169.000 ;
        RECT 1.905 156.760 331.135 167.600 ;
        RECT 4.400 155.360 331.135 156.760 ;
        RECT 1.905 144.520 331.135 155.360 ;
        RECT 4.400 143.120 331.135 144.520 ;
        RECT 1.905 132.280 331.135 143.120 ;
        RECT 4.400 130.880 331.135 132.280 ;
        RECT 1.905 120.040 331.135 130.880 ;
        RECT 4.400 118.640 331.135 120.040 ;
        RECT 1.905 107.800 331.135 118.640 ;
        RECT 4.400 106.400 331.135 107.800 ;
        RECT 1.905 95.560 331.135 106.400 ;
        RECT 4.400 94.160 331.135 95.560 ;
        RECT 1.905 83.320 331.135 94.160 ;
        RECT 4.400 81.920 331.135 83.320 ;
        RECT 1.905 71.080 331.135 81.920 ;
        RECT 4.400 69.680 331.135 71.080 ;
        RECT 1.905 58.840 331.135 69.680 ;
        RECT 4.400 57.440 331.135 58.840 ;
        RECT 1.905 46.600 331.135 57.440 ;
        RECT 4.400 45.200 331.135 46.600 ;
        RECT 1.905 34.360 331.135 45.200 ;
        RECT 4.400 32.960 331.135 34.360 ;
        RECT 1.905 22.120 331.135 32.960 ;
        RECT 4.400 20.720 331.135 22.120 ;
        RECT 1.905 9.880 331.135 20.720 ;
        RECT 4.400 9.015 331.135 9.880 ;
      LAYER met4 ;
        RECT 3.055 15.815 20.640 335.065 ;
        RECT 23.040 15.815 97.440 335.065 ;
        RECT 99.840 15.815 174.240 335.065 ;
        RECT 176.640 15.815 251.040 335.065 ;
        RECT 253.440 15.815 283.065 335.065 ;
  END
END wrapped_as2650
END LIBRARY

