magic
tech sky130B
magscale 1 2
timestamp 1682093612
<< obsli1 >>
rect 1104 2159 10856 15793
<< obsm1 >>
rect 750 2128 11118 15824
<< metal2 >>
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
<< obsm2 >>
rect 756 856 11112 16561
rect 866 800 2170 856
rect 2338 800 3642 856
rect 3810 800 5114 856
rect 5282 800 6586 856
rect 6754 800 8058 856
rect 8226 800 9530 856
rect 9698 800 11002 856
<< metal3 >>
rect 0 16464 800 16584
rect 0 14288 800 14408
rect 0 12112 800 12232
rect 0 9936 800 10056
rect 0 7760 800 7880
rect 0 5584 800 5704
rect 0 3408 800 3528
rect 0 1232 800 1352
<< obsm3 >>
rect 880 16384 11014 16557
rect 800 14488 11014 16384
rect 880 14208 11014 14488
rect 800 12312 11014 14208
rect 880 12032 11014 12312
rect 800 10136 11014 12032
rect 880 9856 11014 10136
rect 800 7960 11014 9856
rect 880 7680 11014 7960
rect 800 5784 11014 7680
rect 880 5504 11014 5784
rect 800 3608 11014 5504
rect 880 3328 11014 3608
rect 800 1432 11014 3328
rect 880 1259 11014 1432
<< metal4 >>
rect 2163 2128 2483 15824
rect 3382 2128 3702 15824
rect 4601 2128 4921 15824
rect 5820 2128 6140 15824
rect 7039 2128 7359 15824
rect 8258 2128 8578 15824
rect 9477 2128 9797 15824
rect 10696 2128 11016 15824
<< labels >>
rlabel metal3 s 0 1232 800 1352 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 io_in[7]
port 8 nsew signal input
rlabel metal2 s 754 0 810 800 6 io_out[0]
port 9 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 io_out[1]
port 10 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 io_out[2]
port 11 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 io_out[3]
port 12 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 io_out[4]
port 13 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 io_out[5]
port 14 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 io_out[6]
port 15 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 io_out[7]
port 16 nsew signal output
rlabel metal4 s 2163 2128 2483 15824 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 15824 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 15824 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 15824 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 3382 2128 3702 15824 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 5820 2128 6140 15824 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 8258 2128 8578 15824 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 10696 2128 11016 15824 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 533758
string GDS_FILE /run/media/tholin/Data/Projects/MPW/TMBoC/openlane/4x4-multiply/runs/23_04_21_18_13/results/signoff/tt2_tholin_multiplier.magic.gds
string GDS_START 232398
<< end >>

