magic
tech sky130B
magscale 1 2
timestamp 1683541604
<< viali >>
rect 4169 15453 4203 15487
rect 10701 15453 10735 15487
rect 14473 15453 14507 15487
rect 15025 15453 15059 15487
rect 4077 15317 4111 15351
rect 10793 15317 10827 15351
rect 14381 15317 14415 15351
rect 15117 15317 15151 15351
rect 4638 14977 4672 15011
rect 4905 14977 4939 15011
rect 6745 14977 6779 15011
rect 9689 14977 9723 15011
rect 10609 14977 10643 15011
rect 11897 14977 11931 15011
rect 12541 14977 12575 15011
rect 13829 14977 13863 15011
rect 14473 14977 14507 15011
rect 15117 14977 15151 15011
rect 15761 14977 15795 15011
rect 3525 14773 3559 14807
rect 6653 14773 6687 14807
rect 9597 14773 9631 14807
rect 10517 14773 10551 14807
rect 11805 14773 11839 14807
rect 12449 14773 12483 14807
rect 13737 14773 13771 14807
rect 14381 14773 14415 14807
rect 15025 14773 15059 14807
rect 15669 14773 15703 14807
rect 7389 14501 7423 14535
rect 5917 14433 5951 14467
rect 11989 14433 12023 14467
rect 12265 14433 12299 14467
rect 14289 14433 14323 14467
rect 16037 14433 16071 14467
rect 2789 14365 2823 14399
rect 4169 14365 4203 14399
rect 4261 14365 4295 14399
rect 5641 14365 5675 14399
rect 9137 14365 9171 14399
rect 9413 14365 9447 14399
rect 10241 14365 10275 14399
rect 13461 14365 13495 14399
rect 16313 14365 16347 14399
rect 3985 14297 4019 14331
rect 2697 14229 2731 14263
rect 9229 14229 9263 14263
rect 13369 14229 13403 14263
rect 5917 14025 5951 14059
rect 6653 14025 6687 14059
rect 2513 13957 2547 13991
rect 13369 13957 13403 13991
rect 15117 13957 15151 13991
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 9505 13889 9539 13923
rect 10425 13889 10459 13923
rect 12449 13889 12483 13923
rect 13093 13889 13127 13923
rect 15761 13889 15795 13923
rect 2237 13821 2271 13855
rect 3985 13821 4019 13855
rect 9229 13821 9263 13855
rect 12265 13821 12299 13855
rect 12633 13821 12667 13855
rect 7757 13685 7791 13719
rect 10333 13685 10367 13719
rect 15669 13685 15703 13719
rect 2513 13481 2547 13515
rect 4169 13481 4203 13515
rect 4353 13481 4387 13515
rect 8493 13481 8527 13515
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 11897 13345 11931 13379
rect 14565 13345 14599 13379
rect 16313 13345 16347 13379
rect 2605 13277 2639 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 14289 13277 14323 13311
rect 3985 13209 4019 13243
rect 4185 13141 4219 13175
rect 7021 12937 7055 12971
rect 7297 12937 7331 12971
rect 8125 12937 8159 12971
rect 11805 12937 11839 12971
rect 14749 12937 14783 12971
rect 15393 12937 15427 12971
rect 7389 12869 7423 12903
rect 2237 12801 2271 12835
rect 2697 12801 2731 12835
rect 5181 12801 5215 12835
rect 7205 12801 7239 12835
rect 8033 12801 8067 12835
rect 11897 12801 11931 12835
rect 14841 12801 14875 12835
rect 15301 12801 15335 12835
rect 2789 12733 2823 12767
rect 4905 12733 4939 12767
rect 7573 12665 7607 12699
rect 2145 12597 2179 12631
rect 3433 12597 3467 12631
rect 6837 12393 6871 12427
rect 4169 12325 4203 12359
rect 1869 12257 1903 12291
rect 1593 12189 1627 12223
rect 4169 12189 4203 12223
rect 4353 12189 4387 12223
rect 6101 12189 6135 12223
rect 6929 12189 6963 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 3341 12053 3375 12087
rect 6193 12053 6227 12087
rect 7481 12053 7515 12087
rect 2421 11849 2455 11883
rect 2973 11781 3007 11815
rect 6837 11781 6871 11815
rect 2513 11713 2547 11747
rect 3157 11713 3191 11747
rect 3341 11713 3375 11747
rect 6009 11713 6043 11747
rect 6561 11713 6595 11747
rect 8953 11713 8987 11747
rect 9137 11713 9171 11747
rect 10885 11713 10919 11747
rect 11897 11713 11931 11747
rect 12541 11713 12575 11747
rect 14841 11713 14875 11747
rect 16037 11713 16071 11747
rect 8953 11577 8987 11611
rect 12449 11577 12483 11611
rect 5917 11509 5951 11543
rect 8309 11509 8343 11543
rect 10793 11509 10827 11543
rect 11805 11509 11839 11543
rect 14933 11509 14967 11543
rect 16129 11509 16163 11543
rect 8033 11237 8067 11271
rect 6561 11169 6595 11203
rect 9781 11169 9815 11203
rect 11805 11169 11839 11203
rect 16037 11169 16071 11203
rect 6285 11101 6319 11135
rect 13645 11101 13679 11135
rect 14289 11101 14323 11135
rect 16313 11101 16347 11135
rect 10057 11033 10091 11067
rect 13553 11033 13587 11067
rect 6653 10761 6687 10795
rect 7665 10761 7699 10795
rect 15301 10761 15335 10795
rect 11161 10693 11195 10727
rect 6745 10625 6779 10659
rect 8953 10625 8987 10659
rect 9413 10625 9447 10659
rect 15393 10625 15427 10659
rect 15853 10625 15887 10659
rect 12265 10557 12299 10591
rect 12541 10557 12575 10591
rect 14289 10557 14323 10591
rect 15945 10421 15979 10455
rect 10057 10217 10091 10251
rect 13277 10217 13311 10251
rect 5273 10081 5307 10115
rect 10609 10081 10643 10115
rect 10885 10081 10919 10115
rect 12633 10081 12667 10115
rect 14289 10081 14323 10115
rect 16313 10081 16347 10115
rect 2421 10013 2455 10047
rect 3249 10013 3283 10047
rect 3433 10013 3467 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 8401 10013 8435 10047
rect 9505 10013 9539 10047
rect 10149 10013 10183 10047
rect 13369 10013 13403 10047
rect 3985 9945 4019 9979
rect 7021 9945 7055 9979
rect 16037 9945 16071 9979
rect 2513 9877 2547 9911
rect 3341 9877 3375 9911
rect 8493 9877 8527 9911
rect 9413 9877 9447 9911
rect 2697 9605 2731 9639
rect 8861 9605 8895 9639
rect 11897 9605 11931 9639
rect 12541 9605 12575 9639
rect 16129 9605 16163 9639
rect 1961 9537 1995 9571
rect 4813 9537 4847 9571
rect 4997 9537 5031 9571
rect 5641 9537 5675 9571
rect 6009 9537 6043 9571
rect 6837 9537 6871 9571
rect 7047 9537 7081 9571
rect 7941 9537 7975 9571
rect 11989 9537 12023 9571
rect 12449 9537 12483 9571
rect 15393 9537 15427 9571
rect 16037 9537 16071 9571
rect 2421 9469 2455 9503
rect 5825 9469 5859 9503
rect 7205 9469 7239 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 10333 9469 10367 9503
rect 15485 9401 15519 9435
rect 1869 9333 1903 9367
rect 4169 9333 4203 9367
rect 4905 9333 4939 9367
rect 5917 9333 5951 9367
rect 6837 9333 6871 9367
rect 1593 8993 1627 9027
rect 6653 8925 6687 8959
rect 7021 8925 7055 8959
rect 7389 8925 7423 8959
rect 7757 8925 7791 8959
rect 11069 8925 11103 8959
rect 14473 8925 14507 8959
rect 1869 8857 1903 8891
rect 5089 8857 5123 8891
rect 5181 8857 5215 8891
rect 5549 8857 5583 8891
rect 5917 8857 5951 8891
rect 8033 8857 8067 8891
rect 3341 8789 3375 8823
rect 4813 8789 4847 8823
rect 6101 8789 6135 8823
rect 9781 8789 9815 8823
rect 14381 8789 14415 8823
rect 2513 8585 2547 8619
rect 7481 8585 7515 8619
rect 10241 8585 10275 8619
rect 7665 8517 7699 8551
rect 8953 8517 8987 8551
rect 2605 8449 2639 8483
rect 12633 8449 12667 8483
rect 15117 8449 15151 8483
rect 12909 8381 12943 8415
rect 14657 8381 14691 8415
rect 8033 8313 8067 8347
rect 7665 8245 7699 8279
rect 15209 8245 15243 8279
rect 13645 8041 13679 8075
rect 5733 7973 5767 8007
rect 16313 7905 16347 7939
rect 4169 7837 4203 7871
rect 7941 7837 7975 7871
rect 8401 7837 8435 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 10425 7837 10459 7871
rect 13737 7837 13771 7871
rect 7021 7769 7055 7803
rect 14289 7769 14323 7803
rect 16037 7769 16071 7803
rect 4077 7701 4111 7735
rect 7849 7701 7883 7735
rect 8493 7701 8527 7735
rect 9229 7701 9263 7735
rect 11713 7701 11747 7735
rect 2973 7497 3007 7531
rect 15301 7497 15335 7531
rect 15945 7497 15979 7531
rect 2881 7429 2915 7463
rect 9321 7429 9355 7463
rect 2145 7361 2179 7395
rect 2789 7361 2823 7395
rect 3617 7361 3651 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 9045 7361 9079 7395
rect 11713 7361 11747 7395
rect 14381 7361 14415 7395
rect 15393 7361 15427 7395
rect 15853 7361 15887 7395
rect 3157 7293 3191 7327
rect 3893 7293 3927 7327
rect 6745 7293 6779 7327
rect 7021 7293 7055 7327
rect 2605 7225 2639 7259
rect 8493 7225 8527 7259
rect 2053 7157 2087 7191
rect 4997 7157 5031 7191
rect 6009 7157 6043 7191
rect 10793 7157 10827 7191
rect 11805 7157 11839 7191
rect 14289 7157 14323 7191
rect 12369 6953 12403 6987
rect 2513 6817 2547 6851
rect 10241 6817 10275 6851
rect 10885 6817 10919 6851
rect 14289 6817 14323 6851
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 5089 6749 5123 6783
rect 6924 6749 6958 6783
rect 7297 6749 7331 6783
rect 8217 6749 8251 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 12633 6749 12667 6783
rect 13369 6749 13403 6783
rect 4813 6681 4847 6715
rect 5181 6681 5215 6715
rect 5549 6681 5583 6715
rect 7021 6681 7055 6715
rect 7113 6681 7147 6715
rect 14565 6681 14599 6715
rect 3157 6613 3191 6647
rect 5917 6613 5951 6647
rect 6101 6613 6135 6647
rect 6728 6613 6762 6647
rect 8125 6613 8159 6647
rect 13277 6613 13311 6647
rect 16037 6613 16071 6647
rect 3985 6409 4019 6443
rect 6561 6409 6595 6443
rect 8309 6409 8343 6443
rect 11805 6409 11839 6443
rect 12449 6409 12483 6443
rect 14473 6409 14507 6443
rect 15853 6409 15887 6443
rect 2513 6341 2547 6375
rect 9597 6341 9631 6375
rect 13338 6341 13372 6375
rect 1777 6273 1811 6307
rect 2237 6273 2271 6307
rect 6929 6273 6963 6307
rect 7021 6273 7055 6307
rect 11897 6273 11931 6307
rect 12357 6273 12391 6307
rect 13093 6273 13127 6307
rect 14933 6273 14967 6307
rect 15117 6273 15151 6307
rect 15761 6273 15795 6307
rect 7205 6205 7239 6239
rect 15209 6137 15243 6171
rect 1685 6069 1719 6103
rect 14565 5865 14599 5899
rect 2513 5661 2547 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 8585 5661 8619 5695
rect 9321 5661 9355 5695
rect 9413 5661 9447 5695
rect 14657 5661 14691 5695
rect 2421 5525 2455 5559
rect 3249 5525 3283 5559
rect 8493 5525 8527 5559
rect 9229 5525 9263 5559
rect 9965 5321 9999 5355
rect 2145 5253 2179 5287
rect 3893 5253 3927 5287
rect 8493 5253 8527 5287
rect 1869 5185 1903 5219
rect 4813 5185 4847 5219
rect 4997 5185 5031 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 7573 5185 7607 5219
rect 7665 5117 7699 5151
rect 8217 5117 8251 5151
rect 5457 5049 5491 5083
rect 4813 4981 4847 5015
rect 5641 4709 5675 4743
rect 14565 4709 14599 4743
rect 9505 4641 9539 4675
rect 14289 4641 14323 4675
rect 4721 4573 4755 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 6653 4573 6687 4607
rect 7297 4573 7331 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 9413 4573 9447 4607
rect 11897 4573 11931 4607
rect 13553 4573 13587 4607
rect 15853 4573 15887 4607
rect 4537 4505 4571 4539
rect 4905 4505 4939 4539
rect 5641 4505 5675 4539
rect 12081 4505 12115 4539
rect 16129 4505 16163 4539
rect 6745 4437 6779 4471
rect 7389 4437 7423 4471
rect 8493 4437 8527 4471
rect 11713 4437 11747 4471
rect 13645 4437 13679 4471
rect 14749 4437 14783 4471
rect 3525 4233 3559 4267
rect 4629 4233 4663 4267
rect 6653 4165 6687 4199
rect 7941 4165 7975 4199
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3801 4097 3835 4131
rect 4445 4097 4479 4131
rect 4721 4097 4755 4131
rect 5457 4097 5491 4131
rect 6561 4097 6595 4131
rect 7665 4097 7699 4131
rect 10977 4097 11011 4131
rect 12357 4097 12391 4131
rect 13001 4097 13035 4131
rect 13921 4097 13955 4131
rect 14177 4097 14211 4131
rect 15761 4097 15795 4131
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 5181 4029 5215 4063
rect 9689 4029 9723 4063
rect 13461 4029 13495 4063
rect 15945 4029 15979 4063
rect 3709 3961 3743 3995
rect 12081 3961 12115 3995
rect 13369 3961 13403 3995
rect 3065 3893 3099 3927
rect 5273 3893 5307 3927
rect 5641 3893 5675 3927
rect 11069 3893 11103 3927
rect 11897 3893 11931 3927
rect 15301 3893 15335 3927
rect 3341 3689 3375 3723
rect 6837 3689 6871 3723
rect 10517 3689 10551 3723
rect 12909 3689 12943 3723
rect 14289 3689 14323 3723
rect 4721 3621 4755 3655
rect 4813 3621 4847 3655
rect 12449 3621 12483 3655
rect 1961 3553 1995 3587
rect 2421 3553 2455 3587
rect 3433 3553 3467 3587
rect 13369 3553 13403 3587
rect 13553 3553 13587 3587
rect 15669 3553 15703 3587
rect 16221 3553 16255 3587
rect 2329 3485 2363 3519
rect 3157 3485 3191 3519
rect 4629 3485 4663 3519
rect 4905 3485 4939 3519
rect 5641 3485 5675 3519
rect 5825 3485 5859 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 6745 3485 6779 3519
rect 7021 3485 7055 3519
rect 9137 3485 9171 3519
rect 9404 3485 9438 3519
rect 11069 3485 11103 3519
rect 11336 3485 11370 3519
rect 15402 3485 15436 3519
rect 16129 3485 16163 3519
rect 2973 3349 3007 3383
rect 5089 3349 5123 3383
rect 6285 3349 6319 3383
rect 7205 3349 7239 3383
rect 13277 3349 13311 3383
rect 5089 3145 5123 3179
rect 6653 3145 6687 3179
rect 9321 3145 9355 3179
rect 11069 3145 11103 3179
rect 13921 3145 13955 3179
rect 14749 3145 14783 3179
rect 3433 3077 3467 3111
rect 4445 3077 4479 3111
rect 5457 3077 5491 3111
rect 14013 3077 14047 3111
rect 2053 3009 2087 3043
rect 3617 3009 3651 3043
rect 3801 3009 3835 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 5549 3009 5583 3043
rect 6745 3009 6779 3043
rect 9413 3009 9447 3043
rect 10977 3009 11011 3043
rect 11713 3009 11747 3043
rect 11980 3009 12014 3043
rect 15117 3009 15151 3043
rect 1777 2941 1811 2975
rect 4261 2941 4295 2975
rect 14197 2941 14231 2975
rect 15209 2941 15243 2975
rect 15301 2941 15335 2975
rect 13553 2873 13587 2907
rect 13093 2805 13127 2839
rect 14473 2601 14507 2635
rect 15025 2465 15059 2499
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 5365 2397 5399 2431
rect 6837 2397 6871 2431
rect 8125 2397 8159 2431
rect 9781 2397 9815 2431
rect 12173 2397 12207 2431
rect 13185 2397 13219 2431
rect 14841 2397 14875 2431
rect 14933 2397 14967 2431
rect 15669 2397 15703 2431
rect 2605 2329 2639 2363
rect 4261 2329 4295 2363
rect 5641 2329 5675 2363
rect 7113 2329 7147 2363
rect 8401 2329 8435 2363
rect 10057 2329 10091 2363
rect 11897 2329 11931 2363
rect 12909 2329 12943 2363
rect 15945 2329 15979 2363
<< metal1 >>
rect 13538 17280 13544 17332
rect 13596 17320 13602 17332
rect 14458 17320 14464 17332
rect 13596 17292 14464 17320
rect 13596 17280 13602 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 1104 15802 16836 15824
rect 1104 15750 2916 15802
rect 2968 15750 2980 15802
rect 3032 15750 3044 15802
rect 3096 15750 3108 15802
rect 3160 15750 3172 15802
rect 3224 15750 6849 15802
rect 6901 15750 6913 15802
rect 6965 15750 6977 15802
rect 7029 15750 7041 15802
rect 7093 15750 7105 15802
rect 7157 15750 10782 15802
rect 10834 15750 10846 15802
rect 10898 15750 10910 15802
rect 10962 15750 10974 15802
rect 11026 15750 11038 15802
rect 11090 15750 14715 15802
rect 14767 15750 14779 15802
rect 14831 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 16836 15802
rect 1104 15728 16836 15750
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 6270 15484 6276 15496
rect 4203 15456 6276 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 14458 15444 14464 15496
rect 14516 15444 14522 15496
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 15028 15416 15056 15447
rect 13872 15388 15056 15416
rect 13872 15376 13878 15388
rect 4065 15351 4123 15357
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4798 15348 4804 15360
rect 4111 15320 4804 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 10781 15351 10839 15357
rect 10781 15317 10793 15351
rect 10827 15348 10839 15351
rect 11974 15348 11980 15360
rect 10827 15320 11980 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 14148 15320 14381 15348
rect 14148 15308 14154 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14369 15311 14427 15317
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 16022 15348 16028 15360
rect 15151 15320 16028 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 1104 15258 16995 15280
rect 1104 15206 4882 15258
rect 4934 15206 4946 15258
rect 4998 15206 5010 15258
rect 5062 15206 5074 15258
rect 5126 15206 5138 15258
rect 5190 15206 8815 15258
rect 8867 15206 8879 15258
rect 8931 15206 8943 15258
rect 8995 15206 9007 15258
rect 9059 15206 9071 15258
rect 9123 15206 12748 15258
rect 12800 15206 12812 15258
rect 12864 15206 12876 15258
rect 12928 15206 12940 15258
rect 12992 15206 13004 15258
rect 13056 15206 16681 15258
rect 16733 15206 16745 15258
rect 16797 15206 16809 15258
rect 16861 15206 16873 15258
rect 16925 15206 16937 15258
rect 16989 15206 16995 15258
rect 1104 15184 16995 15206
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 4626 15011 4684 15017
rect 4626 15008 4638 15011
rect 4396 14980 4638 15008
rect 4396 14968 4402 14980
rect 4626 14977 4638 14980
rect 4672 14977 4684 15011
rect 4626 14971 4684 14977
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4856 14980 4905 15008
rect 4856 14968 4862 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7374 15008 7380 15020
rect 6779 14980 7380 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9692 14940 9720 14971
rect 10594 14968 10600 15020
rect 10652 14968 10658 15020
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 13814 14968 13820 15020
rect 13872 14968 13878 15020
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 15008 15163 15011
rect 15286 15008 15292 15020
rect 15151 14980 15292 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 11146 14940 11152 14952
rect 9692 14912 11152 14940
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 11900 14940 11928 14968
rect 14476 14940 14504 14971
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 15764 14940 15792 14971
rect 11900 14912 15792 14940
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 3970 14804 3976 14816
rect 3559 14776 3976 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 6641 14807 6699 14813
rect 6641 14804 6653 14807
rect 5960 14776 6653 14804
rect 5960 14764 5966 14776
rect 6641 14773 6653 14776
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 9585 14807 9643 14813
rect 9585 14804 9597 14807
rect 9548 14776 9597 14804
rect 9548 14764 9554 14776
rect 9585 14773 9597 14776
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 9858 14764 9864 14816
rect 9916 14804 9922 14816
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 9916 14776 10517 14804
rect 9916 14764 9922 14776
rect 10505 14773 10517 14776
rect 10551 14773 10563 14807
rect 10505 14767 10563 14773
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 11572 14776 11805 14804
rect 11572 14764 11578 14776
rect 11793 14773 11805 14776
rect 11839 14773 11851 14807
rect 11793 14767 11851 14773
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12308 14776 12449 14804
rect 12308 14764 12314 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13725 14807 13783 14813
rect 13725 14804 13737 14807
rect 13136 14776 13737 14804
rect 13136 14764 13142 14776
rect 13725 14773 13737 14776
rect 13771 14773 13783 14807
rect 13725 14767 13783 14773
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 15013 14807 15071 14813
rect 15013 14804 15025 14807
rect 14608 14776 15025 14804
rect 14608 14764 14614 14776
rect 15013 14773 15025 14776
rect 15059 14773 15071 14807
rect 15013 14767 15071 14773
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15620 14776 15669 14804
rect 15620 14764 15626 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 1104 14714 16836 14736
rect 1104 14662 2916 14714
rect 2968 14662 2980 14714
rect 3032 14662 3044 14714
rect 3096 14662 3108 14714
rect 3160 14662 3172 14714
rect 3224 14662 6849 14714
rect 6901 14662 6913 14714
rect 6965 14662 6977 14714
rect 7029 14662 7041 14714
rect 7093 14662 7105 14714
rect 7157 14662 10782 14714
rect 10834 14662 10846 14714
rect 10898 14662 10910 14714
rect 10962 14662 10974 14714
rect 11026 14662 11038 14714
rect 11090 14662 14715 14714
rect 14767 14662 14779 14714
rect 14831 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 16836 14714
rect 1104 14640 16836 14662
rect 4430 14560 4436 14612
rect 4488 14600 4494 14612
rect 8294 14600 8300 14612
rect 4488 14572 8300 14600
rect 4488 14560 4494 14572
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 7374 14492 7380 14544
rect 7432 14492 7438 14544
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4120 14436 4292 14464
rect 4120 14424 4126 14436
rect 4264 14405 4292 14436
rect 5902 14424 5908 14476
rect 5960 14424 5966 14476
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 8478 14464 8484 14476
rect 6604 14436 8484 14464
rect 6604 14424 6610 14436
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 11882 14464 11888 14476
rect 8536 14436 9168 14464
rect 8536 14424 8542 14436
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 4157 14399 4215 14405
rect 2823 14368 3924 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 2556 14232 2697 14260
rect 2556 14220 2562 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 3896 14260 3924 14368
rect 4157 14365 4169 14399
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 3970 14288 3976 14340
rect 4028 14288 4034 14340
rect 4172 14328 4200 14359
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 9140 14405 9168 14436
rect 9416 14436 11888 14464
rect 9416 14405 9444 14436
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 11974 14424 11980 14476
rect 12032 14424 12038 14476
rect 12250 14424 12256 14476
rect 12308 14424 12314 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14277 14467 14335 14473
rect 14277 14464 14289 14467
rect 13872 14436 14289 14464
rect 13872 14424 13878 14436
rect 14277 14433 14289 14436
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 16022 14424 16028 14476
rect 16080 14424 16086 14476
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10594 14396 10600 14408
rect 10275 14368 10600 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 12584 14368 13461 14396
rect 12584 14356 12590 14368
rect 13449 14365 13461 14368
rect 13495 14396 13507 14399
rect 14642 14396 14648 14408
rect 13495 14368 14648 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 16298 14356 16304 14408
rect 16356 14356 16362 14408
rect 4172 14300 4292 14328
rect 4154 14260 4160 14272
rect 3896 14232 4160 14260
rect 2685 14223 2743 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4264 14260 4292 14300
rect 6638 14288 6644 14340
rect 6696 14288 6702 14340
rect 11514 14288 11520 14340
rect 11572 14288 11578 14340
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 6730 14260 6736 14272
rect 4264 14232 6736 14260
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 9214 14220 9220 14272
rect 9272 14220 9278 14272
rect 13354 14220 13360 14272
rect 13412 14220 13418 14272
rect 1104 14170 16995 14192
rect 1104 14118 4882 14170
rect 4934 14118 4946 14170
rect 4998 14118 5010 14170
rect 5062 14118 5074 14170
rect 5126 14118 5138 14170
rect 5190 14118 8815 14170
rect 8867 14118 8879 14170
rect 8931 14118 8943 14170
rect 8995 14118 9007 14170
rect 9059 14118 9071 14170
rect 9123 14118 12748 14170
rect 12800 14118 12812 14170
rect 12864 14118 12876 14170
rect 12928 14118 12940 14170
rect 12992 14118 13004 14170
rect 13056 14118 16681 14170
rect 16733 14118 16745 14170
rect 16797 14118 16809 14170
rect 16861 14118 16873 14170
rect 16925 14118 16937 14170
rect 16989 14118 16995 14170
rect 1104 14096 16995 14118
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5684 14028 5917 14056
rect 5684 14016 5690 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 5905 14019 5963 14025
rect 6638 14016 6644 14068
rect 6696 14016 6702 14068
rect 2498 13948 2504 14000
rect 2556 13948 2562 14000
rect 3970 13988 3976 14000
rect 3726 13960 3976 13988
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 9214 13988 9220 14000
rect 8786 13960 9220 13988
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 13354 13948 13360 14000
rect 13412 13948 13418 14000
rect 14366 13948 14372 14000
rect 14424 13948 14430 14000
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 15105 13991 15163 13997
rect 15105 13988 15117 13991
rect 14700 13960 15117 13988
rect 14700 13948 14706 13960
rect 15105 13957 15117 13960
rect 15151 13957 15163 13991
rect 15105 13951 15163 13957
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 2222 13812 2228 13864
rect 2280 13812 2286 13864
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4154 13852 4160 13864
rect 4019 13824 4160 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 6012 13852 6040 13883
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 9490 13880 9496 13932
rect 9548 13880 9554 13932
rect 10413 13923 10471 13929
rect 10413 13889 10425 13923
rect 10459 13920 10471 13923
rect 11146 13920 11152 13932
rect 10459 13892 11152 13920
rect 10459 13889 10471 13892
rect 10413 13883 10471 13889
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 13078 13880 13084 13932
rect 13136 13880 13142 13932
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15528 13892 15761 13920
rect 15528 13880 15534 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 6012 13824 6914 13852
rect 6886 13716 6914 13824
rect 9214 13812 9220 13864
rect 9272 13812 9278 13864
rect 12250 13812 12256 13864
rect 12308 13812 12314 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 14090 13852 14096 13864
rect 12667 13824 14096 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 7745 13719 7803 13725
rect 7745 13716 7757 13719
rect 6886 13688 7757 13716
rect 7745 13685 7757 13688
rect 7791 13716 7803 13719
rect 7834 13716 7840 13728
rect 7791 13688 7840 13716
rect 7791 13685 7803 13688
rect 7745 13679 7803 13685
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 10192 13688 10333 13716
rect 10192 13676 10198 13688
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 15654 13676 15660 13728
rect 15712 13676 15718 13728
rect 1104 13626 16836 13648
rect 1104 13574 2916 13626
rect 2968 13574 2980 13626
rect 3032 13574 3044 13626
rect 3096 13574 3108 13626
rect 3160 13574 3172 13626
rect 3224 13574 6849 13626
rect 6901 13574 6913 13626
rect 6965 13574 6977 13626
rect 7029 13574 7041 13626
rect 7093 13574 7105 13626
rect 7157 13574 10782 13626
rect 10834 13574 10846 13626
rect 10898 13574 10910 13626
rect 10962 13574 10974 13626
rect 11026 13574 11038 13626
rect 11090 13574 14715 13626
rect 14767 13574 14779 13626
rect 14831 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 16836 13626
rect 1104 13552 16836 13574
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2501 13515 2559 13521
rect 2501 13512 2513 13515
rect 2280 13484 2513 13512
rect 2280 13472 2286 13484
rect 2501 13481 2513 13484
rect 2547 13481 2559 13515
rect 2501 13475 2559 13481
rect 4154 13472 4160 13524
rect 4212 13472 4218 13524
rect 4338 13472 4344 13524
rect 4396 13472 4402 13524
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 4172 13444 4200 13472
rect 4706 13444 4712 13456
rect 4172 13416 4712 13444
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11885 13379 11943 13385
rect 11885 13376 11897 13379
rect 11204 13348 11897 13376
rect 11204 13336 11210 13348
rect 11885 13345 11897 13348
rect 11931 13345 11943 13379
rect 11885 13339 11943 13345
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15344 13348 16313 13376
rect 15344 13336 15350 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2608 13240 2636 13271
rect 6270 13268 6276 13320
rect 6328 13268 6334 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13308 6423 13311
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6411 13280 6929 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 7064 13280 7205 13308
rect 7064 13268 7070 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 2774 13240 2780 13252
rect 2608 13212 2780 13240
rect 2774 13200 2780 13212
rect 2832 13240 2838 13252
rect 3970 13240 3976 13252
rect 2832 13212 3976 13240
rect 2832 13200 2838 13212
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 4173 13175 4231 13181
rect 4173 13172 4185 13175
rect 3936 13144 4185 13172
rect 3936 13132 3942 13144
rect 4173 13141 4185 13144
rect 4219 13141 4231 13175
rect 6288 13172 6316 13268
rect 11790 13240 11796 13252
rect 11362 13212 11796 13240
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 7650 13172 7656 13184
rect 6288 13144 7656 13172
rect 4173 13135 4231 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 1104 13082 16995 13104
rect 1104 13030 4882 13082
rect 4934 13030 4946 13082
rect 4998 13030 5010 13082
rect 5062 13030 5074 13082
rect 5126 13030 5138 13082
rect 5190 13030 8815 13082
rect 8867 13030 8879 13082
rect 8931 13030 8943 13082
rect 8995 13030 9007 13082
rect 9059 13030 9071 13082
rect 9123 13030 12748 13082
rect 12800 13030 12812 13082
rect 12864 13030 12876 13082
rect 12928 13030 12940 13082
rect 12992 13030 13004 13082
rect 13056 13030 16681 13082
rect 16733 13030 16745 13082
rect 16797 13030 16809 13082
rect 16861 13030 16873 13082
rect 16925 13030 16937 13082
rect 16989 13030 16995 13082
rect 1104 13008 16995 13030
rect 7006 12928 7012 12980
rect 7064 12928 7070 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7331 12940 8125 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 8113 12937 8125 12940
rect 8159 12968 8171 12971
rect 9214 12968 9220 12980
rect 8159 12940 9220 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14332 12940 14749 12968
rect 14332 12928 14338 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 16298 12968 16304 12980
rect 15427 12940 16304 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 2774 12900 2780 12912
rect 2240 12872 2780 12900
rect 2240 12841 2268 12872
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 4154 12860 4160 12912
rect 4212 12860 4218 12912
rect 7374 12900 7380 12912
rect 6886 12872 7380 12900
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 6546 12832 6552 12844
rect 5215 12804 6552 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 2498 12656 2504 12708
rect 2556 12696 2562 12708
rect 2700 12696 2728 12795
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 3878 12764 3884 12776
rect 2823 12736 3884 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3878 12724 3884 12736
rect 3936 12764 3942 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 3936 12736 4905 12764
rect 3936 12724 3942 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 6886 12764 6914 12872
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7892 12804 8033 12832
rect 7892 12792 7898 12804
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14332 12804 14841 12832
rect 14332 12792 14338 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 15286 12792 15292 12844
rect 15344 12792 15350 12844
rect 6696 12736 6914 12764
rect 6696 12724 6702 12736
rect 2556 12668 3464 12696
rect 2556 12656 2562 12668
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 3436 12637 3464 12668
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 7340 12668 7573 12696
rect 7340 12656 7346 12668
rect 7561 12665 7573 12668
rect 7607 12665 7619 12699
rect 7561 12659 7619 12665
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 1912 12600 2145 12628
rect 1912 12588 1918 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2133 12591 2191 12597
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 5626 12628 5632 12640
rect 3467 12600 5632 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 1104 12538 16836 12560
rect 1104 12486 2916 12538
rect 2968 12486 2980 12538
rect 3032 12486 3044 12538
rect 3096 12486 3108 12538
rect 3160 12486 3172 12538
rect 3224 12486 6849 12538
rect 6901 12486 6913 12538
rect 6965 12486 6977 12538
rect 7029 12486 7041 12538
rect 7093 12486 7105 12538
rect 7157 12486 10782 12538
rect 10834 12486 10846 12538
rect 10898 12486 10910 12538
rect 10962 12486 10974 12538
rect 11026 12486 11038 12538
rect 11090 12486 14715 12538
rect 14767 12486 14779 12538
rect 14831 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 16836 12538
rect 1104 12464 16836 12486
rect 6825 12427 6883 12433
rect 6825 12393 6837 12427
rect 6871 12424 6883 12427
rect 6914 12424 6920 12436
rect 6871 12396 6920 12424
rect 6871 12393 6883 12396
rect 6825 12387 6883 12393
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 7190 12424 7196 12436
rect 6972 12396 7196 12424
rect 6972 12384 6978 12396
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 4154 12316 4160 12368
rect 4212 12316 4218 12368
rect 1854 12248 1860 12300
rect 1912 12248 1918 12300
rect 6730 12288 6736 12300
rect 4172 12260 6736 12288
rect 1578 12180 1584 12232
rect 1636 12180 1642 12232
rect 2958 12180 2964 12232
rect 3016 12180 3022 12232
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 4172 12229 4200 12260
rect 6730 12248 6736 12260
rect 6788 12288 6794 12300
rect 6788 12260 7604 12288
rect 6788 12248 6794 12260
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 3292 12192 4169 12220
rect 3292 12180 3298 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 4356 12152 4384 12183
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 6052 12192 6101 12220
rect 6052 12180 6058 12192
rect 6089 12189 6101 12192
rect 6135 12220 6147 12223
rect 6638 12220 6644 12232
rect 6135 12192 6644 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 7190 12220 7196 12232
rect 6963 12192 7196 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7576 12229 7604 12260
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 4120 12124 4384 12152
rect 7484 12152 7512 12183
rect 8478 12152 8484 12164
rect 7484 12124 8484 12152
rect 4120 12112 4126 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 3329 12087 3387 12093
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3970 12084 3976 12096
rect 3375 12056 3976 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3970 12044 3976 12056
rect 4028 12084 4034 12096
rect 5534 12084 5540 12096
rect 4028 12056 5540 12084
rect 4028 12044 4034 12056
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 6546 12084 6552 12096
rect 6227 12056 6552 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7466 12044 7472 12096
rect 7524 12044 7530 12096
rect 1104 11994 16995 12016
rect 1104 11942 4882 11994
rect 4934 11942 4946 11994
rect 4998 11942 5010 11994
rect 5062 11942 5074 11994
rect 5126 11942 5138 11994
rect 5190 11942 8815 11994
rect 8867 11942 8879 11994
rect 8931 11942 8943 11994
rect 8995 11942 9007 11994
rect 9059 11942 9071 11994
rect 9123 11942 12748 11994
rect 12800 11942 12812 11994
rect 12864 11942 12876 11994
rect 12928 11942 12940 11994
rect 12992 11942 13004 11994
rect 13056 11942 16681 11994
rect 16733 11942 16745 11994
rect 16797 11942 16809 11994
rect 16861 11942 16873 11994
rect 16925 11942 16937 11994
rect 16989 11942 16995 11994
rect 1104 11920 16995 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 1636 11852 2421 11880
rect 1636 11840 1642 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 6788 11852 8156 11880
rect 6788 11840 6794 11852
rect 2958 11772 2964 11824
rect 3016 11772 3022 11824
rect 6825 11815 6883 11821
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 6914 11812 6920 11824
rect 6871 11784 6920 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 7466 11772 7472 11824
rect 7524 11772 7530 11824
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 3142 11704 3148 11756
rect 3200 11704 3206 11756
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 4062 11744 4068 11756
rect 3384 11716 4068 11744
rect 3384 11704 3390 11716
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 6012 11676 6040 11707
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 8128 11744 8156 11852
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 8536 11784 9168 11812
rect 8536 11772 8542 11784
rect 9140 11753 9168 11784
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8128 11716 8953 11744
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10873 11747 10931 11753
rect 10873 11744 10885 11747
rect 10192 11716 10885 11744
rect 10192 11704 10198 11716
rect 10873 11713 10885 11716
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 14332 11716 14841 11744
rect 14332 11704 14338 11716
rect 14829 11713 14841 11716
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 16025 11747 16083 11753
rect 16025 11744 16037 11747
rect 15436 11716 16037 11744
rect 15436 11704 15442 11716
rect 16025 11713 16037 11716
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 7282 11676 7288 11688
rect 6012 11648 7288 11676
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 8938 11568 8944 11620
rect 8996 11568 9002 11620
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12437 11611 12495 11617
rect 12437 11608 12449 11611
rect 12216 11580 12449 11608
rect 12216 11568 12222 11580
rect 12437 11577 12449 11580
rect 12483 11577 12495 11611
rect 12437 11571 12495 11577
rect 5905 11543 5963 11549
rect 5905 11509 5917 11543
rect 5951 11540 5963 11543
rect 6546 11540 6552 11552
rect 5951 11512 6552 11540
rect 5951 11509 5963 11512
rect 5905 11503 5963 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 8297 11543 8355 11549
rect 8297 11540 8309 11543
rect 7248 11512 8309 11540
rect 7248 11500 7254 11512
rect 8297 11509 8309 11512
rect 8343 11509 8355 11543
rect 8297 11503 8355 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10652 11512 10793 11540
rect 10652 11500 10658 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11388 11512 11805 11540
rect 11388 11500 11394 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 14921 11543 14979 11549
rect 14921 11509 14933 11543
rect 14967 11540 14979 11543
rect 16022 11540 16028 11552
rect 14967 11512 16028 11540
rect 14967 11509 14979 11512
rect 14921 11503 14979 11509
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16114 11500 16120 11552
rect 16172 11500 16178 11552
rect 1104 11450 16836 11472
rect 1104 11398 2916 11450
rect 2968 11398 2980 11450
rect 3032 11398 3044 11450
rect 3096 11398 3108 11450
rect 3160 11398 3172 11450
rect 3224 11398 6849 11450
rect 6901 11398 6913 11450
rect 6965 11398 6977 11450
rect 7029 11398 7041 11450
rect 7093 11398 7105 11450
rect 7157 11398 10782 11450
rect 10834 11398 10846 11450
rect 10898 11398 10910 11450
rect 10962 11398 10974 11450
rect 11026 11398 11038 11450
rect 11090 11398 14715 11450
rect 14767 11398 14779 11450
rect 14831 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 16836 11450
rect 1104 11376 16836 11398
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7340 11308 7696 11336
rect 7340 11296 7346 11308
rect 7668 11280 7696 11308
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10192 11308 11836 11336
rect 10192 11296 10198 11308
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 8021 11271 8079 11277
rect 8021 11268 8033 11271
rect 7708 11240 8033 11268
rect 7708 11228 7714 11240
rect 8021 11237 8033 11240
rect 8067 11237 8079 11271
rect 8021 11231 8079 11237
rect 6546 11160 6552 11212
rect 6604 11160 6610 11212
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 11808 11209 11836 11308
rect 9769 11203 9827 11209
rect 9769 11200 9781 11203
rect 7800 11172 9781 11200
rect 7800 11160 7806 11172
rect 9769 11169 9781 11172
rect 9815 11200 9827 11203
rect 11793 11203 11851 11209
rect 9815 11172 11284 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 8938 11132 8944 11144
rect 7682 11104 8944 11132
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 11256 11132 11284 11172
rect 11793 11169 11805 11203
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 15470 11200 15476 11212
rect 11940 11172 15476 11200
rect 11940 11160 11946 11172
rect 12434 11132 12440 11144
rect 11256 11104 12440 11132
rect 12434 11092 12440 11104
rect 12492 11132 12498 11144
rect 12618 11132 12624 11144
rect 12492 11104 12624 11132
rect 12492 11092 12498 11104
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13648 11141 13676 11172
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16022 11160 16028 11212
rect 16080 11160 16086 11212
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11101 13691 11135
rect 13633 11095 13691 11101
rect 14274 11092 14280 11144
rect 14332 11092 14338 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 10042 11024 10048 11076
rect 10100 11024 10106 11076
rect 11330 11064 11336 11076
rect 11270 11036 11336 11064
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 13538 11024 13544 11076
rect 13596 11024 13602 11076
rect 15286 11024 15292 11076
rect 15344 11024 15350 11076
rect 15746 11024 15752 11076
rect 15804 11064 15810 11076
rect 16316 11064 16344 11095
rect 15804 11036 16344 11064
rect 15804 11024 15810 11036
rect 1104 10906 16995 10928
rect 1104 10854 4882 10906
rect 4934 10854 4946 10906
rect 4998 10854 5010 10906
rect 5062 10854 5074 10906
rect 5126 10854 5138 10906
rect 5190 10854 8815 10906
rect 8867 10854 8879 10906
rect 8931 10854 8943 10906
rect 8995 10854 9007 10906
rect 9059 10854 9071 10906
rect 9123 10854 12748 10906
rect 12800 10854 12812 10906
rect 12864 10854 12876 10906
rect 12928 10854 12940 10906
rect 12992 10854 13004 10906
rect 13056 10854 16681 10906
rect 16733 10854 16745 10906
rect 16797 10854 16809 10906
rect 16861 10854 16873 10906
rect 16925 10854 16937 10906
rect 16989 10854 16995 10906
rect 1104 10832 16995 10854
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6641 10795 6699 10801
rect 6641 10792 6653 10795
rect 6328 10764 6653 10792
rect 6328 10752 6334 10764
rect 6641 10761 6653 10764
rect 6687 10761 6699 10795
rect 6641 10755 6699 10761
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 7742 10792 7748 10804
rect 7699 10764 7748 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 15286 10752 15292 10804
rect 15344 10752 15350 10804
rect 11149 10727 11207 10733
rect 11149 10693 11161 10727
rect 11195 10724 11207 10727
rect 11882 10724 11888 10736
rect 11195 10696 11888 10724
rect 11195 10693 11207 10696
rect 11149 10687 11207 10693
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 13538 10684 13544 10736
rect 13596 10684 13602 10736
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 5868 10628 6745 10656
rect 5868 10616 5874 10628
rect 6733 10625 6745 10628
rect 6779 10656 6791 10659
rect 7190 10656 7196 10668
rect 6779 10628 7196 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9306 10656 9312 10668
rect 8987 10628 9312 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9766 10656 9772 10668
rect 9447 10628 9772 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 15470 10656 15476 10668
rect 15427 10628 15476 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10588 12587 10591
rect 13262 10588 13268 10600
rect 12575 10560 13268 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 12268 10452 12296 10551
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13538 10548 13544 10600
rect 13596 10588 13602 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 13596 10560 14289 10588
rect 13596 10548 13602 10560
rect 14277 10557 14289 10560
rect 14323 10588 14335 10591
rect 15856 10588 15884 10619
rect 14323 10560 15884 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 12526 10452 12532 10464
rect 12268 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 15933 10455 15991 10461
rect 15933 10421 15945 10455
rect 15979 10452 15991 10455
rect 16298 10452 16304 10464
rect 15979 10424 16304 10452
rect 15979 10421 15991 10424
rect 15933 10415 15991 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 1104 10362 16836 10384
rect 1104 10310 2916 10362
rect 2968 10310 2980 10362
rect 3032 10310 3044 10362
rect 3096 10310 3108 10362
rect 3160 10310 3172 10362
rect 3224 10310 6849 10362
rect 6901 10310 6913 10362
rect 6965 10310 6977 10362
rect 7029 10310 7041 10362
rect 7093 10310 7105 10362
rect 7157 10310 10782 10362
rect 10834 10310 10846 10362
rect 10898 10310 10910 10362
rect 10962 10310 10974 10362
rect 11026 10310 11038 10362
rect 11090 10310 14715 10362
rect 14767 10310 14779 10362
rect 14831 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 16836 10362
rect 1104 10288 16836 10310
rect 10042 10208 10048 10260
rect 10100 10208 10106 10260
rect 13262 10208 13268 10260
rect 13320 10208 13326 10260
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 3252 10084 5273 10112
rect 3252 10056 3280 10084
rect 5261 10081 5273 10084
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 10594 10072 10600 10124
rect 10652 10072 10658 10124
rect 10873 10115 10931 10121
rect 10873 10081 10885 10115
rect 10919 10112 10931 10115
rect 12158 10112 12164 10124
rect 10919 10084 12164 10112
rect 10919 10081 10931 10084
rect 10873 10075 10931 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12492 10084 12633 10112
rect 12492 10072 12498 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 15378 10112 15384 10124
rect 14323 10084 15384 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 3234 10004 3240 10056
rect 3292 10004 3298 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 4157 10047 4215 10053
rect 3467 10016 4108 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3970 9936 3976 9988
rect 4028 9936 4034 9988
rect 2501 9911 2559 9917
rect 2501 9877 2513 9911
rect 2547 9908 2559 9911
rect 2682 9908 2688 9920
rect 2547 9880 2688 9908
rect 2547 9877 2559 9880
rect 2501 9871 2559 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 3292 9880 3341 9908
rect 3292 9868 3298 9880
rect 3329 9877 3341 9880
rect 3375 9877 3387 9911
rect 4080 9908 4108 10016
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4172 9976 4200 10007
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 9214 10044 9220 10056
rect 8435 10016 9220 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 9539 10016 10088 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 4522 9976 4528 9988
rect 4172 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 9766 9976 9772 9988
rect 7055 9948 9772 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10060 9976 10088 10016
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 13538 10044 13544 10056
rect 13403 10016 13544 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 10060 9948 10180 9976
rect 4338 9908 4344 9920
rect 4080 9880 4344 9908
rect 3329 9871 3387 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 8478 9868 8484 9920
rect 8536 9868 8542 9920
rect 9401 9911 9459 9917
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9858 9908 9864 9920
rect 9447 9880 9864 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10152 9908 10180 9948
rect 11882 9936 11888 9988
rect 11940 9936 11946 9988
rect 15562 9936 15568 9988
rect 15620 9936 15626 9988
rect 16025 9979 16083 9985
rect 16025 9945 16037 9979
rect 16071 9976 16083 9979
rect 16114 9976 16120 9988
rect 16071 9948 16120 9976
rect 16071 9945 16083 9948
rect 16025 9939 16083 9945
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 11698 9908 11704 9920
rect 10152 9880 11704 9908
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 1104 9818 16995 9840
rect 1104 9766 4882 9818
rect 4934 9766 4946 9818
rect 4998 9766 5010 9818
rect 5062 9766 5074 9818
rect 5126 9766 5138 9818
rect 5190 9766 8815 9818
rect 8867 9766 8879 9818
rect 8931 9766 8943 9818
rect 8995 9766 9007 9818
rect 9059 9766 9071 9818
rect 9123 9766 12748 9818
rect 12800 9766 12812 9818
rect 12864 9766 12876 9818
rect 12928 9766 12940 9818
rect 12992 9766 13004 9818
rect 13056 9766 16681 9818
rect 16733 9766 16745 9818
rect 16797 9766 16809 9818
rect 16861 9766 16873 9818
rect 16925 9766 16937 9818
rect 16989 9766 16995 9818
rect 1104 9744 16995 9766
rect 2406 9596 2412 9648
rect 2464 9596 2470 9648
rect 2682 9596 2688 9648
rect 2740 9596 2746 9648
rect 3970 9636 3976 9648
rect 3910 9608 3976 9636
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 6840 9608 7604 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2424 9568 2452 9596
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 1995 9540 2452 9568
rect 4172 9540 4813 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 3326 9500 3332 9512
rect 2455 9472 3332 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1636 9336 1869 9364
rect 1636 9324 1642 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 4172 9373 4200 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5000 9500 5028 9531
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6840 9577 6868 9608
rect 7576 9580 7604 9608
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 8536 9608 8861 9636
rect 8536 9596 8542 9608
rect 8849 9605 8861 9608
rect 8895 9605 8907 9639
rect 8849 9599 8907 9605
rect 9858 9596 9864 9648
rect 9916 9596 9922 9648
rect 11882 9596 11888 9648
rect 11940 9596 11946 9648
rect 12526 9596 12532 9648
rect 12584 9596 12590 9648
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 15620 9608 16129 9636
rect 15620 9596 15626 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5776 9540 6009 9568
rect 5776 9528 5782 9540
rect 5997 9537 6009 9540
rect 6043 9568 6055 9571
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6043 9540 6837 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 7035 9571 7093 9577
rect 7035 9537 7047 9571
rect 7081 9568 7093 9571
rect 7374 9568 7380 9580
rect 7081 9540 7380 9568
rect 7081 9537 7093 9540
rect 7035 9531 7093 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7616 9540 7941 9568
rect 7616 9528 7622 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11756 9540 11989 9568
rect 11756 9528 11762 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12434 9528 12440 9580
rect 12492 9528 12498 9580
rect 15378 9528 15384 9580
rect 15436 9528 15442 9580
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15528 9540 16037 9568
rect 15528 9528 15534 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 5166 9500 5172 9512
rect 5000 9472 5172 9500
rect 5166 9460 5172 9472
rect 5224 9500 5230 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5224 9472 5825 9500
rect 5224 9460 5230 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7834 9500 7840 9512
rect 7239 9472 7840 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 5828 9432 5856 9463
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 8067 9472 8585 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 9214 9500 9220 9512
rect 8573 9463 8631 9469
rect 8680 9472 9220 9500
rect 6086 9432 6092 9444
rect 5828 9404 6092 9432
rect 6086 9392 6092 9404
rect 6144 9432 6150 9444
rect 6144 9404 6868 9432
rect 6144 9392 6150 9404
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 2464 9336 4169 9364
rect 2464 9324 2470 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4157 9327 4215 9333
rect 4890 9324 4896 9376
rect 4948 9324 4954 9376
rect 5902 9324 5908 9376
rect 5960 9324 5966 9376
rect 6840 9373 6868 9404
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 8386 9364 8392 9376
rect 6871 9336 8392 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 8386 9324 8392 9336
rect 8444 9364 8450 9376
rect 8680 9364 8708 9472
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 9272 9472 10333 9500
rect 9272 9460 9278 9472
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 15473 9435 15531 9441
rect 15473 9401 15485 9435
rect 15519 9432 15531 9435
rect 15746 9432 15752 9444
rect 15519 9404 15752 9432
rect 15519 9401 15531 9404
rect 15473 9395 15531 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 8444 9336 8708 9364
rect 8444 9324 8450 9336
rect 1104 9274 16836 9296
rect 1104 9222 2916 9274
rect 2968 9222 2980 9274
rect 3032 9222 3044 9274
rect 3096 9222 3108 9274
rect 3160 9222 3172 9274
rect 3224 9222 6849 9274
rect 6901 9222 6913 9274
rect 6965 9222 6977 9274
rect 7029 9222 7041 9274
rect 7093 9222 7105 9274
rect 7157 9222 10782 9274
rect 10834 9222 10846 9274
rect 10898 9222 10910 9274
rect 10962 9222 10974 9274
rect 11026 9222 11038 9274
rect 11090 9222 14715 9274
rect 14767 9222 14779 9274
rect 14831 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 16836 9274
rect 1104 9200 16836 9222
rect 1578 8984 1584 9036
rect 1636 8984 1642 9036
rect 5626 8984 5632 9036
rect 5684 8984 5690 9036
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 5960 8996 7052 9024
rect 5960 8984 5966 8996
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 7024 8965 7052 8996
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 4948 8928 6653 8956
rect 4948 8916 4954 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7524 8928 7757 8956
rect 7524 8916 7530 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 12250 8956 12256 8968
rect 11103 8928 12256 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 1854 8848 1860 8900
rect 1912 8848 1918 8900
rect 3234 8888 3240 8900
rect 3082 8860 3240 8888
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 5077 8891 5135 8897
rect 5077 8857 5089 8891
rect 5123 8857 5135 8891
rect 5077 8851 5135 8857
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 2648 8792 3341 8820
rect 2648 8780 2654 8792
rect 3329 8789 3341 8792
rect 3375 8820 3387 8823
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 3375 8792 4813 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 5092 8820 5120 8851
rect 5166 8848 5172 8900
rect 5224 8848 5230 8900
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 5905 8891 5963 8897
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 5994 8888 6000 8900
rect 5951 8860 6000 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 8021 8891 8079 8897
rect 8021 8857 8033 8891
rect 8067 8857 8079 8891
rect 8021 8851 8079 8857
rect 5442 8820 5448 8832
rect 5092 8792 5448 8820
rect 4801 8783 4859 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5684 8792 6101 8820
rect 5684 8780 5690 8792
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 6089 8783 6147 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 8036 8820 8064 8851
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 14476 8888 14504 8919
rect 15378 8888 15384 8900
rect 11756 8860 15384 8888
rect 11756 8848 11762 8860
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 7432 8792 8064 8820
rect 7432 8780 7438 8792
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10410 8820 10416 8832
rect 9824 8792 10416 8820
rect 9824 8780 9830 8792
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 14366 8780 14372 8832
rect 14424 8780 14430 8832
rect 1104 8730 16995 8752
rect 1104 8678 4882 8730
rect 4934 8678 4946 8730
rect 4998 8678 5010 8730
rect 5062 8678 5074 8730
rect 5126 8678 5138 8730
rect 5190 8678 8815 8730
rect 8867 8678 8879 8730
rect 8931 8678 8943 8730
rect 8995 8678 9007 8730
rect 9059 8678 9071 8730
rect 9123 8678 12748 8730
rect 12800 8678 12812 8730
rect 12864 8678 12876 8730
rect 12928 8678 12940 8730
rect 12992 8678 13004 8730
rect 13056 8678 16681 8730
rect 16733 8678 16745 8730
rect 16797 8678 16809 8730
rect 16861 8678 16873 8730
rect 16925 8678 16937 8730
rect 16989 8678 16995 8730
rect 1104 8656 16995 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 1912 8588 2513 8616
rect 1912 8576 1918 8588
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 2501 8579 2559 8585
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 9364 8588 10241 8616
rect 9364 8576 9370 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 7558 8508 7564 8560
rect 7616 8548 7622 8560
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 7616 8520 7665 8548
rect 7616 8508 7622 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8352 8520 8953 8548
rect 8352 8508 8358 8520
rect 8941 8517 8953 8520
rect 8987 8517 8999 8551
rect 14366 8548 14372 8560
rect 14122 8520 14372 8548
rect 8941 8511 8999 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 2590 8440 2596 8492
rect 2648 8440 2654 8492
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 8202 8480 8208 8492
rect 5500 8452 8208 8480
rect 5500 8440 5506 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14660 8452 15117 8480
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14660 8421 14688 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14608 8384 14657 8412
rect 14608 8372 14614 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 7926 8304 7932 8356
rect 7984 8344 7990 8356
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7984 8316 8033 8344
rect 7984 8304 7990 8316
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8386 8344 8392 8356
rect 8021 8307 8079 8313
rect 8128 8316 8392 8344
rect 7653 8279 7711 8285
rect 7653 8245 7665 8279
rect 7699 8276 7711 8279
rect 8128 8276 8156 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 7699 8248 8156 8276
rect 15197 8279 15255 8285
rect 7699 8245 7711 8248
rect 7653 8239 7711 8245
rect 15197 8245 15209 8279
rect 15243 8276 15255 8279
rect 16298 8276 16304 8288
rect 15243 8248 16304 8276
rect 15243 8245 15255 8248
rect 15197 8239 15255 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 1104 8186 16836 8208
rect 1104 8134 2916 8186
rect 2968 8134 2980 8186
rect 3032 8134 3044 8186
rect 3096 8134 3108 8186
rect 3160 8134 3172 8186
rect 3224 8134 6849 8186
rect 6901 8134 6913 8186
rect 6965 8134 6977 8186
rect 7029 8134 7041 8186
rect 7093 8134 7105 8186
rect 7157 8134 10782 8186
rect 10834 8134 10846 8186
rect 10898 8134 10910 8186
rect 10962 8134 10974 8186
rect 11026 8134 11038 8186
rect 11090 8134 14715 8186
rect 14767 8134 14779 8186
rect 14831 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 16836 8186
rect 1104 8112 16836 8134
rect 8294 8072 8300 8084
rect 4172 8044 8300 8072
rect 4172 7877 4200 8044
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 12952 8044 13645 8072
rect 12952 8032 12958 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 7973 5779 8007
rect 5721 7967 5779 7973
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 5736 7936 5764 7967
rect 9490 7936 9496 7948
rect 4580 7908 9496 7936
rect 4580 7896 4586 7908
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 9324 7877 9352 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8260 7840 8401 7868
rect 8260 7828 8266 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9398 7828 9404 7880
rect 9456 7828 9462 7880
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 14550 7868 14556 7880
rect 13771 7840 14556 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 10428 7800 10456 7828
rect 7055 7772 10456 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 14274 7760 14280 7812
rect 14332 7760 14338 7812
rect 15286 7760 15292 7812
rect 15344 7760 15350 7812
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 15988 7772 16037 7800
rect 15988 7760 15994 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3660 7704 4077 7732
rect 3660 7692 3666 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 8386 7732 8392 7744
rect 7883 7704 8392 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 1104 7642 16995 7664
rect 1104 7590 4882 7642
rect 4934 7590 4946 7642
rect 4998 7590 5010 7642
rect 5062 7590 5074 7642
rect 5126 7590 5138 7642
rect 5190 7590 8815 7642
rect 8867 7590 8879 7642
rect 8931 7590 8943 7642
rect 8995 7590 9007 7642
rect 9059 7590 9071 7642
rect 9123 7590 12748 7642
rect 12800 7590 12812 7642
rect 12864 7590 12876 7642
rect 12928 7590 12940 7642
rect 12992 7590 13004 7642
rect 13056 7590 16681 7642
rect 16733 7590 16745 7642
rect 16797 7590 16809 7642
rect 16861 7590 16873 7642
rect 16925 7590 16937 7642
rect 16989 7590 16995 7642
rect 1104 7568 16995 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2832 7500 2973 7528
rect 2832 7488 2838 7500
rect 2961 7497 2973 7500
rect 3007 7497 3019 7531
rect 2961 7491 3019 7497
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8536 7500 9352 7528
rect 8536 7488 8542 7500
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 2869 7463 2927 7469
rect 2869 7460 2881 7463
rect 2740 7432 2881 7460
rect 2740 7420 2746 7432
rect 2869 7429 2881 7432
rect 2915 7429 2927 7463
rect 9214 7460 9220 7472
rect 8234 7432 9220 7460
rect 2869 7423 2927 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 9324 7469 9352 7500
rect 15286 7488 15292 7540
rect 15344 7488 15350 7540
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7429 9367 7463
rect 9309 7423 9367 7429
rect 10318 7420 10324 7472
rect 10376 7420 10382 7472
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 14332 7432 15884 7460
rect 14332 7420 14338 7432
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2590 7392 2596 7404
rect 2179 7364 2596 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2590 7352 2596 7364
rect 2648 7392 2654 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2648 7364 2789 7392
rect 2648 7352 2654 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5718 7392 5724 7404
rect 5592 7364 5724 7392
rect 5592 7352 5598 7364
rect 5718 7352 5724 7364
rect 5776 7392 5782 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5776 7364 5825 7392
rect 5776 7352 5782 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6086 7392 6092 7404
rect 6043 7364 6092 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8444 7364 9045 7392
rect 8444 7352 8450 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 14384 7401 14412 7432
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11204 7364 11713 7392
rect 11204 7352 11210 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15856 7401 15884 7432
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3191 7296 3893 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 6733 7327 6791 7333
rect 6733 7324 6745 7327
rect 3881 7287 3939 7293
rect 5000 7296 6745 7324
rect 2498 7216 2504 7268
rect 2556 7256 2562 7268
rect 2593 7259 2651 7265
rect 2593 7256 2605 7259
rect 2556 7228 2605 7256
rect 2556 7216 2562 7228
rect 2593 7225 2605 7228
rect 2639 7225 2651 7259
rect 2593 7219 2651 7225
rect 2038 7148 2044 7200
rect 2096 7148 2102 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 5000 7197 5028 7296
rect 6733 7293 6745 7296
rect 6779 7293 6791 7327
rect 6733 7287 6791 7293
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 8202 7324 8208 7336
rect 7055 7296 8208 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8018 7216 8024 7268
rect 8076 7256 8082 7268
rect 8481 7259 8539 7265
rect 8481 7256 8493 7259
rect 8076 7228 8493 7256
rect 8076 7216 8082 7228
rect 8481 7225 8493 7228
rect 8527 7225 8539 7259
rect 8481 7219 8539 7225
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4396 7160 4997 7188
rect 4396 7148 4402 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 5997 7191 6055 7197
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 7190 7188 7196 7200
rect 6043 7160 7196 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 10781 7191 10839 7197
rect 10781 7188 10793 7191
rect 8168 7160 10793 7188
rect 8168 7148 8174 7160
rect 10781 7157 10793 7160
rect 10827 7157 10839 7191
rect 10781 7151 10839 7157
rect 11790 7148 11796 7200
rect 11848 7148 11854 7200
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 1104 7098 16836 7120
rect 1104 7046 2916 7098
rect 2968 7046 2980 7098
rect 3032 7046 3044 7098
rect 3096 7046 3108 7098
rect 3160 7046 3172 7098
rect 3224 7046 6849 7098
rect 6901 7046 6913 7098
rect 6965 7046 6977 7098
rect 7029 7046 7041 7098
rect 7093 7046 7105 7098
rect 7157 7046 10782 7098
rect 10834 7046 10846 7098
rect 10898 7046 10910 7098
rect 10962 7046 10974 7098
rect 11026 7046 11038 7098
rect 11090 7046 14715 7098
rect 14767 7046 14779 7098
rect 14831 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 16836 7098
rect 1104 7024 16836 7046
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 12357 6987 12415 6993
rect 12357 6984 12369 6987
rect 11848 6956 12369 6984
rect 11848 6944 11854 6956
rect 12357 6953 12369 6956
rect 12403 6953 12415 6987
rect 12357 6947 12415 6953
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2774 6848 2780 6860
rect 2547 6820 2780 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 4522 6848 4528 6860
rect 3252 6820 4528 6848
rect 2590 6740 2596 6792
rect 2648 6740 2654 6792
rect 3252 6789 3280 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 6086 6848 6092 6860
rect 5842 6820 6092 6848
rect 6086 6808 6092 6820
rect 6144 6848 6150 6860
rect 10229 6851 10287 6857
rect 6144 6820 7328 6848
rect 6144 6808 6150 6820
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 4338 6780 4344 6792
rect 3384 6752 4344 6780
rect 3384 6740 3390 6752
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 6638 6780 6644 6792
rect 5123 6752 6644 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6912 6783 6970 6789
rect 6912 6749 6924 6783
rect 6958 6780 6970 6783
rect 7190 6780 7196 6792
rect 6958 6752 7196 6780
rect 6958 6749 6970 6752
rect 6912 6743 6970 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7300 6789 7328 6820
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10318 6848 10324 6860
rect 10275 6820 10324 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 11146 6848 11152 6860
rect 10919 6820 11152 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 14274 6808 14280 6860
rect 14332 6808 14338 6860
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 8076 6752 8217 6780
rect 8076 6740 8082 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9456 6752 9873 6780
rect 9456 6740 9462 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 4801 6715 4859 6721
rect 4801 6712 4813 6715
rect 4764 6684 4813 6712
rect 4764 6672 4770 6684
rect 4801 6681 4813 6684
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 5169 6715 5227 6721
rect 5169 6681 5181 6715
rect 5215 6712 5227 6715
rect 5442 6712 5448 6724
rect 5215 6684 5448 6712
rect 5215 6681 5227 6684
rect 5169 6675 5227 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 7009 6715 7067 6721
rect 5644 6684 6224 6712
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5644 6644 5672 6684
rect 5316 6616 5672 6644
rect 5316 6604 5322 6616
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5868 6616 5917 6644
rect 5868 6604 5874 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 6086 6604 6092 6656
rect 6144 6604 6150 6656
rect 6196 6644 6224 6684
rect 7009 6681 7021 6715
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 6716 6647 6774 6653
rect 6716 6644 6728 6647
rect 6196 6616 6728 6644
rect 6716 6613 6728 6616
rect 6762 6613 6774 6647
rect 7024 6644 7052 6675
rect 7098 6672 7104 6724
rect 7156 6672 7162 6724
rect 11790 6672 11796 6724
rect 11848 6672 11854 6724
rect 14550 6672 14556 6724
rect 14608 6672 14614 6724
rect 15838 6712 15844 6724
rect 15778 6684 15844 6712
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 7650 6644 7656 6656
rect 7024 6616 7656 6644
rect 6716 6607 6774 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8202 6644 8208 6656
rect 8159 6616 8208 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13136 6616 13277 6644
rect 13136 6604 13142 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 14366 6604 14372 6656
rect 14424 6644 14430 6656
rect 16025 6647 16083 6653
rect 16025 6644 16037 6647
rect 14424 6616 16037 6644
rect 14424 6604 14430 6616
rect 16025 6613 16037 6616
rect 16071 6613 16083 6647
rect 16025 6607 16083 6613
rect 1104 6554 16995 6576
rect 1104 6502 4882 6554
rect 4934 6502 4946 6554
rect 4998 6502 5010 6554
rect 5062 6502 5074 6554
rect 5126 6502 5138 6554
rect 5190 6502 8815 6554
rect 8867 6502 8879 6554
rect 8931 6502 8943 6554
rect 8995 6502 9007 6554
rect 9059 6502 9071 6554
rect 9123 6502 12748 6554
rect 12800 6502 12812 6554
rect 12864 6502 12876 6554
rect 12928 6502 12940 6554
rect 12992 6502 13004 6554
rect 13056 6502 16681 6554
rect 16733 6502 16745 6554
rect 16797 6502 16809 6554
rect 16861 6502 16873 6554
rect 16925 6502 16937 6554
rect 16989 6502 16995 6554
rect 1104 6480 16995 6502
rect 2590 6440 2596 6452
rect 1780 6412 2596 6440
rect 1780 6313 1808 6412
rect 2590 6400 2596 6412
rect 2648 6440 2654 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 2648 6412 3985 6440
rect 2648 6400 2654 6412
rect 3973 6409 3985 6412
rect 4019 6440 4031 6443
rect 5534 6440 5540 6452
rect 4019 6412 5540 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 7098 6440 7104 6452
rect 6595 6412 7104 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 12618 6440 12624 6452
rect 12483 6412 12624 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2774 6372 2780 6384
rect 2547 6344 2780 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 3142 6332 3148 6384
rect 3200 6332 3206 6384
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9585 6375 9643 6381
rect 9585 6372 9597 6375
rect 9364 6344 9597 6372
rect 9364 6332 9370 6344
rect 9585 6341 9597 6344
rect 9631 6341 9643 6375
rect 9585 6335 9643 6341
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 13326 6375 13384 6381
rect 13326 6372 13338 6375
rect 12308 6344 13338 6372
rect 12308 6332 12314 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2096 6276 2237 6304
rect 2096 6264 2102 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 3936 6276 6929 6304
rect 3936 6264 3942 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7282 6304 7288 6316
rect 7055 6276 7288 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 11698 6304 11704 6316
rect 10100 6276 11704 6304
rect 10100 6264 10106 6276
rect 11698 6264 11704 6276
rect 11756 6304 11762 6316
rect 12360 6313 12388 6344
rect 13326 6341 13338 6344
rect 13372 6372 13384 6375
rect 14366 6372 14372 6384
rect 13372 6344 14372 6372
rect 13372 6341 13384 6344
rect 13326 6335 13384 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 14476 6372 14504 6403
rect 15838 6400 15844 6452
rect 15896 6400 15902 6452
rect 14476 6344 15148 6372
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11756 6276 11897 6304
rect 11756 6264 11762 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12391 6276 12425 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 15120 6313 15148 6344
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14608 6276 14933 6304
rect 14608 6264 14614 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 15749 6307 15807 6313
rect 15749 6304 15761 6307
rect 15436 6276 15761 6304
rect 15436 6264 15442 6276
rect 15749 6273 15761 6276
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 7558 6236 7564 6248
rect 7239 6208 7564 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7558 6196 7564 6208
rect 7616 6236 7622 6248
rect 11146 6236 11152 6248
rect 7616 6208 11152 6236
rect 7616 6196 7622 6208
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 15197 6171 15255 6177
rect 15197 6168 15209 6171
rect 14516 6140 15209 6168
rect 14516 6128 14522 6140
rect 15197 6137 15209 6140
rect 15243 6137 15255 6171
rect 15197 6131 15255 6137
rect 1670 6060 1676 6112
rect 1728 6060 1734 6112
rect 1104 6010 16836 6032
rect 1104 5958 2916 6010
rect 2968 5958 2980 6010
rect 3032 5958 3044 6010
rect 3096 5958 3108 6010
rect 3160 5958 3172 6010
rect 3224 5958 6849 6010
rect 6901 5958 6913 6010
rect 6965 5958 6977 6010
rect 7029 5958 7041 6010
rect 7093 5958 7105 6010
rect 7157 5958 10782 6010
rect 10834 5958 10846 6010
rect 10898 5958 10910 6010
rect 10962 5958 10974 6010
rect 11026 5958 11038 6010
rect 11090 5958 14715 6010
rect 14767 5958 14779 6010
rect 14831 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 16836 6010
rect 1104 5936 16836 5958
rect 14550 5856 14556 5908
rect 14608 5856 14614 5908
rect 4522 5760 4528 5772
rect 3160 5732 4528 5760
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 3160 5701 3188 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 9490 5760 9496 5772
rect 9324 5732 9496 5760
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3326 5652 3332 5704
rect 3384 5652 3390 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 9324 5701 9352 5732
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 12308 5664 14657 5692
rect 12308 5652 12314 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 2516 5624 2544 5652
rect 3878 5624 3884 5636
rect 2516 5596 3884 5624
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 2406 5516 2412 5568
rect 2464 5516 2470 5568
rect 3234 5516 3240 5568
rect 3292 5516 3298 5568
rect 8478 5516 8484 5568
rect 8536 5516 8542 5568
rect 9214 5516 9220 5568
rect 9272 5516 9278 5568
rect 1104 5466 16995 5488
rect 1104 5414 4882 5466
rect 4934 5414 4946 5466
rect 4998 5414 5010 5466
rect 5062 5414 5074 5466
rect 5126 5414 5138 5466
rect 5190 5414 8815 5466
rect 8867 5414 8879 5466
rect 8931 5414 8943 5466
rect 8995 5414 9007 5466
rect 9059 5414 9071 5466
rect 9123 5414 12748 5466
rect 12800 5414 12812 5466
rect 12864 5414 12876 5466
rect 12928 5414 12940 5466
rect 12992 5414 13004 5466
rect 13056 5414 16681 5466
rect 16733 5414 16745 5466
rect 16797 5414 16809 5466
rect 16861 5414 16873 5466
rect 16925 5414 16937 5466
rect 16989 5414 16995 5466
rect 1104 5392 16995 5414
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 8570 5352 8576 5364
rect 6696 5324 8576 5352
rect 6696 5312 6702 5324
rect 8570 5312 8576 5324
rect 8628 5352 8634 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 8628 5324 9965 5352
rect 8628 5312 8634 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2406 5284 2412 5296
rect 2179 5256 2412 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 3878 5244 3884 5296
rect 3936 5244 3942 5296
rect 5534 5284 5540 5296
rect 5000 5256 5540 5284
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1728 5188 1869 5216
rect 1728 5176 1734 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 3234 5176 3240 5228
rect 3292 5176 3298 5228
rect 5000 5225 5028 5256
rect 5534 5244 5540 5256
rect 5592 5284 5598 5296
rect 6086 5284 6092 5296
rect 5592 5256 6092 5284
rect 5592 5244 5598 5256
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 8478 5244 8484 5296
rect 8536 5244 8542 5296
rect 9490 5244 9496 5296
rect 9548 5244 9554 5296
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 4816 5148 4844 5179
rect 5350 5148 5356 5160
rect 4816 5120 5356 5148
rect 5350 5108 5356 5120
rect 5408 5148 5414 5160
rect 5460 5148 5488 5179
rect 5626 5176 5632 5228
rect 5684 5176 5690 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8110 5216 8116 5228
rect 7607 5188 8116 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 7374 5148 7380 5160
rect 5408 5120 7380 5148
rect 5408 5108 5414 5120
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7699 5120 8217 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 4488 5052 5457 5080
rect 4488 5040 4494 5052
rect 5445 5049 5457 5052
rect 5491 5049 5503 5083
rect 5445 5043 5503 5049
rect 4798 4972 4804 5024
rect 4856 4972 4862 5024
rect 1104 4922 16836 4944
rect 1104 4870 2916 4922
rect 2968 4870 2980 4922
rect 3032 4870 3044 4922
rect 3096 4870 3108 4922
rect 3160 4870 3172 4922
rect 3224 4870 6849 4922
rect 6901 4870 6913 4922
rect 6965 4870 6977 4922
rect 7029 4870 7041 4922
rect 7093 4870 7105 4922
rect 7157 4870 10782 4922
rect 10834 4870 10846 4922
rect 10898 4870 10910 4922
rect 10962 4870 10974 4922
rect 11026 4870 11038 4922
rect 11090 4870 14715 4922
rect 14767 4870 14779 4922
rect 14831 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 16836 4922
rect 1104 4848 16836 4870
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 14550 4700 14556 4752
rect 14608 4700 14614 4752
rect 5718 4672 5724 4684
rect 4724 4644 5724 4672
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4724 4613 4752 4644
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4672 4576 4721 4604
rect 4672 4564 4678 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 5460 4613 5488 4644
rect 5718 4632 5724 4644
rect 5776 4672 5782 4684
rect 5994 4672 6000 4684
rect 5776 4644 6000 4672
rect 5776 4632 5782 4644
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 9490 4632 9496 4684
rect 9548 4632 9554 4684
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 14240 4644 14289 4672
rect 14240 4632 14246 4644
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 14277 4635 14335 4641
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 7926 4604 7932 4616
rect 7340 4576 7932 4604
rect 7340 4564 7346 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 8202 4564 8208 4616
rect 8260 4564 8266 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8478 4604 8484 4616
rect 8343 4576 8484 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 10042 4604 10048 4616
rect 9447 4576 10048 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 12342 4604 12348 4616
rect 11931 4576 12348 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13412 4576 13553 4604
rect 13412 4564 13418 4576
rect 13541 4573 13553 4576
rect 13587 4604 13599 4607
rect 15562 4604 15568 4616
rect 13587 4576 15568 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 4522 4496 4528 4548
rect 4580 4496 4586 4548
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4536 4951 4539
rect 5534 4536 5540 4548
rect 4939 4508 5540 4536
rect 4939 4505 4951 4508
rect 4893 4499 4951 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 5718 4536 5724 4548
rect 5675 4508 5724 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 12069 4539 12127 4545
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 13446 4536 13452 4548
rect 12115 4508 13452 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 14366 4496 14372 4548
rect 14424 4536 14430 4548
rect 15856 4536 15884 4567
rect 14424 4508 15884 4536
rect 16117 4539 16175 4545
rect 14424 4496 14430 4508
rect 16117 4505 16129 4539
rect 16163 4536 16175 4539
rect 17034 4536 17040 4548
rect 16163 4508 17040 4536
rect 16163 4505 16175 4508
rect 16117 4499 16175 4505
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 7282 4468 7288 4480
rect 6779 4440 7288 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7374 4428 7380 4480
rect 7432 4428 7438 4480
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 9398 4468 9404 4480
rect 8527 4440 9404 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 11701 4471 11759 4477
rect 11701 4468 11713 4471
rect 11388 4440 11713 4468
rect 11388 4428 11394 4440
rect 11701 4437 11713 4440
rect 11747 4437 11759 4471
rect 11701 4431 11759 4437
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 13906 4468 13912 4480
rect 13679 4440 13912 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4468 14795 4471
rect 15378 4468 15384 4480
rect 14783 4440 15384 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 1104 4378 16995 4400
rect 1104 4326 4882 4378
rect 4934 4326 4946 4378
rect 4998 4326 5010 4378
rect 5062 4326 5074 4378
rect 5126 4326 5138 4378
rect 5190 4326 8815 4378
rect 8867 4326 8879 4378
rect 8931 4326 8943 4378
rect 8995 4326 9007 4378
rect 9059 4326 9071 4378
rect 9123 4326 12748 4378
rect 12800 4326 12812 4378
rect 12864 4326 12876 4378
rect 12928 4326 12940 4378
rect 12992 4326 13004 4378
rect 13056 4326 16681 4378
rect 16733 4326 16745 4378
rect 16797 4326 16809 4378
rect 16861 4326 16873 4378
rect 16925 4326 16937 4378
rect 16989 4326 16995 4378
rect 1104 4304 16995 4326
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 3602 4264 3608 4276
rect 3559 4236 3608 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 4430 4224 4436 4276
rect 4488 4224 4494 4276
rect 4614 4224 4620 4276
rect 4672 4224 4678 4276
rect 5350 4264 5356 4276
rect 5000 4236 5356 4264
rect 4448 4196 4476 4224
rect 2976 4168 4476 4196
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 2976 4128 3004 4168
rect 2915 4100 3004 4128
rect 3053 4131 3111 4137
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3326 4128 3332 4140
rect 3099 4100 3332 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3326 4088 3332 4100
rect 3384 4128 3390 4140
rect 3789 4131 3847 4137
rect 3384 4100 3648 4128
rect 3384 4088 3390 4100
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3620 4060 3648 4100
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 4154 4128 4160 4140
rect 3835 4100 4160 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 3620 4032 4261 4060
rect 3513 4023 3571 4029
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4448 4060 4476 4091
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4672 4100 4721 4128
rect 4672 4088 4678 4100
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 5000 4128 5028 4236
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 14182 4264 14188 4276
rect 13464 4236 14188 4264
rect 5718 4196 5724 4208
rect 5368 4168 5724 4196
rect 5368 4128 5396 4168
rect 5718 4156 5724 4168
rect 5776 4196 5782 4208
rect 6641 4199 6699 4205
rect 6641 4196 6653 4199
rect 5776 4168 6653 4196
rect 5776 4156 5782 4168
rect 6641 4165 6653 4168
rect 6687 4165 6699 4199
rect 6641 4159 6699 4165
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7929 4199 7987 4205
rect 7929 4196 7941 4199
rect 7432 4168 7941 4196
rect 7432 4156 7438 4168
rect 7929 4165 7941 4168
rect 7975 4165 7987 4199
rect 9214 4196 9220 4208
rect 9154 4168 9220 4196
rect 7929 4159 7987 4165
rect 9214 4156 9220 4168
rect 9272 4156 9278 4208
rect 13354 4196 13360 4208
rect 12176 4168 13360 4196
rect 4755 4100 5028 4128
rect 5092 4100 5396 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 5092 4060 5120 4100
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 5592 4100 6561 4128
rect 5592 4088 5598 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7340 4100 7665 4128
rect 7340 4088 7346 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 9640 4100 10977 4128
rect 9640 4088 9646 4100
rect 10965 4097 10977 4100
rect 11011 4128 11023 4131
rect 12176 4128 12204 4168
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 11011 4100 12204 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12400 4100 13001 4128
rect 12400 4088 12406 4100
rect 12989 4097 13001 4100
rect 13035 4128 13047 4131
rect 13464 4128 13492 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 13035 4100 13492 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 14165 4131 14223 4137
rect 14165 4128 14177 4131
rect 14016 4100 14177 4128
rect 4448 4032 5120 4060
rect 5169 4063 5227 4069
rect 4249 4023 4307 4029
rect 5169 4029 5181 4063
rect 5215 4060 5227 4063
rect 5626 4060 5632 4072
rect 5215 4032 5632 4060
rect 5215 4029 5227 4032
rect 5169 4023 5227 4029
rect 3528 3992 3556 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 7984 4032 9689 4060
rect 7984 4020 7990 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 14016 4060 14044 4100
rect 14165 4097 14177 4100
rect 14211 4097 14223 4131
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 14165 4091 14223 4097
rect 15304 4100 15761 4128
rect 13495 4032 14044 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 3697 3995 3755 4001
rect 3528 3964 3648 3992
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3510 3924 3516 3936
rect 3099 3896 3516 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3620 3924 3648 3964
rect 3697 3961 3709 3995
rect 3743 3992 3755 3995
rect 4798 3992 4804 4004
rect 3743 3964 4804 3992
rect 3743 3961 3755 3964
rect 3697 3955 3755 3961
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 12069 3995 12127 4001
rect 5644 3964 7788 3992
rect 4246 3924 4252 3936
rect 3620 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3924 4310 3936
rect 4522 3924 4528 3936
rect 4304 3896 4528 3924
rect 4304 3884 4310 3896
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 5644 3933 5672 3964
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 4764 3896 5273 3924
rect 4764 3884 4770 3896
rect 5261 3893 5273 3896
rect 5307 3893 5319 3927
rect 5261 3887 5319 3893
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3893 5687 3927
rect 7760 3924 7788 3964
rect 12069 3961 12081 3995
rect 12115 3992 12127 3995
rect 12894 3992 12900 4004
rect 12115 3964 12900 3992
rect 12115 3961 12127 3964
rect 12069 3955 12127 3961
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 13357 3995 13415 4001
rect 13357 3961 13369 3995
rect 13403 3961 13415 3995
rect 13357 3955 13415 3961
rect 9766 3924 9772 3936
rect 7760 3896 9772 3924
rect 5629 3887 5687 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 11698 3924 11704 3936
rect 11103 3896 11704 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 11974 3924 11980 3936
rect 11931 3896 11980 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 13372 3924 13400 3955
rect 14274 3924 14280 3936
rect 13372 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15304 3933 15332 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15712 4032 15945 4060
rect 15712 4020 15718 4032
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15160 3896 15301 3924
rect 15160 3884 15166 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 1104 3834 16836 3856
rect 1104 3782 2916 3834
rect 2968 3782 2980 3834
rect 3032 3782 3044 3834
rect 3096 3782 3108 3834
rect 3160 3782 3172 3834
rect 3224 3782 6849 3834
rect 6901 3782 6913 3834
rect 6965 3782 6977 3834
rect 7029 3782 7041 3834
rect 7093 3782 7105 3834
rect 7157 3782 10782 3834
rect 10834 3782 10846 3834
rect 10898 3782 10910 3834
rect 10962 3782 10974 3834
rect 11026 3782 11038 3834
rect 11090 3782 14715 3834
rect 14767 3782 14779 3834
rect 14831 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 16836 3834
rect 1104 3760 16836 3782
rect 3326 3680 3332 3732
rect 3384 3680 3390 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5684 3692 6837 3720
rect 5684 3680 5690 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 9364 3692 10517 3720
rect 9364 3680 9370 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 12894 3680 12900 3732
rect 12952 3680 12958 3732
rect 14277 3723 14335 3729
rect 14277 3689 14289 3723
rect 14323 3720 14335 3723
rect 14366 3720 14372 3732
rect 14323 3692 14372 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 4706 3612 4712 3664
rect 4764 3612 4770 3664
rect 4798 3612 4804 3664
rect 4856 3612 4862 3664
rect 12437 3655 12495 3661
rect 12437 3621 12449 3655
rect 12483 3652 12495 3655
rect 12483 3624 13400 3652
rect 12483 3621 12495 3624
rect 12437 3615 12495 3621
rect 13372 3596 13400 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2038 3584 2044 3596
rect 1995 3556 2044 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 2464 3556 3433 3584
rect 2464 3544 2470 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3568 3556 4936 3584
rect 3568 3544 3574 3556
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3326 3516 3332 3528
rect 3191 3488 3332 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 2332 3448 2360 3479
rect 3326 3476 3332 3488
rect 3384 3516 3390 3528
rect 4908 3525 4936 3556
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 5776 3556 5948 3584
rect 5776 3544 5782 3556
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3384 3488 4629 3516
rect 3384 3476 3390 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 4246 3448 4252 3460
rect 2332 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 4632 3448 4660 3479
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5500 3488 5641 3516
rect 5500 3476 5506 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5644 3448 5672 3479
rect 5810 3476 5816 3528
rect 5868 3476 5874 3528
rect 5920 3525 5948 3556
rect 13354 3544 13360 3596
rect 13412 3544 13418 3596
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3584 13599 3587
rect 14458 3584 14464 3596
rect 13587 3556 14464 3584
rect 13587 3553 13599 3556
rect 13541 3547 13599 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 15703 3556 16221 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 16209 3547 16267 3553
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 5994 3476 6000 3528
rect 6052 3476 6058 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6144 3488 6745 3516
rect 6144 3476 6150 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9214 3516 9220 3528
rect 9171 3488 9220 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 7024 3448 7052 3479
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9398 3525 9404 3528
rect 9392 3516 9404 3525
rect 9359 3488 9404 3516
rect 9392 3479 9404 3488
rect 9398 3476 9404 3479
rect 9456 3476 9462 3528
rect 11054 3476 11060 3528
rect 11112 3476 11118 3528
rect 11330 3525 11336 3528
rect 11324 3516 11336 3525
rect 11291 3488 11336 3516
rect 11324 3479 11336 3488
rect 11330 3476 11336 3479
rect 11388 3476 11394 3528
rect 15378 3476 15384 3528
rect 15436 3525 15442 3528
rect 15436 3516 15448 3525
rect 15436 3488 15481 3516
rect 15436 3479 15448 3488
rect 15436 3476 15442 3479
rect 15562 3476 15568 3528
rect 15620 3516 15626 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15620 3488 16129 3516
rect 15620 3476 15626 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 4632 3420 7052 3448
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2832 3352 2973 3380
rect 2832 3340 2838 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 5077 3383 5135 3389
rect 5077 3349 5089 3383
rect 5123 3380 5135 3383
rect 5350 3380 5356 3392
rect 5123 3352 5356 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 6270 3340 6276 3392
rect 6328 3340 6334 3392
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 8110 3380 8116 3392
rect 7239 3352 8116 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 13262 3340 13268 3392
rect 13320 3340 13326 3392
rect 1104 3290 16995 3312
rect 1104 3238 4882 3290
rect 4934 3238 4946 3290
rect 4998 3238 5010 3290
rect 5062 3238 5074 3290
rect 5126 3238 5138 3290
rect 5190 3238 8815 3290
rect 8867 3238 8879 3290
rect 8931 3238 8943 3290
rect 8995 3238 9007 3290
rect 9059 3238 9071 3290
rect 9123 3238 12748 3290
rect 12800 3238 12812 3290
rect 12864 3238 12876 3290
rect 12928 3238 12940 3290
rect 12992 3238 13004 3290
rect 13056 3238 16681 3290
rect 16733 3238 16745 3290
rect 16797 3238 16809 3290
rect 16861 3238 16873 3290
rect 16925 3238 16937 3290
rect 16989 3238 16995 3290
rect 1104 3216 16995 3238
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 4764 3148 5089 3176
rect 4764 3136 4770 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 5868 3148 6653 3176
rect 5868 3136 5874 3148
rect 6641 3145 6653 3148
rect 6687 3145 6699 3179
rect 6641 3139 6699 3145
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 9272 3148 9321 3176
rect 9272 3136 9278 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 9309 3139 9367 3145
rect 11054 3136 11060 3188
rect 11112 3136 11118 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13909 3179 13967 3185
rect 13909 3176 13921 3179
rect 13412 3148 13921 3176
rect 13412 3136 13418 3148
rect 13909 3145 13921 3148
rect 13955 3145 13967 3179
rect 13909 3139 13967 3145
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 14332 3148 14749 3176
rect 14332 3136 14338 3148
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 14737 3139 14795 3145
rect 3326 3068 3332 3120
rect 3384 3108 3390 3120
rect 3421 3111 3479 3117
rect 3421 3108 3433 3111
rect 3384 3080 3433 3108
rect 3384 3068 3390 3080
rect 3421 3077 3433 3080
rect 3467 3077 3479 3111
rect 4246 3108 4252 3120
rect 3421 3071 3479 3077
rect 3620 3080 4252 3108
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 3620 3049 3648 3080
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 4430 3068 4436 3120
rect 4488 3068 4494 3120
rect 5445 3111 5503 3117
rect 5445 3077 5457 3111
rect 5491 3108 5503 3111
rect 5994 3108 6000 3120
rect 5491 3080 6000 3108
rect 5491 3077 5503 3080
rect 5445 3071 5503 3077
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 14001 3111 14059 3117
rect 14001 3077 14013 3111
rect 14047 3108 14059 3111
rect 14366 3108 14372 3120
rect 14047 3080 14372 3108
rect 14047 3077 14059 3080
rect 14001 3071 14059 3077
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4154 3040 4160 3052
rect 3835 3012 4160 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4154 3000 4160 3012
rect 4212 3040 4218 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4212 3012 4629 3040
rect 4212 3000 4218 3012
rect 4617 3009 4629 3012
rect 4663 3040 4675 3043
rect 5258 3040 5264 3052
rect 4663 3012 5264 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5718 3040 5724 3052
rect 5583 3012 5724 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 1762 2932 1768 2984
rect 1820 2932 1826 2984
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 2464 2944 4261 2972
rect 2464 2932 2470 2944
rect 4249 2941 4261 2944
rect 4295 2972 4307 2975
rect 6086 2972 6092 2984
rect 4295 2944 6092 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 6748 2904 6776 3003
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 8352 3012 9413 3040
rect 8352 3000 8358 3012
rect 9401 3009 9413 3012
rect 9447 3040 9459 3043
rect 9582 3040 9588 3052
rect 9447 3012 9588 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9582 3000 9588 3012
rect 9640 3040 9646 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 9640 3012 10977 3040
rect 9640 3000 9646 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11974 3049 11980 3052
rect 11968 3040 11980 3049
rect 11935 3012 11980 3040
rect 11968 3003 11980 3012
rect 11974 3000 11980 3003
rect 12032 3000 12038 3052
rect 15102 3000 15108 3052
rect 15160 3000 15166 3052
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 14458 2972 14464 2984
rect 14231 2944 14464 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 15194 2932 15200 2984
rect 15252 2932 15258 2984
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 4672 2876 6776 2904
rect 4672 2864 4678 2876
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 13541 2907 13599 2913
rect 13541 2904 13553 2907
rect 13504 2876 13553 2904
rect 13504 2864 13510 2876
rect 13541 2873 13553 2876
rect 13587 2873 13599 2907
rect 14476 2904 14504 2932
rect 15304 2904 15332 2935
rect 14476 2876 15332 2904
rect 13541 2867 13599 2873
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13262 2836 13268 2848
rect 13127 2808 13268 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13262 2796 13268 2808
rect 13320 2836 13326 2848
rect 15194 2836 15200 2848
rect 13320 2808 15200 2836
rect 13320 2796 13326 2808
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 1104 2746 16836 2768
rect 1104 2694 2916 2746
rect 2968 2694 2980 2746
rect 3032 2694 3044 2746
rect 3096 2694 3108 2746
rect 3160 2694 3172 2746
rect 3224 2694 6849 2746
rect 6901 2694 6913 2746
rect 6965 2694 6977 2746
rect 7029 2694 7041 2746
rect 7093 2694 7105 2746
rect 7157 2694 10782 2746
rect 10834 2694 10846 2746
rect 10898 2694 10910 2746
rect 10962 2694 10974 2746
rect 11026 2694 11038 2746
rect 11090 2694 14715 2746
rect 14767 2694 14779 2746
rect 14831 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 16836 2746
rect 1104 2672 16836 2694
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 14550 2632 14556 2644
rect 14507 2604 14556 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14516 2468 15025 2496
rect 14516 2456 14522 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2832 2400 2881 2428
rect 2832 2388 2838 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3660 2400 3985 2428
rect 3660 2388 3666 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6328 2400 6837 2428
rect 6328 2388 6334 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2428 12219 2431
rect 12342 2428 12348 2440
rect 12207 2400 12348 2428
rect 12207 2397 12219 2400
rect 12161 2391 12219 2397
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13354 2428 13360 2440
rect 13219 2400 13360 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14424 2400 14841 2428
rect 14424 2388 14430 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15102 2428 15108 2440
rect 14967 2400 15108 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15252 2400 15669 2428
rect 15252 2388 15258 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 2372 2332 2605 2360
rect 2372 2320 2378 2332
rect 2593 2329 2605 2332
rect 2639 2329 2651 2363
rect 2593 2323 2651 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 4212 2332 4261 2360
rect 4212 2320 4218 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 5534 2320 5540 2372
rect 5592 2360 5598 2372
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 5592 2332 5641 2360
rect 5592 2320 5598 2332
rect 5629 2329 5641 2332
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 7101 2363 7159 2369
rect 7101 2360 7113 2363
rect 6972 2332 7113 2360
rect 6972 2320 6978 2332
rect 7101 2329 7113 2332
rect 7147 2329 7159 2363
rect 7101 2323 7159 2329
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 8352 2332 8401 2360
rect 8352 2320 8358 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8389 2323 8447 2329
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 10045 2363 10103 2369
rect 10045 2360 10057 2363
rect 9732 2332 10057 2360
rect 9732 2320 9738 2332
rect 10045 2329 10057 2332
rect 10091 2329 10103 2363
rect 10045 2323 10103 2329
rect 11146 2320 11152 2372
rect 11204 2360 11210 2372
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 11204 2332 11897 2360
rect 11204 2320 11210 2332
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 11885 2323 11943 2329
rect 12618 2320 12624 2372
rect 12676 2360 12682 2372
rect 12897 2363 12955 2369
rect 12897 2360 12909 2363
rect 12676 2332 12909 2360
rect 12676 2320 12682 2332
rect 12897 2329 12909 2332
rect 12943 2329 12955 2363
rect 12897 2323 12955 2329
rect 15930 2320 15936 2372
rect 15988 2320 15994 2372
rect 1104 2202 16995 2224
rect 1104 2150 4882 2202
rect 4934 2150 4946 2202
rect 4998 2150 5010 2202
rect 5062 2150 5074 2202
rect 5126 2150 5138 2202
rect 5190 2150 8815 2202
rect 8867 2150 8879 2202
rect 8931 2150 8943 2202
rect 8995 2150 9007 2202
rect 9059 2150 9071 2202
rect 9123 2150 12748 2202
rect 12800 2150 12812 2202
rect 12864 2150 12876 2202
rect 12928 2150 12940 2202
rect 12992 2150 13004 2202
rect 13056 2150 16681 2202
rect 16733 2150 16745 2202
rect 16797 2150 16809 2202
rect 16861 2150 16873 2202
rect 16925 2150 16937 2202
rect 16989 2150 16995 2202
rect 1104 2128 16995 2150
rect 842 892 848 944
rect 900 932 906 944
rect 1762 932 1768 944
rect 900 904 1768 932
rect 900 892 906 904
rect 1762 892 1768 904
rect 1820 892 1826 944
rect 14090 892 14096 944
rect 14148 932 14154 944
rect 15930 932 15936 944
rect 14148 904 15936 932
rect 14148 892 14154 904
rect 15930 892 15936 904
rect 15988 892 15994 944
<< via1 >>
rect 13544 17280 13596 17332
rect 14464 17280 14516 17332
rect 2916 15750 2968 15802
rect 2980 15750 3032 15802
rect 3044 15750 3096 15802
rect 3108 15750 3160 15802
rect 3172 15750 3224 15802
rect 6849 15750 6901 15802
rect 6913 15750 6965 15802
rect 6977 15750 7029 15802
rect 7041 15750 7093 15802
rect 7105 15750 7157 15802
rect 10782 15750 10834 15802
rect 10846 15750 10898 15802
rect 10910 15750 10962 15802
rect 10974 15750 11026 15802
rect 11038 15750 11090 15802
rect 14715 15750 14767 15802
rect 14779 15750 14831 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 6276 15444 6328 15496
rect 10600 15444 10652 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 13820 15376 13872 15428
rect 4804 15308 4856 15360
rect 11980 15308 12032 15360
rect 14096 15308 14148 15360
rect 16028 15308 16080 15360
rect 4882 15206 4934 15258
rect 4946 15206 4998 15258
rect 5010 15206 5062 15258
rect 5074 15206 5126 15258
rect 5138 15206 5190 15258
rect 8815 15206 8867 15258
rect 8879 15206 8931 15258
rect 8943 15206 8995 15258
rect 9007 15206 9059 15258
rect 9071 15206 9123 15258
rect 12748 15206 12800 15258
rect 12812 15206 12864 15258
rect 12876 15206 12928 15258
rect 12940 15206 12992 15258
rect 13004 15206 13056 15258
rect 16681 15206 16733 15258
rect 16745 15206 16797 15258
rect 16809 15206 16861 15258
rect 16873 15206 16925 15258
rect 16937 15206 16989 15258
rect 4344 14968 4396 15020
rect 4804 14968 4856 15020
rect 7380 14968 7432 15020
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 11152 14900 11204 14952
rect 15292 14968 15344 15020
rect 3976 14764 4028 14816
rect 5908 14764 5960 14816
rect 9496 14764 9548 14816
rect 9864 14764 9916 14816
rect 11520 14764 11572 14816
rect 12256 14764 12308 14816
rect 13084 14764 13136 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 14556 14764 14608 14816
rect 15568 14764 15620 14816
rect 2916 14662 2968 14714
rect 2980 14662 3032 14714
rect 3044 14662 3096 14714
rect 3108 14662 3160 14714
rect 3172 14662 3224 14714
rect 6849 14662 6901 14714
rect 6913 14662 6965 14714
rect 6977 14662 7029 14714
rect 7041 14662 7093 14714
rect 7105 14662 7157 14714
rect 10782 14662 10834 14714
rect 10846 14662 10898 14714
rect 10910 14662 10962 14714
rect 10974 14662 11026 14714
rect 11038 14662 11090 14714
rect 14715 14662 14767 14714
rect 14779 14662 14831 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 4436 14560 4488 14612
rect 8300 14560 8352 14612
rect 7380 14535 7432 14544
rect 7380 14501 7389 14535
rect 7389 14501 7423 14535
rect 7423 14501 7432 14535
rect 7380 14492 7432 14501
rect 4068 14424 4120 14476
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 6552 14424 6604 14476
rect 8484 14424 8536 14476
rect 2504 14220 2556 14272
rect 3976 14331 4028 14340
rect 3976 14297 3985 14331
rect 3985 14297 4019 14331
rect 4019 14297 4028 14331
rect 3976 14288 4028 14297
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 11888 14424 11940 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 12256 14467 12308 14476
rect 12256 14433 12265 14467
rect 12265 14433 12299 14467
rect 12299 14433 12308 14467
rect 12256 14424 12308 14433
rect 13820 14424 13872 14476
rect 16028 14467 16080 14476
rect 16028 14433 16037 14467
rect 16037 14433 16071 14467
rect 16071 14433 16080 14467
rect 16028 14424 16080 14433
rect 10600 14356 10652 14408
rect 12532 14356 12584 14408
rect 14648 14356 14700 14408
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 4160 14220 4212 14272
rect 6644 14288 6696 14340
rect 11520 14288 11572 14340
rect 15568 14288 15620 14340
rect 6736 14220 6788 14272
rect 9220 14263 9272 14272
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 4882 14118 4934 14170
rect 4946 14118 4998 14170
rect 5010 14118 5062 14170
rect 5074 14118 5126 14170
rect 5138 14118 5190 14170
rect 8815 14118 8867 14170
rect 8879 14118 8931 14170
rect 8943 14118 8995 14170
rect 9007 14118 9059 14170
rect 9071 14118 9123 14170
rect 12748 14118 12800 14170
rect 12812 14118 12864 14170
rect 12876 14118 12928 14170
rect 12940 14118 12992 14170
rect 13004 14118 13056 14170
rect 16681 14118 16733 14170
rect 16745 14118 16797 14170
rect 16809 14118 16861 14170
rect 16873 14118 16925 14170
rect 16937 14118 16989 14170
rect 5632 14016 5684 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 2504 13991 2556 14000
rect 2504 13957 2513 13991
rect 2513 13957 2547 13991
rect 2547 13957 2556 13991
rect 2504 13948 2556 13957
rect 3976 13948 4028 14000
rect 9220 13948 9272 14000
rect 13360 13991 13412 14000
rect 13360 13957 13369 13991
rect 13369 13957 13403 13991
rect 13403 13957 13412 13991
rect 13360 13948 13412 13957
rect 14372 13948 14424 14000
rect 14648 13948 14700 14000
rect 2228 13855 2280 13864
rect 2228 13821 2237 13855
rect 2237 13821 2271 13855
rect 2271 13821 2280 13855
rect 2228 13812 2280 13821
rect 4160 13812 4212 13864
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 11152 13880 11204 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 15476 13880 15528 13932
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 14096 13812 14148 13864
rect 7840 13676 7892 13728
rect 10140 13676 10192 13728
rect 15660 13719 15712 13728
rect 15660 13685 15669 13719
rect 15669 13685 15703 13719
rect 15703 13685 15712 13719
rect 15660 13676 15712 13685
rect 2916 13574 2968 13626
rect 2980 13574 3032 13626
rect 3044 13574 3096 13626
rect 3108 13574 3160 13626
rect 3172 13574 3224 13626
rect 6849 13574 6901 13626
rect 6913 13574 6965 13626
rect 6977 13574 7029 13626
rect 7041 13574 7093 13626
rect 7105 13574 7157 13626
rect 10782 13574 10834 13626
rect 10846 13574 10898 13626
rect 10910 13574 10962 13626
rect 10974 13574 11026 13626
rect 11038 13574 11090 13626
rect 14715 13574 14767 13626
rect 14779 13574 14831 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 2228 13472 2280 13524
rect 4160 13515 4212 13524
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 4344 13515 4396 13524
rect 4344 13481 4353 13515
rect 4353 13481 4387 13515
rect 4387 13481 4396 13515
rect 4344 13472 4396 13481
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 4712 13404 4764 13456
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 11152 13336 11204 13388
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 15292 13336 15344 13388
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 7012 13268 7064 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15660 13268 15712 13320
rect 2780 13200 2832 13252
rect 3976 13243 4028 13252
rect 3976 13209 3985 13243
rect 3985 13209 4019 13243
rect 4019 13209 4028 13243
rect 3976 13200 4028 13209
rect 3884 13132 3936 13184
rect 11796 13200 11848 13252
rect 7656 13132 7708 13184
rect 4882 13030 4934 13082
rect 4946 13030 4998 13082
rect 5010 13030 5062 13082
rect 5074 13030 5126 13082
rect 5138 13030 5190 13082
rect 8815 13030 8867 13082
rect 8879 13030 8931 13082
rect 8943 13030 8995 13082
rect 9007 13030 9059 13082
rect 9071 13030 9123 13082
rect 12748 13030 12800 13082
rect 12812 13030 12864 13082
rect 12876 13030 12928 13082
rect 12940 13030 12992 13082
rect 13004 13030 13056 13082
rect 16681 13030 16733 13082
rect 16745 13030 16797 13082
rect 16809 13030 16861 13082
rect 16873 13030 16925 13082
rect 16937 13030 16989 13082
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 9220 12928 9272 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 14280 12928 14332 12980
rect 16304 12928 16356 12980
rect 2780 12860 2832 12912
rect 4160 12860 4212 12912
rect 7380 12903 7432 12912
rect 2504 12656 2556 12708
rect 6552 12792 6604 12844
rect 3884 12724 3936 12776
rect 6644 12724 6696 12776
rect 7380 12869 7389 12903
rect 7389 12869 7423 12903
rect 7423 12869 7432 12903
rect 7380 12860 7432 12869
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7840 12792 7892 12844
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 14280 12792 14332 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 1860 12588 1912 12640
rect 7288 12656 7340 12708
rect 5632 12588 5684 12640
rect 2916 12486 2968 12538
rect 2980 12486 3032 12538
rect 3044 12486 3096 12538
rect 3108 12486 3160 12538
rect 3172 12486 3224 12538
rect 6849 12486 6901 12538
rect 6913 12486 6965 12538
rect 6977 12486 7029 12538
rect 7041 12486 7093 12538
rect 7105 12486 7157 12538
rect 10782 12486 10834 12538
rect 10846 12486 10898 12538
rect 10910 12486 10962 12538
rect 10974 12486 11026 12538
rect 11038 12486 11090 12538
rect 14715 12486 14767 12538
rect 14779 12486 14831 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 6920 12384 6972 12436
rect 7196 12384 7248 12436
rect 4160 12359 4212 12368
rect 4160 12325 4169 12359
rect 4169 12325 4203 12359
rect 4203 12325 4212 12359
rect 4160 12316 4212 12325
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 2964 12180 3016 12232
rect 3240 12180 3292 12232
rect 6736 12248 6788 12300
rect 4068 12112 4120 12164
rect 6000 12180 6052 12232
rect 6644 12180 6696 12232
rect 7196 12180 7248 12232
rect 8484 12112 8536 12164
rect 3976 12044 4028 12096
rect 5540 12044 5592 12096
rect 6552 12044 6604 12096
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 4882 11942 4934 11994
rect 4946 11942 4998 11994
rect 5010 11942 5062 11994
rect 5074 11942 5126 11994
rect 5138 11942 5190 11994
rect 8815 11942 8867 11994
rect 8879 11942 8931 11994
rect 8943 11942 8995 11994
rect 9007 11942 9059 11994
rect 9071 11942 9123 11994
rect 12748 11942 12800 11994
rect 12812 11942 12864 11994
rect 12876 11942 12928 11994
rect 12940 11942 12992 11994
rect 13004 11942 13056 11994
rect 16681 11942 16733 11994
rect 16745 11942 16797 11994
rect 16809 11942 16861 11994
rect 16873 11942 16925 11994
rect 16937 11942 16989 11994
rect 1584 11840 1636 11892
rect 6736 11840 6788 11892
rect 2964 11815 3016 11824
rect 2964 11781 2973 11815
rect 2973 11781 3007 11815
rect 3007 11781 3016 11815
rect 2964 11772 3016 11781
rect 6920 11772 6972 11824
rect 7472 11772 7524 11824
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 4068 11704 4120 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 8484 11772 8536 11824
rect 10140 11704 10192 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 14280 11704 14332 11756
rect 15384 11704 15436 11756
rect 7288 11636 7340 11688
rect 8944 11611 8996 11620
rect 8944 11577 8953 11611
rect 8953 11577 8987 11611
rect 8987 11577 8996 11611
rect 8944 11568 8996 11577
rect 12164 11568 12216 11620
rect 6552 11500 6604 11552
rect 7196 11500 7248 11552
rect 10600 11500 10652 11552
rect 11336 11500 11388 11552
rect 16028 11500 16080 11552
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 2916 11398 2968 11450
rect 2980 11398 3032 11450
rect 3044 11398 3096 11450
rect 3108 11398 3160 11450
rect 3172 11398 3224 11450
rect 6849 11398 6901 11450
rect 6913 11398 6965 11450
rect 6977 11398 7029 11450
rect 7041 11398 7093 11450
rect 7105 11398 7157 11450
rect 10782 11398 10834 11450
rect 10846 11398 10898 11450
rect 10910 11398 10962 11450
rect 10974 11398 11026 11450
rect 11038 11398 11090 11450
rect 14715 11398 14767 11450
rect 14779 11398 14831 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 7288 11296 7340 11348
rect 10140 11296 10192 11348
rect 7656 11228 7708 11280
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 7748 11160 7800 11212
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 8944 11092 8996 11144
rect 11888 11160 11940 11212
rect 12440 11092 12492 11144
rect 12624 11092 12676 11144
rect 15476 11160 15528 11212
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 11336 11024 11388 11076
rect 13544 11067 13596 11076
rect 13544 11033 13553 11067
rect 13553 11033 13587 11067
rect 13587 11033 13596 11067
rect 13544 11024 13596 11033
rect 15292 11024 15344 11076
rect 15752 11024 15804 11076
rect 4882 10854 4934 10906
rect 4946 10854 4998 10906
rect 5010 10854 5062 10906
rect 5074 10854 5126 10906
rect 5138 10854 5190 10906
rect 8815 10854 8867 10906
rect 8879 10854 8931 10906
rect 8943 10854 8995 10906
rect 9007 10854 9059 10906
rect 9071 10854 9123 10906
rect 12748 10854 12800 10906
rect 12812 10854 12864 10906
rect 12876 10854 12928 10906
rect 12940 10854 12992 10906
rect 13004 10854 13056 10906
rect 16681 10854 16733 10906
rect 16745 10854 16797 10906
rect 16809 10854 16861 10906
rect 16873 10854 16925 10906
rect 16937 10854 16989 10906
rect 6276 10752 6328 10804
rect 7748 10752 7800 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 11888 10684 11940 10736
rect 13544 10684 13596 10736
rect 5816 10616 5868 10668
rect 7196 10616 7248 10668
rect 9312 10616 9364 10668
rect 9772 10616 9824 10668
rect 15476 10616 15528 10668
rect 13268 10548 13320 10600
rect 13544 10548 13596 10600
rect 12532 10412 12584 10464
rect 16304 10412 16356 10464
rect 2916 10310 2968 10362
rect 2980 10310 3032 10362
rect 3044 10310 3096 10362
rect 3108 10310 3160 10362
rect 3172 10310 3224 10362
rect 6849 10310 6901 10362
rect 6913 10310 6965 10362
rect 6977 10310 7029 10362
rect 7041 10310 7093 10362
rect 7105 10310 7157 10362
rect 10782 10310 10834 10362
rect 10846 10310 10898 10362
rect 10910 10310 10962 10362
rect 10974 10310 11026 10362
rect 11038 10310 11090 10362
rect 14715 10310 14767 10362
rect 14779 10310 14831 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 10600 10115 10652 10124
rect 10600 10081 10609 10115
rect 10609 10081 10643 10115
rect 10643 10081 10652 10115
rect 10600 10072 10652 10081
rect 12164 10072 12216 10124
rect 12440 10072 12492 10124
rect 15384 10072 15436 10124
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 2688 9868 2740 9920
rect 3240 9868 3292 9920
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 9220 10004 9272 10056
rect 4528 9936 4580 9988
rect 9772 9936 9824 9988
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 13544 10004 13596 10056
rect 4344 9868 4396 9920
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 9864 9868 9916 9920
rect 11888 9936 11940 9988
rect 15568 9936 15620 9988
rect 16120 9936 16172 9988
rect 11704 9868 11756 9920
rect 4882 9766 4934 9818
rect 4946 9766 4998 9818
rect 5010 9766 5062 9818
rect 5074 9766 5126 9818
rect 5138 9766 5190 9818
rect 8815 9766 8867 9818
rect 8879 9766 8931 9818
rect 8943 9766 8995 9818
rect 9007 9766 9059 9818
rect 9071 9766 9123 9818
rect 12748 9766 12800 9818
rect 12812 9766 12864 9818
rect 12876 9766 12928 9818
rect 12940 9766 12992 9818
rect 13004 9766 13056 9818
rect 16681 9766 16733 9818
rect 16745 9766 16797 9818
rect 16809 9766 16861 9818
rect 16873 9766 16925 9818
rect 16937 9766 16989 9818
rect 2412 9596 2464 9648
rect 2688 9639 2740 9648
rect 2688 9605 2697 9639
rect 2697 9605 2731 9639
rect 2731 9605 2740 9639
rect 2688 9596 2740 9605
rect 3976 9596 4028 9648
rect 3332 9460 3384 9512
rect 1584 9324 1636 9376
rect 2412 9324 2464 9376
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 5724 9528 5776 9580
rect 8484 9596 8536 9648
rect 9864 9596 9916 9648
rect 11888 9639 11940 9648
rect 11888 9605 11897 9639
rect 11897 9605 11931 9639
rect 11931 9605 11940 9639
rect 11888 9596 11940 9605
rect 12532 9639 12584 9648
rect 12532 9605 12541 9639
rect 12541 9605 12575 9639
rect 12575 9605 12584 9639
rect 12532 9596 12584 9605
rect 15568 9596 15620 9648
rect 7380 9528 7432 9580
rect 7564 9528 7616 9580
rect 11704 9528 11756 9580
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 15476 9528 15528 9580
rect 5172 9460 5224 9512
rect 7840 9460 7892 9512
rect 6092 9392 6144 9444
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 8392 9324 8444 9376
rect 9220 9460 9272 9512
rect 15752 9392 15804 9444
rect 2916 9222 2968 9274
rect 2980 9222 3032 9274
rect 3044 9222 3096 9274
rect 3108 9222 3160 9274
rect 3172 9222 3224 9274
rect 6849 9222 6901 9274
rect 6913 9222 6965 9274
rect 6977 9222 7029 9274
rect 7041 9222 7093 9274
rect 7105 9222 7157 9274
rect 10782 9222 10834 9274
rect 10846 9222 10898 9274
rect 10910 9222 10962 9274
rect 10974 9222 11026 9274
rect 11038 9222 11090 9274
rect 14715 9222 14767 9274
rect 14779 9222 14831 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 5632 8984 5684 9036
rect 5908 8984 5960 9036
rect 4896 8916 4948 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7472 8916 7524 8968
rect 12256 8916 12308 8968
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 3240 8848 3292 8900
rect 2596 8780 2648 8832
rect 5172 8891 5224 8900
rect 5172 8857 5181 8891
rect 5181 8857 5215 8891
rect 5215 8857 5224 8891
rect 5172 8848 5224 8857
rect 5540 8891 5592 8900
rect 5540 8857 5549 8891
rect 5549 8857 5583 8891
rect 5583 8857 5592 8891
rect 5540 8848 5592 8857
rect 6000 8848 6052 8900
rect 5448 8780 5500 8832
rect 5632 8780 5684 8832
rect 7380 8780 7432 8832
rect 11704 8848 11756 8900
rect 15384 8848 15436 8900
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 10416 8780 10468 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 4882 8678 4934 8730
rect 4946 8678 4998 8730
rect 5010 8678 5062 8730
rect 5074 8678 5126 8730
rect 5138 8678 5190 8730
rect 8815 8678 8867 8730
rect 8879 8678 8931 8730
rect 8943 8678 8995 8730
rect 9007 8678 9059 8730
rect 9071 8678 9123 8730
rect 12748 8678 12800 8730
rect 12812 8678 12864 8730
rect 12876 8678 12928 8730
rect 12940 8678 12992 8730
rect 13004 8678 13056 8730
rect 16681 8678 16733 8730
rect 16745 8678 16797 8730
rect 16809 8678 16861 8730
rect 16873 8678 16925 8730
rect 16937 8678 16989 8730
rect 1860 8576 1912 8628
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 9312 8576 9364 8628
rect 7564 8508 7616 8560
rect 8300 8508 8352 8560
rect 14372 8508 14424 8560
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 5448 8440 5500 8492
rect 8208 8440 8260 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 14556 8372 14608 8424
rect 7932 8304 7984 8356
rect 8392 8304 8444 8356
rect 16304 8236 16356 8288
rect 2916 8134 2968 8186
rect 2980 8134 3032 8186
rect 3044 8134 3096 8186
rect 3108 8134 3160 8186
rect 3172 8134 3224 8186
rect 6849 8134 6901 8186
rect 6913 8134 6965 8186
rect 6977 8134 7029 8186
rect 7041 8134 7093 8186
rect 7105 8134 7157 8186
rect 10782 8134 10834 8186
rect 10846 8134 10898 8186
rect 10910 8134 10962 8186
rect 10974 8134 11026 8186
rect 11038 8134 11090 8186
rect 14715 8134 14767 8186
rect 14779 8134 14831 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 8300 8032 8352 8084
rect 12900 8032 12952 8084
rect 4528 7896 4580 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8208 7828 8260 7880
rect 9496 7896 9548 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 14556 7828 14608 7880
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 15292 7760 15344 7812
rect 15936 7760 15988 7812
rect 3608 7692 3660 7744
rect 8392 7692 8444 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 4882 7590 4934 7642
rect 4946 7590 4998 7642
rect 5010 7590 5062 7642
rect 5074 7590 5126 7642
rect 5138 7590 5190 7642
rect 8815 7590 8867 7642
rect 8879 7590 8931 7642
rect 8943 7590 8995 7642
rect 9007 7590 9059 7642
rect 9071 7590 9123 7642
rect 12748 7590 12800 7642
rect 12812 7590 12864 7642
rect 12876 7590 12928 7642
rect 12940 7590 12992 7642
rect 13004 7590 13056 7642
rect 16681 7590 16733 7642
rect 16745 7590 16797 7642
rect 16809 7590 16861 7642
rect 16873 7590 16925 7642
rect 16937 7590 16989 7642
rect 2780 7488 2832 7540
rect 8484 7488 8536 7540
rect 2688 7420 2740 7472
rect 9220 7420 9272 7472
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 10324 7420 10376 7472
rect 14280 7420 14332 7472
rect 2596 7352 2648 7404
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 5540 7352 5592 7404
rect 5724 7352 5776 7404
rect 6092 7352 6144 7404
rect 8392 7352 8444 7404
rect 11152 7352 11204 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 2504 7216 2556 7268
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 4344 7148 4396 7200
rect 8208 7284 8260 7336
rect 8024 7216 8076 7268
rect 7196 7148 7248 7200
rect 8116 7148 8168 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 2916 7046 2968 7098
rect 2980 7046 3032 7098
rect 3044 7046 3096 7098
rect 3108 7046 3160 7098
rect 3172 7046 3224 7098
rect 6849 7046 6901 7098
rect 6913 7046 6965 7098
rect 6977 7046 7029 7098
rect 7041 7046 7093 7098
rect 7105 7046 7157 7098
rect 10782 7046 10834 7098
rect 10846 7046 10898 7098
rect 10910 7046 10962 7098
rect 10974 7046 11026 7098
rect 11038 7046 11090 7098
rect 14715 7046 14767 7098
rect 14779 7046 14831 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 11796 6944 11848 6996
rect 2780 6808 2832 6860
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 4528 6808 4580 6860
rect 6092 6808 6144 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4344 6740 4396 6792
rect 6644 6740 6696 6792
rect 7196 6740 7248 6792
rect 10324 6808 10376 6860
rect 11152 6808 11204 6860
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 8024 6740 8076 6792
rect 9404 6740 9456 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 4712 6672 4764 6724
rect 5448 6672 5500 6724
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 5264 6604 5316 6656
rect 5816 6604 5868 6656
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 7104 6715 7156 6724
rect 7104 6681 7113 6715
rect 7113 6681 7147 6715
rect 7147 6681 7156 6715
rect 7104 6672 7156 6681
rect 11796 6672 11848 6724
rect 14556 6715 14608 6724
rect 14556 6681 14565 6715
rect 14565 6681 14599 6715
rect 14599 6681 14608 6715
rect 14556 6672 14608 6681
rect 15844 6672 15896 6724
rect 7656 6604 7708 6656
rect 8208 6604 8260 6656
rect 13084 6604 13136 6656
rect 14372 6604 14424 6656
rect 4882 6502 4934 6554
rect 4946 6502 4998 6554
rect 5010 6502 5062 6554
rect 5074 6502 5126 6554
rect 5138 6502 5190 6554
rect 8815 6502 8867 6554
rect 8879 6502 8931 6554
rect 8943 6502 8995 6554
rect 9007 6502 9059 6554
rect 9071 6502 9123 6554
rect 12748 6502 12800 6554
rect 12812 6502 12864 6554
rect 12876 6502 12928 6554
rect 12940 6502 12992 6554
rect 13004 6502 13056 6554
rect 16681 6502 16733 6554
rect 16745 6502 16797 6554
rect 16809 6502 16861 6554
rect 16873 6502 16925 6554
rect 16937 6502 16989 6554
rect 2596 6400 2648 6452
rect 5540 6400 5592 6452
rect 7104 6400 7156 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 12624 6400 12676 6452
rect 2780 6332 2832 6384
rect 3148 6332 3200 6384
rect 9312 6332 9364 6384
rect 12256 6332 12308 6384
rect 2044 6264 2096 6316
rect 3884 6264 3936 6316
rect 7288 6264 7340 6316
rect 10048 6264 10100 6316
rect 11704 6264 11756 6316
rect 14372 6332 14424 6384
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 14556 6264 14608 6316
rect 15384 6264 15436 6316
rect 7564 6196 7616 6248
rect 11152 6196 11204 6248
rect 14464 6128 14516 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 2916 5958 2968 6010
rect 2980 5958 3032 6010
rect 3044 5958 3096 6010
rect 3108 5958 3160 6010
rect 3172 5958 3224 6010
rect 6849 5958 6901 6010
rect 6913 5958 6965 6010
rect 6977 5958 7029 6010
rect 7041 5958 7093 6010
rect 7105 5958 7157 6010
rect 10782 5958 10834 6010
rect 10846 5958 10898 6010
rect 10910 5958 10962 6010
rect 10974 5958 11026 6010
rect 11038 5958 11090 6010
rect 14715 5958 14767 6010
rect 14779 5958 14831 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 4528 5720 4580 5772
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 9496 5720 9548 5772
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 12256 5652 12308 5704
rect 3884 5584 3936 5636
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 4882 5414 4934 5466
rect 4946 5414 4998 5466
rect 5010 5414 5062 5466
rect 5074 5414 5126 5466
rect 5138 5414 5190 5466
rect 8815 5414 8867 5466
rect 8879 5414 8931 5466
rect 8943 5414 8995 5466
rect 9007 5414 9059 5466
rect 9071 5414 9123 5466
rect 12748 5414 12800 5466
rect 12812 5414 12864 5466
rect 12876 5414 12928 5466
rect 12940 5414 12992 5466
rect 13004 5414 13056 5466
rect 16681 5414 16733 5466
rect 16745 5414 16797 5466
rect 16809 5414 16861 5466
rect 16873 5414 16925 5466
rect 16937 5414 16989 5466
rect 6644 5312 6696 5364
rect 8576 5312 8628 5364
rect 2412 5244 2464 5296
rect 3884 5287 3936 5296
rect 3884 5253 3893 5287
rect 3893 5253 3927 5287
rect 3927 5253 3936 5287
rect 3884 5244 3936 5253
rect 1676 5176 1728 5228
rect 3240 5176 3292 5228
rect 5540 5244 5592 5296
rect 6092 5244 6144 5296
rect 8484 5287 8536 5296
rect 8484 5253 8493 5287
rect 8493 5253 8527 5287
rect 8527 5253 8536 5287
rect 8484 5244 8536 5253
rect 9496 5244 9548 5296
rect 5356 5108 5408 5160
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 8116 5176 8168 5228
rect 7380 5108 7432 5160
rect 4436 5040 4488 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 2916 4870 2968 4922
rect 2980 4870 3032 4922
rect 3044 4870 3096 4922
rect 3108 4870 3160 4922
rect 3172 4870 3224 4922
rect 6849 4870 6901 4922
rect 6913 4870 6965 4922
rect 6977 4870 7029 4922
rect 7041 4870 7093 4922
rect 7105 4870 7157 4922
rect 10782 4870 10834 4922
rect 10846 4870 10898 4922
rect 10910 4870 10962 4922
rect 10974 4870 11026 4922
rect 11038 4870 11090 4922
rect 14715 4870 14767 4922
rect 14779 4870 14831 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 14556 4743 14608 4752
rect 14556 4709 14565 4743
rect 14565 4709 14599 4743
rect 14599 4709 14608 4743
rect 14556 4700 14608 4709
rect 4620 4564 4672 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 5724 4632 5776 4684
rect 6000 4632 6052 4684
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 14188 4632 14240 4684
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7932 4607 7984 4616
rect 7288 4564 7340 4573
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8484 4564 8536 4616
rect 9312 4564 9364 4616
rect 10048 4564 10100 4616
rect 12348 4564 12400 4616
rect 13360 4564 13412 4616
rect 15568 4564 15620 4616
rect 4528 4539 4580 4548
rect 4528 4505 4537 4539
rect 4537 4505 4571 4539
rect 4571 4505 4580 4539
rect 4528 4496 4580 4505
rect 5540 4496 5592 4548
rect 5724 4496 5776 4548
rect 13452 4496 13504 4548
rect 14372 4496 14424 4548
rect 17040 4496 17092 4548
rect 7288 4428 7340 4480
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 9404 4428 9456 4480
rect 11336 4428 11388 4480
rect 13912 4428 13964 4480
rect 15384 4428 15436 4480
rect 4882 4326 4934 4378
rect 4946 4326 4998 4378
rect 5010 4326 5062 4378
rect 5074 4326 5126 4378
rect 5138 4326 5190 4378
rect 8815 4326 8867 4378
rect 8879 4326 8931 4378
rect 8943 4326 8995 4378
rect 9007 4326 9059 4378
rect 9071 4326 9123 4378
rect 12748 4326 12800 4378
rect 12812 4326 12864 4378
rect 12876 4326 12928 4378
rect 12940 4326 12992 4378
rect 13004 4326 13056 4378
rect 16681 4326 16733 4378
rect 16745 4326 16797 4378
rect 16809 4326 16861 4378
rect 16873 4326 16925 4378
rect 16937 4326 16989 4378
rect 3608 4224 3660 4276
rect 4436 4224 4488 4276
rect 4620 4267 4672 4276
rect 4620 4233 4629 4267
rect 4629 4233 4663 4267
rect 4663 4233 4672 4267
rect 4620 4224 4672 4233
rect 3332 4088 3384 4140
rect 4160 4088 4212 4140
rect 4620 4088 4672 4140
rect 5356 4224 5408 4276
rect 5724 4156 5776 4208
rect 7380 4156 7432 4208
rect 9220 4156 9272 4208
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 5540 4088 5592 4140
rect 7288 4088 7340 4140
rect 9588 4088 9640 4140
rect 13360 4156 13412 4208
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 14188 4224 14240 4276
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 5632 4020 5684 4072
rect 7932 4020 7984 4072
rect 3516 3884 3568 3936
rect 4804 3952 4856 4004
rect 4252 3884 4304 3936
rect 4528 3884 4580 3936
rect 4712 3884 4764 3936
rect 12900 3952 12952 4004
rect 9772 3884 9824 3936
rect 11704 3884 11756 3936
rect 11980 3884 12032 3936
rect 14280 3884 14332 3936
rect 15108 3884 15160 3936
rect 15660 4020 15712 4072
rect 2916 3782 2968 3834
rect 2980 3782 3032 3834
rect 3044 3782 3096 3834
rect 3108 3782 3160 3834
rect 3172 3782 3224 3834
rect 6849 3782 6901 3834
rect 6913 3782 6965 3834
rect 6977 3782 7029 3834
rect 7041 3782 7093 3834
rect 7105 3782 7157 3834
rect 10782 3782 10834 3834
rect 10846 3782 10898 3834
rect 10910 3782 10962 3834
rect 10974 3782 11026 3834
rect 11038 3782 11090 3834
rect 14715 3782 14767 3834
rect 14779 3782 14831 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 5632 3680 5684 3732
rect 9312 3680 9364 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 14372 3680 14424 3732
rect 4712 3655 4764 3664
rect 4712 3621 4721 3655
rect 4721 3621 4755 3655
rect 4755 3621 4764 3655
rect 4712 3612 4764 3621
rect 4804 3655 4856 3664
rect 4804 3621 4813 3655
rect 4813 3621 4847 3655
rect 4847 3621 4856 3655
rect 4804 3612 4856 3621
rect 2044 3544 2096 3596
rect 2412 3587 2464 3596
rect 2412 3553 2421 3587
rect 2421 3553 2455 3587
rect 2455 3553 2464 3587
rect 2412 3544 2464 3553
rect 3516 3544 3568 3596
rect 3332 3476 3384 3528
rect 5724 3544 5776 3596
rect 4252 3408 4304 3460
rect 5448 3476 5500 3528
rect 5816 3519 5868 3528
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 14464 3544 14516 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6092 3476 6144 3528
rect 9220 3476 9272 3528
rect 9404 3519 9456 3528
rect 9404 3485 9438 3519
rect 9438 3485 9456 3519
rect 9404 3476 9456 3485
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 11336 3519 11388 3528
rect 11336 3485 11370 3519
rect 11370 3485 11388 3519
rect 11336 3476 11388 3485
rect 15384 3519 15436 3528
rect 15384 3485 15402 3519
rect 15402 3485 15436 3519
rect 15384 3476 15436 3485
rect 15568 3476 15620 3528
rect 2780 3340 2832 3392
rect 5356 3340 5408 3392
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 6276 3340 6328 3349
rect 8116 3340 8168 3392
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 4882 3238 4934 3290
rect 4946 3238 4998 3290
rect 5010 3238 5062 3290
rect 5074 3238 5126 3290
rect 5138 3238 5190 3290
rect 8815 3238 8867 3290
rect 8879 3238 8931 3290
rect 8943 3238 8995 3290
rect 9007 3238 9059 3290
rect 9071 3238 9123 3290
rect 12748 3238 12800 3290
rect 12812 3238 12864 3290
rect 12876 3238 12928 3290
rect 12940 3238 12992 3290
rect 13004 3238 13056 3290
rect 16681 3238 16733 3290
rect 16745 3238 16797 3290
rect 16809 3238 16861 3290
rect 16873 3238 16925 3290
rect 16937 3238 16989 3290
rect 4712 3136 4764 3188
rect 5816 3136 5868 3188
rect 9220 3136 9272 3188
rect 11060 3179 11112 3188
rect 11060 3145 11069 3179
rect 11069 3145 11103 3179
rect 11103 3145 11112 3179
rect 11060 3136 11112 3145
rect 13360 3136 13412 3188
rect 14280 3136 14332 3188
rect 3332 3068 3384 3120
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 4252 3068 4304 3120
rect 4436 3111 4488 3120
rect 4436 3077 4445 3111
rect 4445 3077 4479 3111
rect 4479 3077 4488 3111
rect 4436 3068 4488 3077
rect 6000 3068 6052 3120
rect 14372 3068 14424 3120
rect 4160 3000 4212 3052
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5724 3000 5776 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2412 2932 2464 2984
rect 6092 2932 6144 2984
rect 4620 2864 4672 2916
rect 8300 3000 8352 3052
rect 9588 3000 9640 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 11980 3043 12032 3052
rect 11980 3009 12014 3043
rect 12014 3009 12032 3043
rect 11980 3000 12032 3009
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 14464 2932 14516 2984
rect 15200 2975 15252 2984
rect 15200 2941 15209 2975
rect 15209 2941 15243 2975
rect 15243 2941 15252 2975
rect 15200 2932 15252 2941
rect 13452 2864 13504 2916
rect 13268 2796 13320 2848
rect 15200 2796 15252 2848
rect 2916 2694 2968 2746
rect 2980 2694 3032 2746
rect 3044 2694 3096 2746
rect 3108 2694 3160 2746
rect 3172 2694 3224 2746
rect 6849 2694 6901 2746
rect 6913 2694 6965 2746
rect 6977 2694 7029 2746
rect 7041 2694 7093 2746
rect 7105 2694 7157 2746
rect 10782 2694 10834 2746
rect 10846 2694 10898 2746
rect 10910 2694 10962 2746
rect 10974 2694 11026 2746
rect 11038 2694 11090 2746
rect 14715 2694 14767 2746
rect 14779 2694 14831 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 14556 2592 14608 2644
rect 14464 2456 14516 2508
rect 2780 2388 2832 2440
rect 3608 2388 3660 2440
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 6276 2388 6328 2440
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 12348 2388 12400 2440
rect 13360 2388 13412 2440
rect 14372 2388 14424 2440
rect 15108 2388 15160 2440
rect 15200 2388 15252 2440
rect 2320 2320 2372 2372
rect 4160 2320 4212 2372
rect 5540 2320 5592 2372
rect 6920 2320 6972 2372
rect 8300 2320 8352 2372
rect 9680 2320 9732 2372
rect 11152 2320 11204 2372
rect 12624 2320 12676 2372
rect 15936 2363 15988 2372
rect 15936 2329 15945 2363
rect 15945 2329 15979 2363
rect 15979 2329 15988 2363
rect 15936 2320 15988 2329
rect 4882 2150 4934 2202
rect 4946 2150 4998 2202
rect 5010 2150 5062 2202
rect 5074 2150 5126 2202
rect 5138 2150 5190 2202
rect 8815 2150 8867 2202
rect 8879 2150 8931 2202
rect 8943 2150 8995 2202
rect 9007 2150 9059 2202
rect 9071 2150 9123 2202
rect 12748 2150 12800 2202
rect 12812 2150 12864 2202
rect 12876 2150 12928 2202
rect 12940 2150 12992 2202
rect 13004 2150 13056 2202
rect 16681 2150 16733 2202
rect 16745 2150 16797 2202
rect 16809 2150 16861 2202
rect 16873 2150 16925 2202
rect 16937 2150 16989 2202
rect 848 892 900 944
rect 1768 892 1820 944
rect 14096 892 14148 944
rect 15936 892 15988 944
<< metal2 >>
rect 4434 17200 4490 18000
rect 13450 17354 13506 18000
rect 13450 17338 13584 17354
rect 13450 17332 13596 17338
rect 13450 17326 13544 17332
rect 13450 17200 13506 17326
rect 13544 17274 13596 17280
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 2916 15804 3224 15813
rect 2916 15802 2922 15804
rect 2978 15802 3002 15804
rect 3058 15802 3082 15804
rect 3138 15802 3162 15804
rect 3218 15802 3224 15804
rect 2978 15750 2980 15802
rect 3160 15750 3162 15802
rect 2916 15748 2922 15750
rect 2978 15748 3002 15750
rect 3058 15748 3082 15750
rect 3138 15748 3162 15750
rect 3218 15748 3224 15750
rect 2916 15739 3224 15748
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 3976 14816 4028 14822
rect 4028 14764 4108 14770
rect 3976 14758 4108 14764
rect 3988 14742 4108 14758
rect 2916 14716 3224 14725
rect 2916 14714 2922 14716
rect 2978 14714 3002 14716
rect 3058 14714 3082 14716
rect 3138 14714 3162 14716
rect 3218 14714 3224 14716
rect 2978 14662 2980 14714
rect 3160 14662 3162 14714
rect 2916 14660 2922 14662
rect 2978 14660 3002 14662
rect 3058 14660 3082 14662
rect 3138 14660 3162 14662
rect 3218 14660 3224 14662
rect 2916 14651 3224 14660
rect 4080 14482 4108 14742
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 14006 2544 14214
rect 3988 14006 4016 14282
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2240 13530 2268 13806
rect 2916 13628 3224 13637
rect 2916 13626 2922 13628
rect 2978 13626 3002 13628
rect 3058 13626 3082 13628
rect 3138 13626 3162 13628
rect 3218 13626 3224 13628
rect 2978 13574 2980 13626
rect 3160 13574 3162 13626
rect 2916 13572 2922 13574
rect 2978 13572 3002 13574
rect 3058 13572 3082 13574
rect 3138 13572 3162 13574
rect 3218 13572 3224 13574
rect 2916 13563 3224 13572
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 2792 12918 2820 13194
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 3896 12782 3924 13126
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1872 12306 1900 12582
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11898 1624 12174
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 2516 11762 2544 12650
rect 2916 12540 3224 12549
rect 2916 12538 2922 12540
rect 2978 12538 3002 12540
rect 3058 12538 3082 12540
rect 3138 12538 3162 12540
rect 3218 12538 3224 12540
rect 2978 12486 2980 12538
rect 3160 12486 3162 12538
rect 2916 12484 2922 12486
rect 2978 12484 3002 12486
rect 3058 12484 3082 12486
rect 3138 12484 3162 12486
rect 3218 12484 3224 12486
rect 2916 12475 3224 12484
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2976 11830 3004 12174
rect 2964 11824 3016 11830
rect 2964 11766 3016 11772
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 3148 11756 3200 11762
rect 3252 11744 3280 12174
rect 3988 12102 4016 13194
rect 4080 12170 4108 14418
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13870 4200 14214
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4356 13530 4384 14962
rect 4448 14618 4476 17200
rect 6849 15804 7157 15813
rect 6849 15802 6855 15804
rect 6911 15802 6935 15804
rect 6991 15802 7015 15804
rect 7071 15802 7095 15804
rect 7151 15802 7157 15804
rect 6911 15750 6913 15802
rect 7093 15750 7095 15802
rect 6849 15748 6855 15750
rect 6911 15748 6935 15750
rect 6991 15748 7015 15750
rect 7071 15748 7095 15750
rect 7151 15748 7157 15750
rect 6849 15739 7157 15748
rect 10782 15804 11090 15813
rect 10782 15802 10788 15804
rect 10844 15802 10868 15804
rect 10924 15802 10948 15804
rect 11004 15802 11028 15804
rect 11084 15802 11090 15804
rect 10844 15750 10846 15802
rect 11026 15750 11028 15802
rect 10782 15748 10788 15750
rect 10844 15748 10868 15750
rect 10924 15748 10948 15750
rect 11004 15748 11028 15750
rect 11084 15748 11090 15750
rect 10782 15739 11090 15748
rect 14476 15502 14504 17274
rect 14715 15804 15023 15813
rect 14715 15802 14721 15804
rect 14777 15802 14801 15804
rect 14857 15802 14881 15804
rect 14937 15802 14961 15804
rect 15017 15802 15023 15804
rect 14777 15750 14779 15802
rect 14959 15750 14961 15802
rect 14715 15748 14721 15750
rect 14777 15748 14801 15750
rect 14857 15748 14881 15750
rect 14937 15748 14961 15750
rect 15017 15748 15023 15750
rect 14715 15739 15023 15748
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 15026 4844 15302
rect 4882 15260 5190 15269
rect 4882 15258 4888 15260
rect 4944 15258 4968 15260
rect 5024 15258 5048 15260
rect 5104 15258 5128 15260
rect 5184 15258 5190 15260
rect 4944 15206 4946 15258
rect 5126 15206 5128 15258
rect 4882 15204 4888 15206
rect 4944 15204 4968 15206
rect 5024 15204 5048 15206
rect 5104 15204 5128 15206
rect 5184 15204 5190 15206
rect 4882 15195 5190 15204
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 5920 14482 5948 14758
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 4882 14172 5190 14181
rect 4882 14170 4888 14172
rect 4944 14170 4968 14172
rect 5024 14170 5048 14172
rect 5104 14170 5128 14172
rect 5184 14170 5190 14172
rect 4944 14118 4946 14170
rect 5126 14118 5128 14170
rect 4882 14116 4888 14118
rect 4944 14116 4968 14118
rect 5024 14116 5048 14118
rect 5104 14116 5128 14118
rect 5184 14116 5190 14118
rect 4882 14107 5190 14116
rect 5644 14074 5672 14350
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12374 4200 12854
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4080 11762 4108 12106
rect 3200 11716 3280 11744
rect 3148 11698 3200 11704
rect 2916 11452 3224 11461
rect 2916 11450 2922 11452
rect 2978 11450 3002 11452
rect 3058 11450 3082 11452
rect 3138 11450 3162 11452
rect 3218 11450 3224 11452
rect 2978 11398 2980 11450
rect 3160 11398 3162 11450
rect 2916 11396 2922 11398
rect 2978 11396 3002 11398
rect 3058 11396 3082 11398
rect 3138 11396 3162 11398
rect 3218 11396 3224 11398
rect 2916 11387 3224 11396
rect 2916 10364 3224 10373
rect 2916 10362 2922 10364
rect 2978 10362 3002 10364
rect 3058 10362 3082 10364
rect 3138 10362 3162 10364
rect 3218 10362 3224 10364
rect 2978 10310 2980 10362
rect 3160 10310 3162 10362
rect 2916 10308 2922 10310
rect 2978 10308 3002 10310
rect 3058 10308 3082 10310
rect 3138 10308 3162 10310
rect 3218 10308 3224 10310
rect 2916 10299 3224 10308
rect 3252 10062 3280 11716
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2424 9654 2452 9998
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 2700 9654 2728 9862
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2424 9382 2452 9590
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1596 9042 1624 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8634 1900 8842
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2608 8498 2636 8774
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2608 7410 2636 8434
rect 2700 7478 2728 9590
rect 2916 9276 3224 9285
rect 2916 9274 2922 9276
rect 2978 9274 3002 9276
rect 3058 9274 3082 9276
rect 3138 9274 3162 9276
rect 3218 9274 3224 9276
rect 2978 9222 2980 9274
rect 3160 9222 3162 9274
rect 2916 9220 2922 9222
rect 2978 9220 3002 9222
rect 3058 9220 3082 9222
rect 3138 9220 3162 9222
rect 3218 9220 3224 9222
rect 2916 9211 3224 9220
rect 3252 8906 3280 9862
rect 3344 9518 3372 11698
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3988 9654 4016 9930
rect 4356 9926 4384 9998
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 2916 8188 3224 8197
rect 2916 8186 2922 8188
rect 2978 8186 3002 8188
rect 3058 8186 3082 8188
rect 3138 8186 3162 8188
rect 3218 8186 3224 8188
rect 2978 8134 2980 8186
rect 3160 8134 3162 8186
rect 2916 8132 2922 8134
rect 2978 8132 3002 8134
rect 3058 8132 3082 8134
rect 3138 8132 3162 8134
rect 3218 8132 3224 8134
rect 2916 8123 3224 8132
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6322 2084 7142
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5234 1716 6054
rect 2516 5710 2544 7210
rect 2792 6866 2820 7482
rect 3620 7410 3648 7686
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 4356 7206 4384 9862
rect 4540 7954 4568 9930
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 2916 7100 3224 7109
rect 2916 7098 2922 7100
rect 2978 7098 3002 7100
rect 3058 7098 3082 7100
rect 3138 7098 3162 7100
rect 3218 7098 3224 7100
rect 2978 7046 2980 7098
rect 3160 7046 3162 7098
rect 2916 7044 2922 7046
rect 2978 7044 3002 7046
rect 3058 7044 3082 7046
rect 3138 7044 3162 7046
rect 3218 7044 3224 7046
rect 2916 7035 3224 7044
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6458 2636 6734
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2792 6390 2820 6802
rect 4356 6798 4384 7142
rect 4540 6866 4568 7890
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6390 3188 6598
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 2916 6012 3224 6021
rect 2916 6010 2922 6012
rect 2978 6010 3002 6012
rect 3058 6010 3082 6012
rect 3138 6010 3162 6012
rect 3218 6010 3224 6012
rect 2978 5958 2980 6010
rect 3160 5958 3162 6010
rect 2916 5956 2922 5958
rect 2978 5956 3002 5958
rect 3058 5956 3082 5958
rect 3138 5956 3162 5958
rect 3218 5956 3224 5958
rect 2916 5947 3224 5956
rect 3344 5710 3372 6734
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3896 5642 3924 6258
rect 4540 5778 4568 6802
rect 4724 6730 4752 13398
rect 6288 13326 6316 15438
rect 8815 15260 9123 15269
rect 8815 15258 8821 15260
rect 8877 15258 8901 15260
rect 8957 15258 8981 15260
rect 9037 15258 9061 15260
rect 9117 15258 9123 15260
rect 8877 15206 8879 15258
rect 9059 15206 9061 15258
rect 8815 15204 8821 15206
rect 8877 15204 8901 15206
rect 8957 15204 8981 15206
rect 9037 15204 9061 15206
rect 9117 15204 9123 15206
rect 8815 15195 9123 15204
rect 10612 15026 10640 15438
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 6849 14716 7157 14725
rect 6849 14714 6855 14716
rect 6911 14714 6935 14716
rect 6991 14714 7015 14716
rect 7071 14714 7095 14716
rect 7151 14714 7157 14716
rect 6911 14662 6913 14714
rect 7093 14662 7095 14714
rect 6849 14660 6855 14662
rect 6911 14660 6935 14662
rect 6991 14660 7015 14662
rect 7071 14660 7095 14662
rect 7151 14660 7157 14662
rect 6849 14651 7157 14660
rect 7392 14550 7420 14962
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 13938 6592 14418
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6656 14074 6684 14282
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6748 13938 6776 14214
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 4882 13084 5190 13093
rect 4882 13082 4888 13084
rect 4944 13082 4968 13084
rect 5024 13082 5048 13084
rect 5104 13082 5128 13084
rect 5184 13082 5190 13084
rect 4944 13030 4946 13082
rect 5126 13030 5128 13082
rect 4882 13028 4888 13030
rect 4944 13028 4968 13030
rect 5024 13028 5048 13030
rect 5104 13028 5128 13030
rect 5184 13028 5190 13030
rect 4882 13019 5190 13028
rect 6564 12850 6592 13874
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 4882 11996 5190 12005
rect 4882 11994 4888 11996
rect 4944 11994 4968 11996
rect 5024 11994 5048 11996
rect 5104 11994 5128 11996
rect 5184 11994 5190 11996
rect 4944 11942 4946 11994
rect 5126 11942 5128 11994
rect 4882 11940 4888 11942
rect 4944 11940 4968 11942
rect 5024 11940 5048 11942
rect 5104 11940 5128 11942
rect 5184 11940 5190 11942
rect 4882 11931 5190 11940
rect 4882 10908 5190 10917
rect 4882 10906 4888 10908
rect 4944 10906 4968 10908
rect 5024 10906 5048 10908
rect 5104 10906 5128 10908
rect 5184 10906 5190 10908
rect 4944 10854 4946 10906
rect 5126 10854 5128 10906
rect 4882 10852 4888 10854
rect 4944 10852 4968 10854
rect 5024 10852 5048 10854
rect 5104 10852 5128 10854
rect 5184 10852 5190 10854
rect 4882 10843 5190 10852
rect 4882 9820 5190 9829
rect 4882 9818 4888 9820
rect 4944 9818 4968 9820
rect 5024 9818 5048 9820
rect 5104 9818 5128 9820
rect 5184 9818 5190 9820
rect 4944 9766 4946 9818
rect 5126 9766 5128 9818
rect 4882 9764 4888 9766
rect 4944 9764 4968 9766
rect 5024 9764 5048 9766
rect 5104 9764 5128 9766
rect 5184 9764 5190 9766
rect 4882 9755 5190 9764
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8974 4936 9318
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5184 8906 5212 9454
rect 5552 8906 5580 12038
rect 5644 9586 5672 12582
rect 6656 12238 6684 12718
rect 6748 12306 6776 13874
rect 6849 13628 7157 13637
rect 6849 13626 6855 13628
rect 6911 13626 6935 13628
rect 6991 13626 7015 13628
rect 7071 13626 7095 13628
rect 7151 13626 7157 13628
rect 6911 13574 6913 13626
rect 7093 13574 7095 13626
rect 6849 13572 6855 13574
rect 6911 13572 6935 13574
rect 6991 13572 7015 13574
rect 7071 13572 7095 13574
rect 7151 13572 7157 13574
rect 6849 13563 7157 13572
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12986 7052 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7392 12918 7420 14486
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7656 13184 7708 13190
rect 7708 13132 7788 13138
rect 7656 13126 7788 13132
rect 7668 13110 7788 13126
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 6849 12540 7157 12549
rect 6849 12538 6855 12540
rect 6911 12538 6935 12540
rect 6991 12538 7015 12540
rect 7071 12538 7095 12540
rect 7151 12538 7157 12540
rect 6911 12486 6913 12538
rect 7093 12486 7095 12538
rect 6849 12484 6855 12486
rect 6911 12484 6935 12486
rect 6991 12484 7015 12486
rect 7071 12484 7095 12486
rect 7151 12484 7157 12486
rect 6849 12475 7157 12484
rect 7208 12442 7236 12786
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9058 5764 9522
rect 5644 9042 5764 9058
rect 5632 9036 5764 9042
rect 5684 9030 5764 9036
rect 5632 8978 5684 8984
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 4882 8732 5190 8741
rect 4882 8730 4888 8732
rect 4944 8730 4968 8732
rect 5024 8730 5048 8732
rect 5104 8730 5128 8732
rect 5184 8730 5190 8732
rect 4944 8678 4946 8730
rect 5126 8678 5128 8730
rect 4882 8676 4888 8678
rect 4944 8676 4968 8678
rect 5024 8676 5048 8678
rect 5104 8676 5128 8678
rect 5184 8676 5190 8678
rect 4882 8667 5190 8676
rect 5460 8498 5488 8774
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 4882 7644 5190 7653
rect 4882 7642 4888 7644
rect 4944 7642 4968 7644
rect 5024 7642 5048 7644
rect 5104 7642 5128 7644
rect 5184 7642 5190 7644
rect 4944 7590 4946 7642
rect 5126 7590 5128 7642
rect 4882 7588 4888 7590
rect 4944 7588 4968 7590
rect 5024 7588 5048 7590
rect 5104 7588 5128 7590
rect 5184 7588 5190 7590
rect 4882 7579 5190 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5552 6882 5580 7346
rect 5460 6854 5580 6882
rect 5460 6730 5488 6854
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4882 6556 5190 6565
rect 4882 6554 4888 6556
rect 4944 6554 4968 6556
rect 5024 6554 5048 6556
rect 5104 6554 5128 6556
rect 5184 6554 5190 6556
rect 4944 6502 4946 6554
rect 5126 6502 5128 6554
rect 4882 6500 4888 6502
rect 4944 6500 4968 6502
rect 5024 6500 5048 6502
rect 5104 6500 5128 6502
rect 5184 6500 5190 6502
rect 4882 6491 5190 6500
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 2424 5302 2452 5510
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 3252 5234 3280 5510
rect 3896 5302 3924 5578
rect 4882 5468 5190 5477
rect 4882 5466 4888 5468
rect 4944 5466 4968 5468
rect 5024 5466 5048 5468
rect 5104 5466 5128 5468
rect 5184 5466 5190 5468
rect 4944 5414 4946 5466
rect 5126 5414 5128 5466
rect 4882 5412 4888 5414
rect 4944 5412 4968 5414
rect 5024 5412 5048 5414
rect 5104 5412 5128 5414
rect 5184 5412 5190 5414
rect 4882 5403 5190 5412
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 2916 4924 3224 4933
rect 2916 4922 2922 4924
rect 2978 4922 3002 4924
rect 3058 4922 3082 4924
rect 3138 4922 3162 4924
rect 3218 4922 3224 4924
rect 2978 4870 2980 4922
rect 3160 4870 3162 4922
rect 2916 4868 2922 4870
rect 2978 4868 3002 4870
rect 3058 4868 3082 4870
rect 3138 4868 3162 4870
rect 3218 4868 3224 4870
rect 2916 4859 3224 4868
rect 4448 4282 4476 5034
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 2916 3836 3224 3845
rect 2916 3834 2922 3836
rect 2978 3834 3002 3836
rect 3058 3834 3082 3836
rect 3138 3834 3162 3836
rect 3218 3834 3224 3836
rect 2978 3782 2980 3834
rect 3160 3782 3162 3834
rect 2916 3780 2922 3782
rect 2978 3780 3002 3782
rect 3058 3780 3082 3782
rect 3138 3780 3162 3782
rect 3218 3780 3224 3782
rect 2916 3771 3224 3780
rect 3344 3738 3372 4082
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3528 3602 3556 3878
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 2056 3058 2084 3538
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2424 2990 2452 3538
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 1780 950 1808 2926
rect 2792 2446 2820 3334
rect 3344 3126 3372 3470
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 2916 2748 3224 2757
rect 2916 2746 2922 2748
rect 2978 2746 3002 2748
rect 3058 2746 3082 2748
rect 3138 2746 3162 2748
rect 3218 2746 3224 2748
rect 2978 2694 2980 2746
rect 3160 2694 3162 2746
rect 2916 2692 2922 2694
rect 2978 2692 3002 2694
rect 3058 2692 3082 2694
rect 3138 2692 3162 2694
rect 3218 2692 3224 2694
rect 2916 2683 3224 2692
rect 3620 2446 3648 4218
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 3058 4200 4082
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 3466 4292 3878
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4264 3126 4292 3402
rect 4448 3126 4476 4218
rect 4540 3942 4568 4490
rect 4632 4282 4660 4558
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4632 2922 4660 4082
rect 4816 4010 4844 4966
rect 4882 4380 5190 4389
rect 4882 4378 4888 4380
rect 4944 4378 4968 4380
rect 5024 4378 5048 4380
rect 5104 4378 5128 4380
rect 5184 4378 5190 4380
rect 4944 4326 4946 4378
rect 5126 4326 5128 4378
rect 4882 4324 4888 4326
rect 4944 4324 4968 4326
rect 5024 4324 5048 4326
rect 5104 4324 5128 4326
rect 5184 4324 5190 4326
rect 4882 4315 5190 4324
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3670 4752 3878
rect 4816 3670 4844 3946
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4724 3194 4752 3606
rect 4882 3292 5190 3301
rect 4882 3290 4888 3292
rect 4944 3290 4968 3292
rect 5024 3290 5048 3292
rect 5104 3290 5128 3292
rect 5184 3290 5190 3292
rect 4944 3238 4946 3290
rect 5126 3238 5128 3290
rect 4882 3236 4888 3238
rect 4944 3236 4968 3238
rect 5024 3236 5048 3238
rect 5104 3236 5128 3238
rect 5184 3236 5190 3238
rect 4882 3227 5190 3236
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5276 3058 5304 6598
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4622 5396 5102
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4282 5396 4558
rect 5552 4554 5580 5238
rect 5644 5234 5672 8774
rect 5736 7410 5764 9030
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5828 6662 5856 10610
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9042 5948 9318
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6012 8906 6040 12174
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11762 6592 12038
rect 6748 11898 6776 12242
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6932 11830 6960 12378
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 7208 11558 7236 12174
rect 7300 11694 7328 12650
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11830 7512 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6564 11218 6592 11494
rect 6849 11452 7157 11461
rect 6849 11450 6855 11452
rect 6911 11450 6935 11452
rect 6991 11450 7015 11452
rect 7071 11450 7095 11452
rect 7151 11450 7157 11452
rect 6911 11398 6913 11450
rect 7093 11398 7095 11450
rect 6849 11396 6855 11398
rect 6911 11396 6935 11398
rect 6991 11396 7015 11398
rect 7071 11396 7095 11398
rect 7151 11396 7157 11398
rect 6849 11387 7157 11396
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10810 6316 11086
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 7208 10674 7236 11494
rect 7300 11354 7328 11630
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 6849 10364 7157 10373
rect 6849 10362 6855 10364
rect 6911 10362 6935 10364
rect 6991 10362 7015 10364
rect 7071 10362 7095 10364
rect 7151 10362 7157 10364
rect 6911 10310 6913 10362
rect 7093 10310 7095 10362
rect 6849 10308 6855 10310
rect 6911 10308 6935 10310
rect 6991 10308 7015 10310
rect 7071 10308 7095 10310
rect 7151 10308 7157 10310
rect 6849 10299 7157 10308
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6104 7410 6132 9386
rect 6849 9276 7157 9285
rect 6849 9274 6855 9276
rect 6911 9274 6935 9276
rect 6991 9274 7015 9276
rect 7071 9274 7095 9276
rect 7151 9274 7157 9276
rect 6911 9222 6913 9274
rect 7093 9222 7095 9274
rect 6849 9220 6855 9222
rect 6911 9220 6935 9222
rect 6991 9220 7015 9222
rect 7071 9220 7095 9222
rect 7151 9220 7157 9222
rect 6849 9211 7157 9220
rect 7392 8974 7420 9522
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 6849 8188 7157 8197
rect 6849 8186 6855 8188
rect 6911 8186 6935 8188
rect 6991 8186 7015 8188
rect 7071 8186 7095 8188
rect 7151 8186 7157 8188
rect 6911 8134 6913 8186
rect 7093 8134 7095 8186
rect 6849 8132 6855 8134
rect 6911 8132 6935 8134
rect 6991 8132 7015 8134
rect 7071 8132 7095 8134
rect 7151 8132 7157 8134
rect 6849 8123 7157 8132
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 6866 6132 7346
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6849 7100 7157 7109
rect 6849 7098 6855 7100
rect 6911 7098 6935 7100
rect 6991 7098 7015 7100
rect 7071 7098 7095 7100
rect 7151 7098 7157 7100
rect 6911 7046 6913 7098
rect 7093 7046 7095 7098
rect 6849 7044 6855 7046
rect 6911 7044 6935 7046
rect 6991 7044 7015 7046
rect 7071 7044 7095 7046
rect 7151 7044 7157 7046
rect 6849 7035 7157 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 7208 6798 7236 7142
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 5302 6132 6598
rect 6656 5370 6684 6734
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7116 6458 7144 6666
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 6849 6012 7157 6021
rect 6849 6010 6855 6012
rect 6911 6010 6935 6012
rect 6991 6010 7015 6012
rect 7071 6010 7095 6012
rect 7151 6010 7157 6012
rect 6911 5958 6913 6010
rect 7093 5958 7095 6010
rect 6849 5956 6855 5958
rect 6911 5956 6935 5958
rect 6991 5956 7015 5958
rect 7071 5956 7095 5958
rect 7151 5956 7157 5958
rect 6849 5947 7157 5956
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4842 5672 5170
rect 5644 4814 5764 4842
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5552 4146 5580 4490
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5460 3534 5488 4082
rect 5644 4078 5672 4694
rect 5736 4690 5764 4814
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5736 4214 5764 4490
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 3738 5672 4014
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5736 3602 5764 4150
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 5368 2446 5396 3334
rect 5736 3058 5764 3538
rect 6012 3534 6040 4626
rect 6656 4622 6684 5306
rect 6849 4924 7157 4933
rect 6849 4922 6855 4924
rect 6911 4922 6935 4924
rect 6991 4922 7015 4924
rect 7071 4922 7095 4924
rect 7151 4922 7157 4924
rect 6911 4870 6913 4922
rect 7093 4870 7095 4922
rect 6849 4868 6855 4870
rect 6911 4868 6935 4870
rect 6991 4868 7015 4870
rect 7071 4868 7095 4870
rect 7151 4868 7157 4870
rect 6849 4859 7157 4868
rect 7300 4622 7328 6258
rect 7392 5166 7420 8774
rect 7484 8634 7512 8910
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8566 7604 9522
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7576 6254 7604 8502
rect 7668 6662 7696 11222
rect 7760 11218 7788 13110
rect 7852 12850 7880 13670
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10810 7788 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7852 9518 7880 12786
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 8312 8566 8340 14554
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8496 13530 8524 14418
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8815 14172 9123 14181
rect 8815 14170 8821 14172
rect 8877 14170 8901 14172
rect 8957 14170 8981 14172
rect 9037 14170 9061 14172
rect 9117 14170 9123 14172
rect 8877 14118 8879 14170
rect 9059 14118 9061 14170
rect 8815 14116 8821 14118
rect 8877 14116 8901 14118
rect 8957 14116 8981 14118
rect 9037 14116 9061 14118
rect 9117 14116 9123 14118
rect 8815 14107 9123 14116
rect 9232 14006 9260 14214
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9508 13938 9536 14758
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8496 12170 8524 13466
rect 8815 13084 9123 13093
rect 8815 13082 8821 13084
rect 8877 13082 8901 13084
rect 8957 13082 8981 13084
rect 9037 13082 9061 13084
rect 9117 13082 9123 13084
rect 8877 13030 8879 13082
rect 9059 13030 9061 13082
rect 8815 13028 8821 13030
rect 8877 13028 8901 13030
rect 8957 13028 8981 13030
rect 9037 13028 9061 13030
rect 9117 13028 9123 13030
rect 8815 13019 9123 13028
rect 9232 12986 9260 13806
rect 9876 13394 9904 14758
rect 10612 14414 10640 14962
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 10782 14716 11090 14725
rect 10782 14714 10788 14716
rect 10844 14714 10868 14716
rect 10924 14714 10948 14716
rect 11004 14714 11028 14716
rect 11084 14714 11090 14716
rect 10844 14662 10846 14714
rect 11026 14662 11028 14714
rect 10782 14660 10788 14662
rect 10844 14660 10868 14662
rect 10924 14660 10948 14662
rect 11004 14660 11028 14662
rect 11084 14660 11090 14662
rect 10782 14651 11090 14660
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 11164 13938 11192 14894
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14346 11560 14758
rect 11900 14482 11928 14962
rect 11992 14482 12020 15302
rect 12748 15260 13056 15269
rect 12748 15258 12754 15260
rect 12810 15258 12834 15260
rect 12890 15258 12914 15260
rect 12970 15258 12994 15260
rect 13050 15258 13056 15260
rect 12810 15206 12812 15258
rect 12992 15206 12994 15258
rect 12748 15204 12754 15206
rect 12810 15204 12834 15206
rect 12890 15204 12914 15206
rect 12970 15204 12994 15206
rect 13050 15204 13056 15206
rect 12748 15195 13056 15204
rect 13832 15026 13860 15370
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 14482 12296 14758
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13394 10180 13670
rect 10782 13628 11090 13637
rect 10782 13626 10788 13628
rect 10844 13626 10868 13628
rect 10924 13626 10948 13628
rect 11004 13626 11028 13628
rect 11084 13626 11090 13628
rect 10844 13574 10846 13626
rect 11026 13574 11028 13626
rect 10782 13572 10788 13574
rect 10844 13572 10868 13574
rect 10924 13572 10948 13574
rect 11004 13572 11028 13574
rect 11084 13572 11090 13574
rect 10782 13563 11090 13572
rect 11164 13394 11192 13874
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12850 11928 14418
rect 12544 14414 12572 14962
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12748 14172 13056 14181
rect 12748 14170 12754 14172
rect 12810 14170 12834 14172
rect 12890 14170 12914 14172
rect 12970 14170 12994 14172
rect 13050 14170 13056 14172
rect 12810 14118 12812 14170
rect 12992 14118 12994 14170
rect 12748 14116 12754 14118
rect 12810 14116 12834 14118
rect 12890 14116 12914 14118
rect 12970 14116 12994 14118
rect 13050 14116 13056 14118
rect 12748 14107 13056 14116
rect 13096 13938 13124 14758
rect 13832 14482 13860 14962
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 14006 13400 14214
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 10782 12540 11090 12549
rect 10782 12538 10788 12540
rect 10844 12538 10868 12540
rect 10924 12538 10948 12540
rect 11004 12538 11028 12540
rect 11084 12538 11090 12540
rect 10844 12486 10846 12538
rect 11026 12486 11028 12538
rect 10782 12484 10788 12486
rect 10844 12484 10868 12486
rect 10924 12484 10948 12486
rect 11004 12484 11028 12486
rect 11084 12484 11090 12486
rect 10782 12475 11090 12484
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11830 8524 12106
rect 8815 11996 9123 12005
rect 8815 11994 8821 11996
rect 8877 11994 8901 11996
rect 8957 11994 8981 11996
rect 9037 11994 9061 11996
rect 9117 11994 9123 11996
rect 8877 11942 8879 11994
rect 9059 11942 9061 11994
rect 8815 11940 8821 11942
rect 8877 11940 8901 11942
rect 8957 11940 8981 11942
rect 9037 11940 9061 11942
rect 9117 11940 9123 11942
rect 8815 11931 9123 11940
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 11900 11762 11928 12786
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11150 8984 11562
rect 10152 11354 10180 11698
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 8815 10908 9123 10917
rect 8815 10906 8821 10908
rect 8877 10906 8901 10908
rect 8957 10906 8981 10908
rect 9037 10906 9061 10908
rect 9117 10906 9123 10908
rect 8877 10854 8879 10906
rect 9059 10854 9061 10906
rect 8815 10852 8821 10854
rect 8877 10852 8901 10854
rect 8957 10852 8981 10854
rect 9037 10852 9061 10854
rect 9117 10852 9123 10854
rect 8815 10843 9123 10852
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9654 8524 9862
rect 8815 9820 9123 9829
rect 8815 9818 8821 9820
rect 8877 9818 8901 9820
rect 8957 9818 8981 9820
rect 9037 9818 9061 9820
rect 9117 9818 9123 9820
rect 8877 9766 8879 9818
rect 9059 9766 9061 9818
rect 8815 9764 8821 9766
rect 8877 9764 8901 9766
rect 8957 9764 8981 9766
rect 9037 9764 9061 9766
rect 9117 9764 9123 9766
rect 8815 9755 9123 9764
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 9232 9518 9260 9998
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7944 7886 7972 8298
rect 8220 7886 8248 8434
rect 8404 8362 8432 9318
rect 8815 8732 9123 8741
rect 8815 8730 8821 8732
rect 8877 8730 8901 8732
rect 8957 8730 8981 8732
rect 9037 8730 9061 8732
rect 9117 8730 9123 8732
rect 8877 8678 8879 8730
rect 9059 8678 9061 8730
rect 8815 8676 8821 8678
rect 8877 8676 8901 8678
rect 8957 8676 8981 8678
rect 9037 8676 9061 8678
rect 9117 8676 9123 8678
rect 8815 8667 9123 8676
rect 9324 8634 9352 10610
rect 9784 9994 9812 10610
rect 10060 10266 10088 11018
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10152 10062 10180 11290
rect 10612 10130 10640 11494
rect 10782 11452 11090 11461
rect 10782 11450 10788 11452
rect 10844 11450 10868 11452
rect 10924 11450 10948 11452
rect 11004 11450 11028 11452
rect 11084 11450 11090 11452
rect 10844 11398 10846 11450
rect 11026 11398 11028 11450
rect 10782 11396 10788 11398
rect 10844 11396 10868 11398
rect 10924 11396 10948 11398
rect 11004 11396 11028 11398
rect 11084 11396 11090 11398
rect 10782 11387 11090 11396
rect 11348 11082 11376 11494
rect 11900 11218 11928 11698
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11900 10742 11928 11154
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 10782 10364 11090 10373
rect 10782 10362 10788 10364
rect 10844 10362 10868 10364
rect 10924 10362 10948 10364
rect 11004 10362 11028 10364
rect 11084 10362 11090 10364
rect 10844 10310 10846 10362
rect 11026 10310 11028 10362
rect 10782 10308 10788 10310
rect 10844 10308 10868 10310
rect 10924 10308 10948 10310
rect 11004 10308 11028 10310
rect 11084 10308 11090 10310
rect 10782 10299 11090 10308
rect 12176 10130 12204 11562
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 9784 8838 9812 9930
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 9876 9654 9904 9862
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 11716 9586 11744 9862
rect 11900 9654 11928 9930
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 10782 9276 11090 9285
rect 10782 9274 10788 9276
rect 10844 9274 10868 9276
rect 10924 9274 10948 9276
rect 11004 9274 11028 9276
rect 11084 9274 11090 9276
rect 10844 9222 10846 9274
rect 11026 9222 11028 9274
rect 10782 9220 10788 9222
rect 10844 9220 10868 9222
rect 10924 9220 10948 9222
rect 11004 9220 11028 9222
rect 11084 9220 11090 9222
rect 10782 9211 11090 9220
rect 11716 8906 11744 9522
rect 12268 8974 12296 13806
rect 12452 11150 12480 13874
rect 14108 13870 14136 15302
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14384 14006 14412 14758
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 12748 13084 13056 13093
rect 12748 13082 12754 13084
rect 12810 13082 12834 13084
rect 12890 13082 12914 13084
rect 12970 13082 12994 13084
rect 13050 13082 13056 13084
rect 12810 13030 12812 13082
rect 12992 13030 12994 13082
rect 12748 13028 12754 13030
rect 12810 13028 12834 13030
rect 12890 13028 12914 13030
rect 12970 13028 12994 13030
rect 13050 13028 13056 13030
rect 12748 13019 13056 13028
rect 12748 11996 13056 12005
rect 12748 11994 12754 11996
rect 12810 11994 12834 11996
rect 12890 11994 12914 11996
rect 12970 11994 12994 11996
rect 13050 11994 13056 11996
rect 12810 11942 12812 11994
rect 12992 11942 12994 11994
rect 12748 11940 12754 11942
rect 12810 11940 12834 11942
rect 12890 11940 12914 11942
rect 12970 11940 12994 11942
rect 13050 11940 13056 11942
rect 12748 11931 13056 11940
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12544 10554 12572 11698
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12452 10526 12572 10554
rect 12452 10130 12480 10526
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9586 12480 10066
rect 12544 9654 12572 10406
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7944 7256 7972 7822
rect 8220 7426 8248 7822
rect 8128 7398 8248 7426
rect 8024 7268 8076 7274
rect 7944 7228 8024 7256
rect 8024 7210 8076 7216
rect 8036 6798 8064 7210
rect 8128 7206 8156 7398
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8128 5234 8156 7142
rect 8220 6662 8248 7278
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 8128 4622 8156 5170
rect 8220 4622 8248 6598
rect 8312 6458 8340 8026
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8404 7410 8432 7686
rect 8496 7546 8524 7686
rect 8815 7644 9123 7653
rect 8815 7642 8821 7644
rect 8877 7642 8901 7644
rect 8957 7642 8981 7644
rect 9037 7642 9061 7644
rect 9117 7642 9123 7644
rect 8877 7590 8879 7642
rect 9059 7590 9061 7642
rect 8815 7588 8821 7590
rect 8877 7588 8901 7590
rect 8957 7588 8981 7590
rect 9037 7588 9061 7590
rect 9117 7588 9123 7590
rect 8815 7579 9123 7588
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 9232 7478 9260 7686
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8815 6556 9123 6565
rect 8815 6554 8821 6556
rect 8877 6554 8901 6556
rect 8957 6554 8981 6556
rect 9037 6554 9061 6556
rect 9117 6554 9123 6556
rect 8877 6502 8879 6554
rect 9059 6502 9061 6554
rect 8815 6500 8821 6502
rect 8877 6500 8901 6502
rect 8957 6500 8981 6502
rect 9037 6500 9061 6502
rect 9117 6500 9123 6502
rect 8815 6491 9123 6500
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7300 4146 7328 4422
rect 7392 4214 7420 4422
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7944 4078 7972 4558
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 6849 3836 7157 3845
rect 6849 3834 6855 3836
rect 6911 3834 6935 3836
rect 6991 3834 7015 3836
rect 7071 3834 7095 3836
rect 7151 3834 7157 3836
rect 6911 3782 6913 3834
rect 7093 3782 7095 3834
rect 6849 3780 6855 3782
rect 6911 3780 6935 3782
rect 6991 3780 7015 3782
rect 7071 3780 7095 3782
rect 7151 3780 7157 3782
rect 6849 3771 7157 3780
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5828 3194 5856 3470
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6012 3126 6040 3470
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6104 2990 6132 3470
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6288 2446 6316 3334
rect 6849 2748 7157 2757
rect 6849 2746 6855 2748
rect 6911 2746 6935 2748
rect 6991 2746 7015 2748
rect 7071 2746 7095 2748
rect 7151 2746 7157 2748
rect 6911 2694 6913 2746
rect 7093 2694 7095 2746
rect 6849 2692 6855 2694
rect 6911 2692 6935 2694
rect 6991 2692 7015 2694
rect 7071 2692 7095 2694
rect 7151 2692 7157 2694
rect 6849 2683 7157 2692
rect 8128 2446 8156 3334
rect 8312 3058 8340 6394
rect 9324 6390 9352 8570
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 6798 9444 7822
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9416 5710 9444 6734
rect 9508 5778 9536 7890
rect 10428 7886 10456 8774
rect 10782 8188 11090 8197
rect 10782 8186 10788 8188
rect 10844 8186 10868 8188
rect 10924 8186 10948 8188
rect 11004 8186 11028 8188
rect 11084 8186 11090 8188
rect 10844 8134 10846 8186
rect 11026 8134 11028 8186
rect 10782 8132 10788 8134
rect 10844 8132 10868 8134
rect 10924 8132 10948 8134
rect 11004 8132 11028 8134
rect 11084 8132 11090 8134
rect 10782 8123 11090 8132
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 11716 7750 11744 8842
rect 12636 8498 12664 11086
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 12748 10908 13056 10917
rect 12748 10906 12754 10908
rect 12810 10906 12834 10908
rect 12890 10906 12914 10908
rect 12970 10906 12994 10908
rect 13050 10906 13056 10908
rect 12810 10854 12812 10906
rect 12992 10854 12994 10906
rect 12748 10852 12754 10854
rect 12810 10852 12834 10854
rect 12890 10852 12914 10854
rect 12970 10852 12994 10854
rect 13050 10852 13056 10854
rect 12748 10843 13056 10852
rect 13556 10742 13584 11018
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13280 10266 13308 10542
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13556 10062 13584 10542
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 12748 9820 13056 9829
rect 12748 9818 12754 9820
rect 12810 9818 12834 9820
rect 12890 9818 12914 9820
rect 12970 9818 12994 9820
rect 13050 9818 13056 9820
rect 12810 9766 12812 9818
rect 12992 9766 12994 9818
rect 12748 9764 12754 9766
rect 12810 9764 12834 9766
rect 12890 9764 12914 9766
rect 12970 9764 12994 9766
rect 13050 9764 13056 9766
rect 12748 9755 13056 9764
rect 12748 8732 13056 8741
rect 12748 8730 12754 8732
rect 12810 8730 12834 8732
rect 12890 8730 12914 8732
rect 12970 8730 12994 8732
rect 13050 8730 13056 8732
rect 12810 8678 12812 8730
rect 12992 8678 12994 8730
rect 12748 8676 12754 8678
rect 12810 8676 12834 8678
rect 12890 8676 12914 8678
rect 12970 8676 12994 8678
rect 13050 8676 13056 8678
rect 12748 8667 13056 8676
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 8090 12940 8366
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10336 6866 10364 7414
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10782 7100 11090 7109
rect 10782 7098 10788 7100
rect 10844 7098 10868 7100
rect 10924 7098 10948 7100
rect 11004 7098 11028 7100
rect 11084 7098 11090 7100
rect 10844 7046 10846 7098
rect 11026 7046 11028 7098
rect 10782 7044 10788 7046
rect 10844 7044 10868 7046
rect 10924 7044 10948 7046
rect 11004 7044 11028 7046
rect 11084 7044 11090 7046
rect 10782 7035 11090 7044
rect 11164 6866 11192 7346
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6322 10088 6734
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 8576 5704 8628 5710
rect 9404 5704 9456 5710
rect 8576 5646 8628 5652
rect 9324 5664 9404 5692
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5302 8524 5510
rect 8588 5370 8616 5646
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 8815 5468 9123 5477
rect 8815 5466 8821 5468
rect 8877 5466 8901 5468
rect 8957 5466 8981 5468
rect 9037 5466 9061 5468
rect 9117 5466 9123 5468
rect 8877 5414 8879 5466
rect 9059 5414 9061 5466
rect 8815 5412 8821 5414
rect 8877 5412 8901 5414
rect 8957 5412 8981 5414
rect 9037 5412 9061 5414
rect 9117 5412 9123 5414
rect 8815 5403 9123 5412
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8496 4622 8524 5238
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8815 4380 9123 4389
rect 8815 4378 8821 4380
rect 8877 4378 8901 4380
rect 8957 4378 8981 4380
rect 9037 4378 9061 4380
rect 9117 4378 9123 4380
rect 8877 4326 8879 4378
rect 9059 4326 9061 4378
rect 8815 4324 8821 4326
rect 8877 4324 8901 4326
rect 8957 4324 8981 4326
rect 9037 4324 9061 4326
rect 9117 4324 9123 4326
rect 8815 4315 9123 4324
rect 9232 4214 9260 5510
rect 9324 4622 9352 5664
rect 9404 5646 9456 5652
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9508 4690 9536 5238
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 10060 4622 10088 6258
rect 11164 6254 11192 6802
rect 11716 6322 11744 7686
rect 12748 7644 13056 7653
rect 12748 7642 12754 7644
rect 12810 7642 12834 7644
rect 12890 7642 12914 7644
rect 12970 7642 12994 7644
rect 13050 7642 13056 7644
rect 12810 7590 12812 7642
rect 12992 7590 12994 7642
rect 12748 7588 12754 7590
rect 12810 7588 12834 7590
rect 12890 7588 12914 7590
rect 12970 7588 12994 7590
rect 13050 7588 13056 7590
rect 12748 7579 13056 7588
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 7002 11836 7142
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 14108 6914 14136 13806
rect 14568 13394 14596 14758
rect 14715 14716 15023 14725
rect 14715 14714 14721 14716
rect 14777 14714 14801 14716
rect 14857 14714 14881 14716
rect 14937 14714 14961 14716
rect 15017 14714 15023 14716
rect 14777 14662 14779 14714
rect 14959 14662 14961 14714
rect 14715 14660 14721 14662
rect 14777 14660 14801 14662
rect 14857 14660 14881 14662
rect 14937 14660 14961 14662
rect 15017 14660 15023 14662
rect 14715 14651 15023 14660
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 14006 14688 14350
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14715 13628 15023 13637
rect 14715 13626 14721 13628
rect 14777 13626 14801 13628
rect 14857 13626 14881 13628
rect 14937 13626 14961 13628
rect 15017 13626 15023 13628
rect 14777 13574 14779 13626
rect 14959 13574 14961 13626
rect 14715 13572 14721 13574
rect 14777 13572 14801 13574
rect 14857 13572 14881 13574
rect 14937 13572 14961 13574
rect 15017 13572 15023 13574
rect 14715 13563 15023 13572
rect 15304 13394 15332 14962
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14346 15608 14758
rect 16040 14482 16068 15302
rect 16681 15260 16989 15269
rect 16681 15258 16687 15260
rect 16743 15258 16767 15260
rect 16823 15258 16847 15260
rect 16903 15258 16927 15260
rect 16983 15258 16989 15260
rect 16743 15206 16745 15258
rect 16925 15206 16927 15258
rect 16681 15204 16687 15206
rect 16743 15204 16767 15206
rect 16823 15204 16847 15206
rect 16903 15204 16927 15206
rect 16983 15204 16989 15206
rect 16681 15195 16989 15204
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12986 14320 13262
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 15304 12850 15332 13330
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14292 11762 14320 12786
rect 14715 12540 15023 12549
rect 14715 12538 14721 12540
rect 14777 12538 14801 12540
rect 14857 12538 14881 12540
rect 14937 12538 14961 12540
rect 15017 12538 15023 12540
rect 14777 12486 14779 12538
rect 14959 12486 14961 12538
rect 14715 12484 14721 12486
rect 14777 12484 14801 12486
rect 14857 12484 14881 12486
rect 14937 12484 14961 12486
rect 15017 12484 15023 12486
rect 14715 12475 15023 12484
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 14292 11150 14320 11698
rect 14715 11452 15023 11461
rect 14715 11450 14721 11452
rect 14777 11450 14801 11452
rect 14857 11450 14881 11452
rect 14937 11450 14961 11452
rect 15017 11450 15023 11452
rect 14777 11398 14779 11450
rect 14959 11398 14961 11450
rect 14715 11396 14721 11398
rect 14777 11396 14801 11398
rect 14857 11396 14881 11398
rect 14937 11396 14961 11398
rect 15017 11396 15023 11398
rect 14715 11387 15023 11396
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 14715 10364 15023 10373
rect 14715 10362 14721 10364
rect 14777 10362 14801 10364
rect 14857 10362 14881 10364
rect 14937 10362 14961 10364
rect 15017 10362 15023 10364
rect 14777 10310 14779 10362
rect 14959 10310 14961 10362
rect 14715 10308 14721 10310
rect 14777 10308 14801 10310
rect 14857 10308 14881 10310
rect 14937 10308 14961 10310
rect 15017 10308 15023 10310
rect 14715 10299 15023 10308
rect 15396 10130 15424 11698
rect 15488 11218 15516 13874
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13326 15700 13670
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 16316 12986 16344 14350
rect 16681 14172 16989 14181
rect 16681 14170 16687 14172
rect 16743 14170 16767 14172
rect 16823 14170 16847 14172
rect 16903 14170 16927 14172
rect 16983 14170 16989 14172
rect 16743 14118 16745 14170
rect 16925 14118 16927 14170
rect 16681 14116 16687 14118
rect 16743 14116 16767 14118
rect 16823 14116 16847 14118
rect 16903 14116 16927 14118
rect 16983 14116 16989 14118
rect 16681 14107 16989 14116
rect 16681 13084 16989 13093
rect 16681 13082 16687 13084
rect 16743 13082 16767 13084
rect 16823 13082 16847 13084
rect 16903 13082 16927 13084
rect 16983 13082 16989 13084
rect 16743 13030 16745 13082
rect 16925 13030 16927 13082
rect 16681 13028 16687 13030
rect 16743 13028 16767 13030
rect 16823 13028 16847 13030
rect 16903 13028 16927 13030
rect 16983 13028 16989 13030
rect 16681 13019 16989 13028
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16681 11996 16989 12005
rect 16681 11994 16687 11996
rect 16743 11994 16767 11996
rect 16823 11994 16847 11996
rect 16903 11994 16927 11996
rect 16983 11994 16989 11996
rect 16743 11942 16745 11994
rect 16925 11942 16927 11994
rect 16681 11940 16687 11942
rect 16743 11940 16767 11942
rect 16823 11940 16847 11942
rect 16903 11940 16927 11942
rect 16983 11940 16989 11942
rect 16681 11931 16989 11940
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16040 11218 16068 11494
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15488 10674 15516 11154
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9586 15424 10066
rect 15488 9586 15516 10610
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15580 9654 15608 9930
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15764 9450 15792 11018
rect 16132 9994 16160 11494
rect 16681 10908 16989 10917
rect 16681 10906 16687 10908
rect 16743 10906 16767 10908
rect 16823 10906 16847 10908
rect 16903 10906 16927 10908
rect 16983 10906 16989 10908
rect 16743 10854 16745 10906
rect 16925 10854 16927 10906
rect 16681 10852 16687 10854
rect 16743 10852 16767 10854
rect 16823 10852 16847 10854
rect 16903 10852 16927 10854
rect 16983 10852 16989 10854
rect 16681 10843 16989 10852
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10130 16344 10406
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16681 9820 16989 9829
rect 16681 9818 16687 9820
rect 16743 9818 16767 9820
rect 16823 9818 16847 9820
rect 16903 9818 16927 9820
rect 16983 9818 16989 9820
rect 16743 9766 16745 9818
rect 16925 9766 16927 9818
rect 16681 9764 16687 9766
rect 16743 9764 16767 9766
rect 16823 9764 16847 9766
rect 16903 9764 16927 9766
rect 16983 9764 16989 9766
rect 16681 9755 16989 9764
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 14715 9276 15023 9285
rect 14715 9274 14721 9276
rect 14777 9274 14801 9276
rect 14857 9274 14881 9276
rect 14937 9274 14961 9276
rect 15017 9274 15023 9276
rect 14777 9222 14779 9274
rect 14959 9222 14961 9274
rect 14715 9220 14721 9222
rect 14777 9220 14801 9222
rect 14857 9220 14881 9222
rect 14937 9220 14961 9222
rect 15017 9220 15023 9222
rect 14715 9211 15023 9220
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8566 14412 8774
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7886 14596 8366
rect 14715 8188 15023 8197
rect 14715 8186 14721 8188
rect 14777 8186 14801 8188
rect 14857 8186 14881 8188
rect 14937 8186 14961 8188
rect 15017 8186 15023 8188
rect 14777 8134 14779 8186
rect 14959 8134 14961 8186
rect 14715 8132 14721 8134
rect 14777 8132 14801 8134
rect 14857 8132 14881 8134
rect 14937 8132 14961 8134
rect 15017 8132 15023 8134
rect 14715 8123 15023 8132
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 14292 7478 14320 7754
rect 15304 7546 15332 7754
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 15396 7410 15424 8842
rect 16681 8732 16989 8741
rect 16681 8730 16687 8732
rect 16743 8730 16767 8732
rect 16823 8730 16847 8732
rect 16903 8730 16927 8732
rect 16983 8730 16989 8732
rect 16743 8678 16745 8730
rect 16925 8678 16927 8730
rect 16681 8676 16687 8678
rect 16743 8676 16767 8678
rect 16823 8676 16847 8678
rect 16903 8676 16927 8678
rect 16983 8676 16989 8678
rect 16681 8667 16989 8676
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7954 16344 8230
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7546 15976 7754
rect 16681 7644 16989 7653
rect 16681 7642 16687 7644
rect 16743 7642 16767 7644
rect 16823 7642 16847 7644
rect 16903 7642 16927 7644
rect 16983 7642 16989 7644
rect 16743 7590 16745 7642
rect 16925 7590 16927 7642
rect 16681 7588 16687 7590
rect 16743 7588 16767 7590
rect 16823 7588 16847 7590
rect 16903 7588 16927 7590
rect 16983 7588 16989 7590
rect 16681 7579 16989 7588
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14108 6886 14228 6914
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11808 6458 11836 6666
rect 12636 6458 12664 6734
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12748 6556 13056 6565
rect 12748 6554 12754 6556
rect 12810 6554 12834 6556
rect 12890 6554 12914 6556
rect 12970 6554 12994 6556
rect 13050 6554 13056 6556
rect 12810 6502 12812 6554
rect 12992 6502 12994 6554
rect 12748 6500 12754 6502
rect 12810 6500 12834 6502
rect 12890 6500 12914 6502
rect 12970 6500 12994 6502
rect 13050 6500 13056 6502
rect 12748 6491 13056 6500
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10782 6012 11090 6021
rect 10782 6010 10788 6012
rect 10844 6010 10868 6012
rect 10924 6010 10948 6012
rect 11004 6010 11028 6012
rect 11084 6010 11090 6012
rect 10844 5958 10846 6010
rect 11026 5958 11028 6010
rect 10782 5956 10788 5958
rect 10844 5956 10868 5958
rect 10924 5956 10948 5958
rect 11004 5956 11028 5958
rect 11084 5956 11090 5958
rect 10782 5947 11090 5956
rect 12268 5710 12296 6326
rect 13096 6322 13124 6598
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 10782 4924 11090 4933
rect 10782 4922 10788 4924
rect 10844 4922 10868 4924
rect 10924 4922 10948 4924
rect 11004 4922 11028 4924
rect 11084 4922 11090 4924
rect 10844 4870 10846 4922
rect 11026 4870 11028 4922
rect 10782 4868 10788 4870
rect 10844 4868 10868 4870
rect 10924 4868 10948 4870
rect 11004 4868 11028 4870
rect 11084 4868 11090 4870
rect 10782 4859 11090 4868
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 9324 3738 9352 4558
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3534 9444 4422
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8815 3292 9123 3301
rect 8815 3290 8821 3292
rect 8877 3290 8901 3292
rect 8957 3290 8981 3292
rect 9037 3290 9061 3292
rect 9117 3290 9123 3292
rect 8877 3238 8879 3290
rect 9059 3238 9061 3290
rect 8815 3236 8821 3238
rect 8877 3236 8901 3238
rect 8957 3236 8981 3238
rect 9037 3236 9061 3238
rect 9117 3236 9123 3238
rect 8815 3227 9123 3236
rect 9232 3194 9260 3470
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9600 3058 9628 4082
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 2446 9812 3878
rect 10782 3836 11090 3845
rect 10782 3834 10788 3836
rect 10844 3834 10868 3836
rect 10924 3834 10948 3836
rect 11004 3834 11028 3836
rect 11084 3834 11090 3836
rect 10844 3782 10846 3834
rect 11026 3782 11028 3834
rect 10782 3780 10788 3782
rect 10844 3780 10868 3782
rect 10924 3780 10948 3782
rect 11004 3780 11028 3782
rect 11084 3780 11090 3782
rect 10782 3771 11090 3780
rect 11348 3534 11376 4422
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11072 3194 11100 3470
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11716 3058 11744 3878
rect 11992 3058 12020 3878
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12268 2774 12296 5646
rect 12748 5468 13056 5477
rect 12748 5466 12754 5468
rect 12810 5466 12834 5468
rect 12890 5466 12914 5468
rect 12970 5466 12994 5468
rect 13050 5466 13056 5468
rect 12810 5414 12812 5466
rect 12992 5414 12994 5466
rect 12748 5412 12754 5414
rect 12810 5412 12834 5414
rect 12890 5412 12914 5414
rect 12970 5412 12994 5414
rect 13050 5412 13056 5414
rect 12748 5403 13056 5412
rect 13372 4622 13400 6734
rect 14200 4690 14228 6886
rect 14292 6866 14320 7142
rect 14715 7100 15023 7109
rect 14715 7098 14721 7100
rect 14777 7098 14801 7100
rect 14857 7098 14881 7100
rect 14937 7098 14961 7100
rect 15017 7098 15023 7100
rect 14777 7046 14779 7098
rect 14959 7046 14961 7098
rect 14715 7044 14721 7046
rect 14777 7044 14801 7046
rect 14857 7044 14881 7046
rect 14937 7044 14961 7046
rect 15017 7044 15023 7046
rect 14715 7035 15023 7044
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6390 14412 6598
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14568 6322 14596 6666
rect 15396 6322 15424 7346
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15856 6458 15884 6666
rect 16681 6556 16989 6565
rect 16681 6554 16687 6556
rect 16743 6554 16767 6556
rect 16823 6554 16847 6556
rect 16903 6554 16927 6556
rect 16983 6554 16989 6556
rect 16743 6502 16745 6554
rect 16925 6502 16927 6554
rect 16681 6500 16687 6502
rect 16743 6500 16767 6502
rect 16823 6500 16847 6502
rect 16903 6500 16927 6502
rect 16983 6500 16989 6502
rect 16681 6491 16989 6500
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12360 4146 12388 4558
rect 12748 4380 13056 4389
rect 12748 4378 12754 4380
rect 12810 4378 12834 4380
rect 12890 4378 12914 4380
rect 12970 4378 12994 4380
rect 13050 4378 13056 4380
rect 12810 4326 12812 4378
rect 12992 4326 12994 4378
rect 12748 4324 12754 4326
rect 12810 4324 12834 4326
rect 12890 4324 12914 4326
rect 12970 4324 12994 4326
rect 13050 4324 13056 4326
rect 12748 4315 13056 4324
rect 13372 4214 13400 4558
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12912 3738 12940 3946
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 12748 3292 13056 3301
rect 12748 3290 12754 3292
rect 12810 3290 12834 3292
rect 12890 3290 12914 3292
rect 12970 3290 12994 3292
rect 13050 3290 13056 3292
rect 12810 3238 12812 3290
rect 12992 3238 12994 3290
rect 12748 3236 12754 3238
rect 12810 3236 12834 3238
rect 12890 3236 12914 3238
rect 12970 3236 12994 3238
rect 13050 3236 13056 3238
rect 12748 3227 13056 3236
rect 13280 2854 13308 3334
rect 13372 3194 13400 3538
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 10782 2748 11090 2757
rect 10782 2746 10788 2748
rect 10844 2746 10868 2748
rect 10924 2746 10948 2748
rect 11004 2746 11028 2748
rect 11084 2746 11090 2748
rect 12268 2746 12388 2774
rect 10844 2694 10846 2746
rect 11026 2694 11028 2746
rect 10782 2692 10788 2694
rect 10844 2692 10868 2694
rect 10924 2692 10948 2694
rect 11004 2692 11028 2694
rect 11084 2692 11090 2694
rect 10782 2683 11090 2692
rect 12360 2446 12388 2746
rect 13372 2446 13400 3130
rect 13464 2922 13492 4490
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 4146 13952 4422
rect 14200 4282 14228 4626
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3194 14320 3878
rect 14384 3738 14412 4490
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14384 3126 14412 3674
rect 14476 3602 14504 6122
rect 14568 5914 14596 6258
rect 14715 6012 15023 6021
rect 14715 6010 14721 6012
rect 14777 6010 14801 6012
rect 14857 6010 14881 6012
rect 14937 6010 14961 6012
rect 15017 6010 15023 6012
rect 14777 5958 14779 6010
rect 14959 5958 14961 6010
rect 14715 5956 14721 5958
rect 14777 5956 14801 5958
rect 14857 5956 14881 5958
rect 14937 5956 14961 5958
rect 15017 5956 15023 5958
rect 14715 5947 15023 5956
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 16681 5468 16989 5477
rect 16681 5466 16687 5468
rect 16743 5466 16767 5468
rect 16823 5466 16847 5468
rect 16903 5466 16927 5468
rect 16983 5466 16989 5468
rect 16743 5414 16745 5466
rect 16925 5414 16927 5466
rect 16681 5412 16687 5414
rect 16743 5412 16767 5414
rect 16823 5412 16847 5414
rect 16903 5412 16927 5414
rect 16983 5412 16989 5414
rect 16681 5403 16989 5412
rect 14715 4924 15023 4933
rect 14715 4922 14721 4924
rect 14777 4922 14801 4924
rect 14857 4922 14881 4924
rect 14937 4922 14961 4924
rect 15017 4922 15023 4924
rect 14777 4870 14779 4922
rect 14959 4870 14961 4922
rect 14715 4868 14721 4870
rect 14777 4868 14801 4870
rect 14857 4868 14881 4870
rect 14937 4868 14961 4870
rect 15017 4868 15023 4870
rect 14715 4859 15023 4868
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 14384 2446 14412 3062
rect 14476 2990 14504 3538
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14476 2514 14504 2926
rect 14568 2650 14596 4694
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14715 3836 15023 3845
rect 14715 3834 14721 3836
rect 14777 3834 14801 3836
rect 14857 3834 14881 3836
rect 14937 3834 14961 3836
rect 15017 3834 15023 3836
rect 14777 3782 14779 3834
rect 14959 3782 14961 3834
rect 14715 3780 14721 3782
rect 14777 3780 14801 3782
rect 14857 3780 14881 3782
rect 14937 3780 14961 3782
rect 15017 3780 15023 3782
rect 14715 3771 15023 3780
rect 15120 3058 15148 3878
rect 15396 3534 15424 4422
rect 15580 3534 15608 4558
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16681 4380 16989 4389
rect 16681 4378 16687 4380
rect 16743 4378 16767 4380
rect 16823 4378 16847 4380
rect 16903 4378 16927 4380
rect 16983 4378 16989 4380
rect 16743 4326 16745 4378
rect 16925 4326 16927 4378
rect 16681 4324 16687 4326
rect 16743 4324 16767 4326
rect 16823 4324 16847 4326
rect 16903 4324 16927 4326
rect 16983 4324 16989 4326
rect 16681 4315 16989 4324
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 14715 2748 15023 2757
rect 14715 2746 14721 2748
rect 14777 2746 14801 2748
rect 14857 2746 14881 2748
rect 14937 2746 14961 2748
rect 15017 2746 15023 2748
rect 14777 2694 14779 2746
rect 14959 2694 14961 2746
rect 14715 2692 14721 2694
rect 14777 2692 14801 2694
rect 14857 2692 14881 2694
rect 14937 2692 14961 2694
rect 15017 2692 15023 2694
rect 14715 2683 15023 2692
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15120 2446 15148 2994
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2854 15240 2926
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2446 15240 2790
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 848 944 900 950
rect 848 886 900 892
rect 1768 944 1820 950
rect 1768 886 1820 892
rect 860 800 888 886
rect 2332 800 2360 2314
rect 3804 870 3924 898
rect 3804 800 3832 870
rect 846 0 902 800
rect 2318 0 2374 800
rect 3790 0 3846 800
rect 3896 762 3924 870
rect 4172 762 4200 2314
rect 4882 2204 5190 2213
rect 4882 2202 4888 2204
rect 4944 2202 4968 2204
rect 5024 2202 5048 2204
rect 5104 2202 5128 2204
rect 5184 2202 5190 2204
rect 4944 2150 4946 2202
rect 5126 2150 5128 2202
rect 4882 2148 4888 2150
rect 4944 2148 4968 2150
rect 5024 2148 5048 2150
rect 5104 2148 5128 2150
rect 5184 2148 5190 2150
rect 4882 2139 5190 2148
rect 5552 898 5580 2314
rect 6932 898 6960 2314
rect 8312 898 8340 2314
rect 8815 2204 9123 2213
rect 8815 2202 8821 2204
rect 8877 2202 8901 2204
rect 8957 2202 8981 2204
rect 9037 2202 9061 2204
rect 9117 2202 9123 2204
rect 8877 2150 8879 2202
rect 9059 2150 9061 2202
rect 8815 2148 8821 2150
rect 8877 2148 8901 2150
rect 8957 2148 8981 2150
rect 9037 2148 9061 2150
rect 9117 2148 9123 2150
rect 8815 2139 9123 2148
rect 5276 870 5580 898
rect 6748 870 6960 898
rect 8220 870 8340 898
rect 5276 800 5304 870
rect 6748 800 6776 870
rect 8220 800 8248 870
rect 9692 800 9720 2314
rect 11164 800 11192 2314
rect 12636 800 12664 2314
rect 12748 2204 13056 2213
rect 12748 2202 12754 2204
rect 12810 2202 12834 2204
rect 12890 2202 12914 2204
rect 12970 2202 12994 2204
rect 13050 2202 13056 2204
rect 12810 2150 12812 2202
rect 12992 2150 12994 2202
rect 12748 2148 12754 2150
rect 12810 2148 12834 2150
rect 12890 2148 12914 2150
rect 12970 2148 12994 2150
rect 13050 2148 13056 2150
rect 12748 2139 13056 2148
rect 15672 2122 15700 4014
rect 16681 3292 16989 3301
rect 16681 3290 16687 3292
rect 16743 3290 16767 3292
rect 16823 3290 16847 3292
rect 16903 3290 16927 3292
rect 16983 3290 16989 3292
rect 16743 3238 16745 3290
rect 16925 3238 16927 3290
rect 16681 3236 16687 3238
rect 16743 3236 16767 3238
rect 16823 3236 16847 3238
rect 16903 3236 16927 3238
rect 16983 3236 16989 3238
rect 16681 3227 16989 3236
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15580 2094 15700 2122
rect 14096 944 14148 950
rect 14096 886 14148 892
rect 14108 800 14136 886
rect 15580 800 15608 2094
rect 15948 950 15976 2314
rect 16681 2204 16989 2213
rect 16681 2202 16687 2204
rect 16743 2202 16767 2204
rect 16823 2202 16847 2204
rect 16903 2202 16927 2204
rect 16983 2202 16989 2204
rect 16743 2150 16745 2202
rect 16925 2150 16927 2202
rect 16681 2148 16687 2150
rect 16743 2148 16767 2150
rect 16823 2148 16847 2150
rect 16903 2148 16927 2150
rect 16983 2148 16989 2150
rect 16681 2139 16989 2148
rect 15936 944 15988 950
rect 15936 886 15988 892
rect 17052 800 17080 4490
rect 3896 734 4200 762
rect 5262 0 5318 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 14094 0 14150 800
rect 15566 0 15622 800
rect 17038 0 17094 800
<< via2 >>
rect 2922 15802 2978 15804
rect 3002 15802 3058 15804
rect 3082 15802 3138 15804
rect 3162 15802 3218 15804
rect 2922 15750 2968 15802
rect 2968 15750 2978 15802
rect 3002 15750 3032 15802
rect 3032 15750 3044 15802
rect 3044 15750 3058 15802
rect 3082 15750 3096 15802
rect 3096 15750 3108 15802
rect 3108 15750 3138 15802
rect 3162 15750 3172 15802
rect 3172 15750 3218 15802
rect 2922 15748 2978 15750
rect 3002 15748 3058 15750
rect 3082 15748 3138 15750
rect 3162 15748 3218 15750
rect 2922 14714 2978 14716
rect 3002 14714 3058 14716
rect 3082 14714 3138 14716
rect 3162 14714 3218 14716
rect 2922 14662 2968 14714
rect 2968 14662 2978 14714
rect 3002 14662 3032 14714
rect 3032 14662 3044 14714
rect 3044 14662 3058 14714
rect 3082 14662 3096 14714
rect 3096 14662 3108 14714
rect 3108 14662 3138 14714
rect 3162 14662 3172 14714
rect 3172 14662 3218 14714
rect 2922 14660 2978 14662
rect 3002 14660 3058 14662
rect 3082 14660 3138 14662
rect 3162 14660 3218 14662
rect 2922 13626 2978 13628
rect 3002 13626 3058 13628
rect 3082 13626 3138 13628
rect 3162 13626 3218 13628
rect 2922 13574 2968 13626
rect 2968 13574 2978 13626
rect 3002 13574 3032 13626
rect 3032 13574 3044 13626
rect 3044 13574 3058 13626
rect 3082 13574 3096 13626
rect 3096 13574 3108 13626
rect 3108 13574 3138 13626
rect 3162 13574 3172 13626
rect 3172 13574 3218 13626
rect 2922 13572 2978 13574
rect 3002 13572 3058 13574
rect 3082 13572 3138 13574
rect 3162 13572 3218 13574
rect 2922 12538 2978 12540
rect 3002 12538 3058 12540
rect 3082 12538 3138 12540
rect 3162 12538 3218 12540
rect 2922 12486 2968 12538
rect 2968 12486 2978 12538
rect 3002 12486 3032 12538
rect 3032 12486 3044 12538
rect 3044 12486 3058 12538
rect 3082 12486 3096 12538
rect 3096 12486 3108 12538
rect 3108 12486 3138 12538
rect 3162 12486 3172 12538
rect 3172 12486 3218 12538
rect 2922 12484 2978 12486
rect 3002 12484 3058 12486
rect 3082 12484 3138 12486
rect 3162 12484 3218 12486
rect 6855 15802 6911 15804
rect 6935 15802 6991 15804
rect 7015 15802 7071 15804
rect 7095 15802 7151 15804
rect 6855 15750 6901 15802
rect 6901 15750 6911 15802
rect 6935 15750 6965 15802
rect 6965 15750 6977 15802
rect 6977 15750 6991 15802
rect 7015 15750 7029 15802
rect 7029 15750 7041 15802
rect 7041 15750 7071 15802
rect 7095 15750 7105 15802
rect 7105 15750 7151 15802
rect 6855 15748 6911 15750
rect 6935 15748 6991 15750
rect 7015 15748 7071 15750
rect 7095 15748 7151 15750
rect 10788 15802 10844 15804
rect 10868 15802 10924 15804
rect 10948 15802 11004 15804
rect 11028 15802 11084 15804
rect 10788 15750 10834 15802
rect 10834 15750 10844 15802
rect 10868 15750 10898 15802
rect 10898 15750 10910 15802
rect 10910 15750 10924 15802
rect 10948 15750 10962 15802
rect 10962 15750 10974 15802
rect 10974 15750 11004 15802
rect 11028 15750 11038 15802
rect 11038 15750 11084 15802
rect 10788 15748 10844 15750
rect 10868 15748 10924 15750
rect 10948 15748 11004 15750
rect 11028 15748 11084 15750
rect 14721 15802 14777 15804
rect 14801 15802 14857 15804
rect 14881 15802 14937 15804
rect 14961 15802 15017 15804
rect 14721 15750 14767 15802
rect 14767 15750 14777 15802
rect 14801 15750 14831 15802
rect 14831 15750 14843 15802
rect 14843 15750 14857 15802
rect 14881 15750 14895 15802
rect 14895 15750 14907 15802
rect 14907 15750 14937 15802
rect 14961 15750 14971 15802
rect 14971 15750 15017 15802
rect 14721 15748 14777 15750
rect 14801 15748 14857 15750
rect 14881 15748 14937 15750
rect 14961 15748 15017 15750
rect 4888 15258 4944 15260
rect 4968 15258 5024 15260
rect 5048 15258 5104 15260
rect 5128 15258 5184 15260
rect 4888 15206 4934 15258
rect 4934 15206 4944 15258
rect 4968 15206 4998 15258
rect 4998 15206 5010 15258
rect 5010 15206 5024 15258
rect 5048 15206 5062 15258
rect 5062 15206 5074 15258
rect 5074 15206 5104 15258
rect 5128 15206 5138 15258
rect 5138 15206 5184 15258
rect 4888 15204 4944 15206
rect 4968 15204 5024 15206
rect 5048 15204 5104 15206
rect 5128 15204 5184 15206
rect 4888 14170 4944 14172
rect 4968 14170 5024 14172
rect 5048 14170 5104 14172
rect 5128 14170 5184 14172
rect 4888 14118 4934 14170
rect 4934 14118 4944 14170
rect 4968 14118 4998 14170
rect 4998 14118 5010 14170
rect 5010 14118 5024 14170
rect 5048 14118 5062 14170
rect 5062 14118 5074 14170
rect 5074 14118 5104 14170
rect 5128 14118 5138 14170
rect 5138 14118 5184 14170
rect 4888 14116 4944 14118
rect 4968 14116 5024 14118
rect 5048 14116 5104 14118
rect 5128 14116 5184 14118
rect 2922 11450 2978 11452
rect 3002 11450 3058 11452
rect 3082 11450 3138 11452
rect 3162 11450 3218 11452
rect 2922 11398 2968 11450
rect 2968 11398 2978 11450
rect 3002 11398 3032 11450
rect 3032 11398 3044 11450
rect 3044 11398 3058 11450
rect 3082 11398 3096 11450
rect 3096 11398 3108 11450
rect 3108 11398 3138 11450
rect 3162 11398 3172 11450
rect 3172 11398 3218 11450
rect 2922 11396 2978 11398
rect 3002 11396 3058 11398
rect 3082 11396 3138 11398
rect 3162 11396 3218 11398
rect 2922 10362 2978 10364
rect 3002 10362 3058 10364
rect 3082 10362 3138 10364
rect 3162 10362 3218 10364
rect 2922 10310 2968 10362
rect 2968 10310 2978 10362
rect 3002 10310 3032 10362
rect 3032 10310 3044 10362
rect 3044 10310 3058 10362
rect 3082 10310 3096 10362
rect 3096 10310 3108 10362
rect 3108 10310 3138 10362
rect 3162 10310 3172 10362
rect 3172 10310 3218 10362
rect 2922 10308 2978 10310
rect 3002 10308 3058 10310
rect 3082 10308 3138 10310
rect 3162 10308 3218 10310
rect 2922 9274 2978 9276
rect 3002 9274 3058 9276
rect 3082 9274 3138 9276
rect 3162 9274 3218 9276
rect 2922 9222 2968 9274
rect 2968 9222 2978 9274
rect 3002 9222 3032 9274
rect 3032 9222 3044 9274
rect 3044 9222 3058 9274
rect 3082 9222 3096 9274
rect 3096 9222 3108 9274
rect 3108 9222 3138 9274
rect 3162 9222 3172 9274
rect 3172 9222 3218 9274
rect 2922 9220 2978 9222
rect 3002 9220 3058 9222
rect 3082 9220 3138 9222
rect 3162 9220 3218 9222
rect 2922 8186 2978 8188
rect 3002 8186 3058 8188
rect 3082 8186 3138 8188
rect 3162 8186 3218 8188
rect 2922 8134 2968 8186
rect 2968 8134 2978 8186
rect 3002 8134 3032 8186
rect 3032 8134 3044 8186
rect 3044 8134 3058 8186
rect 3082 8134 3096 8186
rect 3096 8134 3108 8186
rect 3108 8134 3138 8186
rect 3162 8134 3172 8186
rect 3172 8134 3218 8186
rect 2922 8132 2978 8134
rect 3002 8132 3058 8134
rect 3082 8132 3138 8134
rect 3162 8132 3218 8134
rect 2922 7098 2978 7100
rect 3002 7098 3058 7100
rect 3082 7098 3138 7100
rect 3162 7098 3218 7100
rect 2922 7046 2968 7098
rect 2968 7046 2978 7098
rect 3002 7046 3032 7098
rect 3032 7046 3044 7098
rect 3044 7046 3058 7098
rect 3082 7046 3096 7098
rect 3096 7046 3108 7098
rect 3108 7046 3138 7098
rect 3162 7046 3172 7098
rect 3172 7046 3218 7098
rect 2922 7044 2978 7046
rect 3002 7044 3058 7046
rect 3082 7044 3138 7046
rect 3162 7044 3218 7046
rect 2922 6010 2978 6012
rect 3002 6010 3058 6012
rect 3082 6010 3138 6012
rect 3162 6010 3218 6012
rect 2922 5958 2968 6010
rect 2968 5958 2978 6010
rect 3002 5958 3032 6010
rect 3032 5958 3044 6010
rect 3044 5958 3058 6010
rect 3082 5958 3096 6010
rect 3096 5958 3108 6010
rect 3108 5958 3138 6010
rect 3162 5958 3172 6010
rect 3172 5958 3218 6010
rect 2922 5956 2978 5958
rect 3002 5956 3058 5958
rect 3082 5956 3138 5958
rect 3162 5956 3218 5958
rect 8821 15258 8877 15260
rect 8901 15258 8957 15260
rect 8981 15258 9037 15260
rect 9061 15258 9117 15260
rect 8821 15206 8867 15258
rect 8867 15206 8877 15258
rect 8901 15206 8931 15258
rect 8931 15206 8943 15258
rect 8943 15206 8957 15258
rect 8981 15206 8995 15258
rect 8995 15206 9007 15258
rect 9007 15206 9037 15258
rect 9061 15206 9071 15258
rect 9071 15206 9117 15258
rect 8821 15204 8877 15206
rect 8901 15204 8957 15206
rect 8981 15204 9037 15206
rect 9061 15204 9117 15206
rect 6855 14714 6911 14716
rect 6935 14714 6991 14716
rect 7015 14714 7071 14716
rect 7095 14714 7151 14716
rect 6855 14662 6901 14714
rect 6901 14662 6911 14714
rect 6935 14662 6965 14714
rect 6965 14662 6977 14714
rect 6977 14662 6991 14714
rect 7015 14662 7029 14714
rect 7029 14662 7041 14714
rect 7041 14662 7071 14714
rect 7095 14662 7105 14714
rect 7105 14662 7151 14714
rect 6855 14660 6911 14662
rect 6935 14660 6991 14662
rect 7015 14660 7071 14662
rect 7095 14660 7151 14662
rect 4888 13082 4944 13084
rect 4968 13082 5024 13084
rect 5048 13082 5104 13084
rect 5128 13082 5184 13084
rect 4888 13030 4934 13082
rect 4934 13030 4944 13082
rect 4968 13030 4998 13082
rect 4998 13030 5010 13082
rect 5010 13030 5024 13082
rect 5048 13030 5062 13082
rect 5062 13030 5074 13082
rect 5074 13030 5104 13082
rect 5128 13030 5138 13082
rect 5138 13030 5184 13082
rect 4888 13028 4944 13030
rect 4968 13028 5024 13030
rect 5048 13028 5104 13030
rect 5128 13028 5184 13030
rect 4888 11994 4944 11996
rect 4968 11994 5024 11996
rect 5048 11994 5104 11996
rect 5128 11994 5184 11996
rect 4888 11942 4934 11994
rect 4934 11942 4944 11994
rect 4968 11942 4998 11994
rect 4998 11942 5010 11994
rect 5010 11942 5024 11994
rect 5048 11942 5062 11994
rect 5062 11942 5074 11994
rect 5074 11942 5104 11994
rect 5128 11942 5138 11994
rect 5138 11942 5184 11994
rect 4888 11940 4944 11942
rect 4968 11940 5024 11942
rect 5048 11940 5104 11942
rect 5128 11940 5184 11942
rect 4888 10906 4944 10908
rect 4968 10906 5024 10908
rect 5048 10906 5104 10908
rect 5128 10906 5184 10908
rect 4888 10854 4934 10906
rect 4934 10854 4944 10906
rect 4968 10854 4998 10906
rect 4998 10854 5010 10906
rect 5010 10854 5024 10906
rect 5048 10854 5062 10906
rect 5062 10854 5074 10906
rect 5074 10854 5104 10906
rect 5128 10854 5138 10906
rect 5138 10854 5184 10906
rect 4888 10852 4944 10854
rect 4968 10852 5024 10854
rect 5048 10852 5104 10854
rect 5128 10852 5184 10854
rect 4888 9818 4944 9820
rect 4968 9818 5024 9820
rect 5048 9818 5104 9820
rect 5128 9818 5184 9820
rect 4888 9766 4934 9818
rect 4934 9766 4944 9818
rect 4968 9766 4998 9818
rect 4998 9766 5010 9818
rect 5010 9766 5024 9818
rect 5048 9766 5062 9818
rect 5062 9766 5074 9818
rect 5074 9766 5104 9818
rect 5128 9766 5138 9818
rect 5138 9766 5184 9818
rect 4888 9764 4944 9766
rect 4968 9764 5024 9766
rect 5048 9764 5104 9766
rect 5128 9764 5184 9766
rect 6855 13626 6911 13628
rect 6935 13626 6991 13628
rect 7015 13626 7071 13628
rect 7095 13626 7151 13628
rect 6855 13574 6901 13626
rect 6901 13574 6911 13626
rect 6935 13574 6965 13626
rect 6965 13574 6977 13626
rect 6977 13574 6991 13626
rect 7015 13574 7029 13626
rect 7029 13574 7041 13626
rect 7041 13574 7071 13626
rect 7095 13574 7105 13626
rect 7105 13574 7151 13626
rect 6855 13572 6911 13574
rect 6935 13572 6991 13574
rect 7015 13572 7071 13574
rect 7095 13572 7151 13574
rect 6855 12538 6911 12540
rect 6935 12538 6991 12540
rect 7015 12538 7071 12540
rect 7095 12538 7151 12540
rect 6855 12486 6901 12538
rect 6901 12486 6911 12538
rect 6935 12486 6965 12538
rect 6965 12486 6977 12538
rect 6977 12486 6991 12538
rect 7015 12486 7029 12538
rect 7029 12486 7041 12538
rect 7041 12486 7071 12538
rect 7095 12486 7105 12538
rect 7105 12486 7151 12538
rect 6855 12484 6911 12486
rect 6935 12484 6991 12486
rect 7015 12484 7071 12486
rect 7095 12484 7151 12486
rect 4888 8730 4944 8732
rect 4968 8730 5024 8732
rect 5048 8730 5104 8732
rect 5128 8730 5184 8732
rect 4888 8678 4934 8730
rect 4934 8678 4944 8730
rect 4968 8678 4998 8730
rect 4998 8678 5010 8730
rect 5010 8678 5024 8730
rect 5048 8678 5062 8730
rect 5062 8678 5074 8730
rect 5074 8678 5104 8730
rect 5128 8678 5138 8730
rect 5138 8678 5184 8730
rect 4888 8676 4944 8678
rect 4968 8676 5024 8678
rect 5048 8676 5104 8678
rect 5128 8676 5184 8678
rect 4888 7642 4944 7644
rect 4968 7642 5024 7644
rect 5048 7642 5104 7644
rect 5128 7642 5184 7644
rect 4888 7590 4934 7642
rect 4934 7590 4944 7642
rect 4968 7590 4998 7642
rect 4998 7590 5010 7642
rect 5010 7590 5024 7642
rect 5048 7590 5062 7642
rect 5062 7590 5074 7642
rect 5074 7590 5104 7642
rect 5128 7590 5138 7642
rect 5138 7590 5184 7642
rect 4888 7588 4944 7590
rect 4968 7588 5024 7590
rect 5048 7588 5104 7590
rect 5128 7588 5184 7590
rect 4888 6554 4944 6556
rect 4968 6554 5024 6556
rect 5048 6554 5104 6556
rect 5128 6554 5184 6556
rect 4888 6502 4934 6554
rect 4934 6502 4944 6554
rect 4968 6502 4998 6554
rect 4998 6502 5010 6554
rect 5010 6502 5024 6554
rect 5048 6502 5062 6554
rect 5062 6502 5074 6554
rect 5074 6502 5104 6554
rect 5128 6502 5138 6554
rect 5138 6502 5184 6554
rect 4888 6500 4944 6502
rect 4968 6500 5024 6502
rect 5048 6500 5104 6502
rect 5128 6500 5184 6502
rect 4888 5466 4944 5468
rect 4968 5466 5024 5468
rect 5048 5466 5104 5468
rect 5128 5466 5184 5468
rect 4888 5414 4934 5466
rect 4934 5414 4944 5466
rect 4968 5414 4998 5466
rect 4998 5414 5010 5466
rect 5010 5414 5024 5466
rect 5048 5414 5062 5466
rect 5062 5414 5074 5466
rect 5074 5414 5104 5466
rect 5128 5414 5138 5466
rect 5138 5414 5184 5466
rect 4888 5412 4944 5414
rect 4968 5412 5024 5414
rect 5048 5412 5104 5414
rect 5128 5412 5184 5414
rect 2922 4922 2978 4924
rect 3002 4922 3058 4924
rect 3082 4922 3138 4924
rect 3162 4922 3218 4924
rect 2922 4870 2968 4922
rect 2968 4870 2978 4922
rect 3002 4870 3032 4922
rect 3032 4870 3044 4922
rect 3044 4870 3058 4922
rect 3082 4870 3096 4922
rect 3096 4870 3108 4922
rect 3108 4870 3138 4922
rect 3162 4870 3172 4922
rect 3172 4870 3218 4922
rect 2922 4868 2978 4870
rect 3002 4868 3058 4870
rect 3082 4868 3138 4870
rect 3162 4868 3218 4870
rect 2922 3834 2978 3836
rect 3002 3834 3058 3836
rect 3082 3834 3138 3836
rect 3162 3834 3218 3836
rect 2922 3782 2968 3834
rect 2968 3782 2978 3834
rect 3002 3782 3032 3834
rect 3032 3782 3044 3834
rect 3044 3782 3058 3834
rect 3082 3782 3096 3834
rect 3096 3782 3108 3834
rect 3108 3782 3138 3834
rect 3162 3782 3172 3834
rect 3172 3782 3218 3834
rect 2922 3780 2978 3782
rect 3002 3780 3058 3782
rect 3082 3780 3138 3782
rect 3162 3780 3218 3782
rect 2922 2746 2978 2748
rect 3002 2746 3058 2748
rect 3082 2746 3138 2748
rect 3162 2746 3218 2748
rect 2922 2694 2968 2746
rect 2968 2694 2978 2746
rect 3002 2694 3032 2746
rect 3032 2694 3044 2746
rect 3044 2694 3058 2746
rect 3082 2694 3096 2746
rect 3096 2694 3108 2746
rect 3108 2694 3138 2746
rect 3162 2694 3172 2746
rect 3172 2694 3218 2746
rect 2922 2692 2978 2694
rect 3002 2692 3058 2694
rect 3082 2692 3138 2694
rect 3162 2692 3218 2694
rect 4888 4378 4944 4380
rect 4968 4378 5024 4380
rect 5048 4378 5104 4380
rect 5128 4378 5184 4380
rect 4888 4326 4934 4378
rect 4934 4326 4944 4378
rect 4968 4326 4998 4378
rect 4998 4326 5010 4378
rect 5010 4326 5024 4378
rect 5048 4326 5062 4378
rect 5062 4326 5074 4378
rect 5074 4326 5104 4378
rect 5128 4326 5138 4378
rect 5138 4326 5184 4378
rect 4888 4324 4944 4326
rect 4968 4324 5024 4326
rect 5048 4324 5104 4326
rect 5128 4324 5184 4326
rect 4888 3290 4944 3292
rect 4968 3290 5024 3292
rect 5048 3290 5104 3292
rect 5128 3290 5184 3292
rect 4888 3238 4934 3290
rect 4934 3238 4944 3290
rect 4968 3238 4998 3290
rect 4998 3238 5010 3290
rect 5010 3238 5024 3290
rect 5048 3238 5062 3290
rect 5062 3238 5074 3290
rect 5074 3238 5104 3290
rect 5128 3238 5138 3290
rect 5138 3238 5184 3290
rect 4888 3236 4944 3238
rect 4968 3236 5024 3238
rect 5048 3236 5104 3238
rect 5128 3236 5184 3238
rect 6855 11450 6911 11452
rect 6935 11450 6991 11452
rect 7015 11450 7071 11452
rect 7095 11450 7151 11452
rect 6855 11398 6901 11450
rect 6901 11398 6911 11450
rect 6935 11398 6965 11450
rect 6965 11398 6977 11450
rect 6977 11398 6991 11450
rect 7015 11398 7029 11450
rect 7029 11398 7041 11450
rect 7041 11398 7071 11450
rect 7095 11398 7105 11450
rect 7105 11398 7151 11450
rect 6855 11396 6911 11398
rect 6935 11396 6991 11398
rect 7015 11396 7071 11398
rect 7095 11396 7151 11398
rect 6855 10362 6911 10364
rect 6935 10362 6991 10364
rect 7015 10362 7071 10364
rect 7095 10362 7151 10364
rect 6855 10310 6901 10362
rect 6901 10310 6911 10362
rect 6935 10310 6965 10362
rect 6965 10310 6977 10362
rect 6977 10310 6991 10362
rect 7015 10310 7029 10362
rect 7029 10310 7041 10362
rect 7041 10310 7071 10362
rect 7095 10310 7105 10362
rect 7105 10310 7151 10362
rect 6855 10308 6911 10310
rect 6935 10308 6991 10310
rect 7015 10308 7071 10310
rect 7095 10308 7151 10310
rect 6855 9274 6911 9276
rect 6935 9274 6991 9276
rect 7015 9274 7071 9276
rect 7095 9274 7151 9276
rect 6855 9222 6901 9274
rect 6901 9222 6911 9274
rect 6935 9222 6965 9274
rect 6965 9222 6977 9274
rect 6977 9222 6991 9274
rect 7015 9222 7029 9274
rect 7029 9222 7041 9274
rect 7041 9222 7071 9274
rect 7095 9222 7105 9274
rect 7105 9222 7151 9274
rect 6855 9220 6911 9222
rect 6935 9220 6991 9222
rect 7015 9220 7071 9222
rect 7095 9220 7151 9222
rect 6855 8186 6911 8188
rect 6935 8186 6991 8188
rect 7015 8186 7071 8188
rect 7095 8186 7151 8188
rect 6855 8134 6901 8186
rect 6901 8134 6911 8186
rect 6935 8134 6965 8186
rect 6965 8134 6977 8186
rect 6977 8134 6991 8186
rect 7015 8134 7029 8186
rect 7029 8134 7041 8186
rect 7041 8134 7071 8186
rect 7095 8134 7105 8186
rect 7105 8134 7151 8186
rect 6855 8132 6911 8134
rect 6935 8132 6991 8134
rect 7015 8132 7071 8134
rect 7095 8132 7151 8134
rect 6855 7098 6911 7100
rect 6935 7098 6991 7100
rect 7015 7098 7071 7100
rect 7095 7098 7151 7100
rect 6855 7046 6901 7098
rect 6901 7046 6911 7098
rect 6935 7046 6965 7098
rect 6965 7046 6977 7098
rect 6977 7046 6991 7098
rect 7015 7046 7029 7098
rect 7029 7046 7041 7098
rect 7041 7046 7071 7098
rect 7095 7046 7105 7098
rect 7105 7046 7151 7098
rect 6855 7044 6911 7046
rect 6935 7044 6991 7046
rect 7015 7044 7071 7046
rect 7095 7044 7151 7046
rect 6855 6010 6911 6012
rect 6935 6010 6991 6012
rect 7015 6010 7071 6012
rect 7095 6010 7151 6012
rect 6855 5958 6901 6010
rect 6901 5958 6911 6010
rect 6935 5958 6965 6010
rect 6965 5958 6977 6010
rect 6977 5958 6991 6010
rect 7015 5958 7029 6010
rect 7029 5958 7041 6010
rect 7041 5958 7071 6010
rect 7095 5958 7105 6010
rect 7105 5958 7151 6010
rect 6855 5956 6911 5958
rect 6935 5956 6991 5958
rect 7015 5956 7071 5958
rect 7095 5956 7151 5958
rect 6855 4922 6911 4924
rect 6935 4922 6991 4924
rect 7015 4922 7071 4924
rect 7095 4922 7151 4924
rect 6855 4870 6901 4922
rect 6901 4870 6911 4922
rect 6935 4870 6965 4922
rect 6965 4870 6977 4922
rect 6977 4870 6991 4922
rect 7015 4870 7029 4922
rect 7029 4870 7041 4922
rect 7041 4870 7071 4922
rect 7095 4870 7105 4922
rect 7105 4870 7151 4922
rect 6855 4868 6911 4870
rect 6935 4868 6991 4870
rect 7015 4868 7071 4870
rect 7095 4868 7151 4870
rect 8821 14170 8877 14172
rect 8901 14170 8957 14172
rect 8981 14170 9037 14172
rect 9061 14170 9117 14172
rect 8821 14118 8867 14170
rect 8867 14118 8877 14170
rect 8901 14118 8931 14170
rect 8931 14118 8943 14170
rect 8943 14118 8957 14170
rect 8981 14118 8995 14170
rect 8995 14118 9007 14170
rect 9007 14118 9037 14170
rect 9061 14118 9071 14170
rect 9071 14118 9117 14170
rect 8821 14116 8877 14118
rect 8901 14116 8957 14118
rect 8981 14116 9037 14118
rect 9061 14116 9117 14118
rect 8821 13082 8877 13084
rect 8901 13082 8957 13084
rect 8981 13082 9037 13084
rect 9061 13082 9117 13084
rect 8821 13030 8867 13082
rect 8867 13030 8877 13082
rect 8901 13030 8931 13082
rect 8931 13030 8943 13082
rect 8943 13030 8957 13082
rect 8981 13030 8995 13082
rect 8995 13030 9007 13082
rect 9007 13030 9037 13082
rect 9061 13030 9071 13082
rect 9071 13030 9117 13082
rect 8821 13028 8877 13030
rect 8901 13028 8957 13030
rect 8981 13028 9037 13030
rect 9061 13028 9117 13030
rect 10788 14714 10844 14716
rect 10868 14714 10924 14716
rect 10948 14714 11004 14716
rect 11028 14714 11084 14716
rect 10788 14662 10834 14714
rect 10834 14662 10844 14714
rect 10868 14662 10898 14714
rect 10898 14662 10910 14714
rect 10910 14662 10924 14714
rect 10948 14662 10962 14714
rect 10962 14662 10974 14714
rect 10974 14662 11004 14714
rect 11028 14662 11038 14714
rect 11038 14662 11084 14714
rect 10788 14660 10844 14662
rect 10868 14660 10924 14662
rect 10948 14660 11004 14662
rect 11028 14660 11084 14662
rect 12754 15258 12810 15260
rect 12834 15258 12890 15260
rect 12914 15258 12970 15260
rect 12994 15258 13050 15260
rect 12754 15206 12800 15258
rect 12800 15206 12810 15258
rect 12834 15206 12864 15258
rect 12864 15206 12876 15258
rect 12876 15206 12890 15258
rect 12914 15206 12928 15258
rect 12928 15206 12940 15258
rect 12940 15206 12970 15258
rect 12994 15206 13004 15258
rect 13004 15206 13050 15258
rect 12754 15204 12810 15206
rect 12834 15204 12890 15206
rect 12914 15204 12970 15206
rect 12994 15204 13050 15206
rect 10788 13626 10844 13628
rect 10868 13626 10924 13628
rect 10948 13626 11004 13628
rect 11028 13626 11084 13628
rect 10788 13574 10834 13626
rect 10834 13574 10844 13626
rect 10868 13574 10898 13626
rect 10898 13574 10910 13626
rect 10910 13574 10924 13626
rect 10948 13574 10962 13626
rect 10962 13574 10974 13626
rect 10974 13574 11004 13626
rect 11028 13574 11038 13626
rect 11038 13574 11084 13626
rect 10788 13572 10844 13574
rect 10868 13572 10924 13574
rect 10948 13572 11004 13574
rect 11028 13572 11084 13574
rect 12754 14170 12810 14172
rect 12834 14170 12890 14172
rect 12914 14170 12970 14172
rect 12994 14170 13050 14172
rect 12754 14118 12800 14170
rect 12800 14118 12810 14170
rect 12834 14118 12864 14170
rect 12864 14118 12876 14170
rect 12876 14118 12890 14170
rect 12914 14118 12928 14170
rect 12928 14118 12940 14170
rect 12940 14118 12970 14170
rect 12994 14118 13004 14170
rect 13004 14118 13050 14170
rect 12754 14116 12810 14118
rect 12834 14116 12890 14118
rect 12914 14116 12970 14118
rect 12994 14116 13050 14118
rect 10788 12538 10844 12540
rect 10868 12538 10924 12540
rect 10948 12538 11004 12540
rect 11028 12538 11084 12540
rect 10788 12486 10834 12538
rect 10834 12486 10844 12538
rect 10868 12486 10898 12538
rect 10898 12486 10910 12538
rect 10910 12486 10924 12538
rect 10948 12486 10962 12538
rect 10962 12486 10974 12538
rect 10974 12486 11004 12538
rect 11028 12486 11038 12538
rect 11038 12486 11084 12538
rect 10788 12484 10844 12486
rect 10868 12484 10924 12486
rect 10948 12484 11004 12486
rect 11028 12484 11084 12486
rect 8821 11994 8877 11996
rect 8901 11994 8957 11996
rect 8981 11994 9037 11996
rect 9061 11994 9117 11996
rect 8821 11942 8867 11994
rect 8867 11942 8877 11994
rect 8901 11942 8931 11994
rect 8931 11942 8943 11994
rect 8943 11942 8957 11994
rect 8981 11942 8995 11994
rect 8995 11942 9007 11994
rect 9007 11942 9037 11994
rect 9061 11942 9071 11994
rect 9071 11942 9117 11994
rect 8821 11940 8877 11942
rect 8901 11940 8957 11942
rect 8981 11940 9037 11942
rect 9061 11940 9117 11942
rect 8821 10906 8877 10908
rect 8901 10906 8957 10908
rect 8981 10906 9037 10908
rect 9061 10906 9117 10908
rect 8821 10854 8867 10906
rect 8867 10854 8877 10906
rect 8901 10854 8931 10906
rect 8931 10854 8943 10906
rect 8943 10854 8957 10906
rect 8981 10854 8995 10906
rect 8995 10854 9007 10906
rect 9007 10854 9037 10906
rect 9061 10854 9071 10906
rect 9071 10854 9117 10906
rect 8821 10852 8877 10854
rect 8901 10852 8957 10854
rect 8981 10852 9037 10854
rect 9061 10852 9117 10854
rect 8821 9818 8877 9820
rect 8901 9818 8957 9820
rect 8981 9818 9037 9820
rect 9061 9818 9117 9820
rect 8821 9766 8867 9818
rect 8867 9766 8877 9818
rect 8901 9766 8931 9818
rect 8931 9766 8943 9818
rect 8943 9766 8957 9818
rect 8981 9766 8995 9818
rect 8995 9766 9007 9818
rect 9007 9766 9037 9818
rect 9061 9766 9071 9818
rect 9071 9766 9117 9818
rect 8821 9764 8877 9766
rect 8901 9764 8957 9766
rect 8981 9764 9037 9766
rect 9061 9764 9117 9766
rect 8821 8730 8877 8732
rect 8901 8730 8957 8732
rect 8981 8730 9037 8732
rect 9061 8730 9117 8732
rect 8821 8678 8867 8730
rect 8867 8678 8877 8730
rect 8901 8678 8931 8730
rect 8931 8678 8943 8730
rect 8943 8678 8957 8730
rect 8981 8678 8995 8730
rect 8995 8678 9007 8730
rect 9007 8678 9037 8730
rect 9061 8678 9071 8730
rect 9071 8678 9117 8730
rect 8821 8676 8877 8678
rect 8901 8676 8957 8678
rect 8981 8676 9037 8678
rect 9061 8676 9117 8678
rect 10788 11450 10844 11452
rect 10868 11450 10924 11452
rect 10948 11450 11004 11452
rect 11028 11450 11084 11452
rect 10788 11398 10834 11450
rect 10834 11398 10844 11450
rect 10868 11398 10898 11450
rect 10898 11398 10910 11450
rect 10910 11398 10924 11450
rect 10948 11398 10962 11450
rect 10962 11398 10974 11450
rect 10974 11398 11004 11450
rect 11028 11398 11038 11450
rect 11038 11398 11084 11450
rect 10788 11396 10844 11398
rect 10868 11396 10924 11398
rect 10948 11396 11004 11398
rect 11028 11396 11084 11398
rect 10788 10362 10844 10364
rect 10868 10362 10924 10364
rect 10948 10362 11004 10364
rect 11028 10362 11084 10364
rect 10788 10310 10834 10362
rect 10834 10310 10844 10362
rect 10868 10310 10898 10362
rect 10898 10310 10910 10362
rect 10910 10310 10924 10362
rect 10948 10310 10962 10362
rect 10962 10310 10974 10362
rect 10974 10310 11004 10362
rect 11028 10310 11038 10362
rect 11038 10310 11084 10362
rect 10788 10308 10844 10310
rect 10868 10308 10924 10310
rect 10948 10308 11004 10310
rect 11028 10308 11084 10310
rect 10788 9274 10844 9276
rect 10868 9274 10924 9276
rect 10948 9274 11004 9276
rect 11028 9274 11084 9276
rect 10788 9222 10834 9274
rect 10834 9222 10844 9274
rect 10868 9222 10898 9274
rect 10898 9222 10910 9274
rect 10910 9222 10924 9274
rect 10948 9222 10962 9274
rect 10962 9222 10974 9274
rect 10974 9222 11004 9274
rect 11028 9222 11038 9274
rect 11038 9222 11084 9274
rect 10788 9220 10844 9222
rect 10868 9220 10924 9222
rect 10948 9220 11004 9222
rect 11028 9220 11084 9222
rect 12754 13082 12810 13084
rect 12834 13082 12890 13084
rect 12914 13082 12970 13084
rect 12994 13082 13050 13084
rect 12754 13030 12800 13082
rect 12800 13030 12810 13082
rect 12834 13030 12864 13082
rect 12864 13030 12876 13082
rect 12876 13030 12890 13082
rect 12914 13030 12928 13082
rect 12928 13030 12940 13082
rect 12940 13030 12970 13082
rect 12994 13030 13004 13082
rect 13004 13030 13050 13082
rect 12754 13028 12810 13030
rect 12834 13028 12890 13030
rect 12914 13028 12970 13030
rect 12994 13028 13050 13030
rect 12754 11994 12810 11996
rect 12834 11994 12890 11996
rect 12914 11994 12970 11996
rect 12994 11994 13050 11996
rect 12754 11942 12800 11994
rect 12800 11942 12810 11994
rect 12834 11942 12864 11994
rect 12864 11942 12876 11994
rect 12876 11942 12890 11994
rect 12914 11942 12928 11994
rect 12928 11942 12940 11994
rect 12940 11942 12970 11994
rect 12994 11942 13004 11994
rect 13004 11942 13050 11994
rect 12754 11940 12810 11942
rect 12834 11940 12890 11942
rect 12914 11940 12970 11942
rect 12994 11940 13050 11942
rect 8821 7642 8877 7644
rect 8901 7642 8957 7644
rect 8981 7642 9037 7644
rect 9061 7642 9117 7644
rect 8821 7590 8867 7642
rect 8867 7590 8877 7642
rect 8901 7590 8931 7642
rect 8931 7590 8943 7642
rect 8943 7590 8957 7642
rect 8981 7590 8995 7642
rect 8995 7590 9007 7642
rect 9007 7590 9037 7642
rect 9061 7590 9071 7642
rect 9071 7590 9117 7642
rect 8821 7588 8877 7590
rect 8901 7588 8957 7590
rect 8981 7588 9037 7590
rect 9061 7588 9117 7590
rect 8821 6554 8877 6556
rect 8901 6554 8957 6556
rect 8981 6554 9037 6556
rect 9061 6554 9117 6556
rect 8821 6502 8867 6554
rect 8867 6502 8877 6554
rect 8901 6502 8931 6554
rect 8931 6502 8943 6554
rect 8943 6502 8957 6554
rect 8981 6502 8995 6554
rect 8995 6502 9007 6554
rect 9007 6502 9037 6554
rect 9061 6502 9071 6554
rect 9071 6502 9117 6554
rect 8821 6500 8877 6502
rect 8901 6500 8957 6502
rect 8981 6500 9037 6502
rect 9061 6500 9117 6502
rect 6855 3834 6911 3836
rect 6935 3834 6991 3836
rect 7015 3834 7071 3836
rect 7095 3834 7151 3836
rect 6855 3782 6901 3834
rect 6901 3782 6911 3834
rect 6935 3782 6965 3834
rect 6965 3782 6977 3834
rect 6977 3782 6991 3834
rect 7015 3782 7029 3834
rect 7029 3782 7041 3834
rect 7041 3782 7071 3834
rect 7095 3782 7105 3834
rect 7105 3782 7151 3834
rect 6855 3780 6911 3782
rect 6935 3780 6991 3782
rect 7015 3780 7071 3782
rect 7095 3780 7151 3782
rect 6855 2746 6911 2748
rect 6935 2746 6991 2748
rect 7015 2746 7071 2748
rect 7095 2746 7151 2748
rect 6855 2694 6901 2746
rect 6901 2694 6911 2746
rect 6935 2694 6965 2746
rect 6965 2694 6977 2746
rect 6977 2694 6991 2746
rect 7015 2694 7029 2746
rect 7029 2694 7041 2746
rect 7041 2694 7071 2746
rect 7095 2694 7105 2746
rect 7105 2694 7151 2746
rect 6855 2692 6911 2694
rect 6935 2692 6991 2694
rect 7015 2692 7071 2694
rect 7095 2692 7151 2694
rect 10788 8186 10844 8188
rect 10868 8186 10924 8188
rect 10948 8186 11004 8188
rect 11028 8186 11084 8188
rect 10788 8134 10834 8186
rect 10834 8134 10844 8186
rect 10868 8134 10898 8186
rect 10898 8134 10910 8186
rect 10910 8134 10924 8186
rect 10948 8134 10962 8186
rect 10962 8134 10974 8186
rect 10974 8134 11004 8186
rect 11028 8134 11038 8186
rect 11038 8134 11084 8186
rect 10788 8132 10844 8134
rect 10868 8132 10924 8134
rect 10948 8132 11004 8134
rect 11028 8132 11084 8134
rect 12754 10906 12810 10908
rect 12834 10906 12890 10908
rect 12914 10906 12970 10908
rect 12994 10906 13050 10908
rect 12754 10854 12800 10906
rect 12800 10854 12810 10906
rect 12834 10854 12864 10906
rect 12864 10854 12876 10906
rect 12876 10854 12890 10906
rect 12914 10854 12928 10906
rect 12928 10854 12940 10906
rect 12940 10854 12970 10906
rect 12994 10854 13004 10906
rect 13004 10854 13050 10906
rect 12754 10852 12810 10854
rect 12834 10852 12890 10854
rect 12914 10852 12970 10854
rect 12994 10852 13050 10854
rect 12754 9818 12810 9820
rect 12834 9818 12890 9820
rect 12914 9818 12970 9820
rect 12994 9818 13050 9820
rect 12754 9766 12800 9818
rect 12800 9766 12810 9818
rect 12834 9766 12864 9818
rect 12864 9766 12876 9818
rect 12876 9766 12890 9818
rect 12914 9766 12928 9818
rect 12928 9766 12940 9818
rect 12940 9766 12970 9818
rect 12994 9766 13004 9818
rect 13004 9766 13050 9818
rect 12754 9764 12810 9766
rect 12834 9764 12890 9766
rect 12914 9764 12970 9766
rect 12994 9764 13050 9766
rect 12754 8730 12810 8732
rect 12834 8730 12890 8732
rect 12914 8730 12970 8732
rect 12994 8730 13050 8732
rect 12754 8678 12800 8730
rect 12800 8678 12810 8730
rect 12834 8678 12864 8730
rect 12864 8678 12876 8730
rect 12876 8678 12890 8730
rect 12914 8678 12928 8730
rect 12928 8678 12940 8730
rect 12940 8678 12970 8730
rect 12994 8678 13004 8730
rect 13004 8678 13050 8730
rect 12754 8676 12810 8678
rect 12834 8676 12890 8678
rect 12914 8676 12970 8678
rect 12994 8676 13050 8678
rect 10788 7098 10844 7100
rect 10868 7098 10924 7100
rect 10948 7098 11004 7100
rect 11028 7098 11084 7100
rect 10788 7046 10834 7098
rect 10834 7046 10844 7098
rect 10868 7046 10898 7098
rect 10898 7046 10910 7098
rect 10910 7046 10924 7098
rect 10948 7046 10962 7098
rect 10962 7046 10974 7098
rect 10974 7046 11004 7098
rect 11028 7046 11038 7098
rect 11038 7046 11084 7098
rect 10788 7044 10844 7046
rect 10868 7044 10924 7046
rect 10948 7044 11004 7046
rect 11028 7044 11084 7046
rect 8821 5466 8877 5468
rect 8901 5466 8957 5468
rect 8981 5466 9037 5468
rect 9061 5466 9117 5468
rect 8821 5414 8867 5466
rect 8867 5414 8877 5466
rect 8901 5414 8931 5466
rect 8931 5414 8943 5466
rect 8943 5414 8957 5466
rect 8981 5414 8995 5466
rect 8995 5414 9007 5466
rect 9007 5414 9037 5466
rect 9061 5414 9071 5466
rect 9071 5414 9117 5466
rect 8821 5412 8877 5414
rect 8901 5412 8957 5414
rect 8981 5412 9037 5414
rect 9061 5412 9117 5414
rect 8821 4378 8877 4380
rect 8901 4378 8957 4380
rect 8981 4378 9037 4380
rect 9061 4378 9117 4380
rect 8821 4326 8867 4378
rect 8867 4326 8877 4378
rect 8901 4326 8931 4378
rect 8931 4326 8943 4378
rect 8943 4326 8957 4378
rect 8981 4326 8995 4378
rect 8995 4326 9007 4378
rect 9007 4326 9037 4378
rect 9061 4326 9071 4378
rect 9071 4326 9117 4378
rect 8821 4324 8877 4326
rect 8901 4324 8957 4326
rect 8981 4324 9037 4326
rect 9061 4324 9117 4326
rect 12754 7642 12810 7644
rect 12834 7642 12890 7644
rect 12914 7642 12970 7644
rect 12994 7642 13050 7644
rect 12754 7590 12800 7642
rect 12800 7590 12810 7642
rect 12834 7590 12864 7642
rect 12864 7590 12876 7642
rect 12876 7590 12890 7642
rect 12914 7590 12928 7642
rect 12928 7590 12940 7642
rect 12940 7590 12970 7642
rect 12994 7590 13004 7642
rect 13004 7590 13050 7642
rect 12754 7588 12810 7590
rect 12834 7588 12890 7590
rect 12914 7588 12970 7590
rect 12994 7588 13050 7590
rect 14721 14714 14777 14716
rect 14801 14714 14857 14716
rect 14881 14714 14937 14716
rect 14961 14714 15017 14716
rect 14721 14662 14767 14714
rect 14767 14662 14777 14714
rect 14801 14662 14831 14714
rect 14831 14662 14843 14714
rect 14843 14662 14857 14714
rect 14881 14662 14895 14714
rect 14895 14662 14907 14714
rect 14907 14662 14937 14714
rect 14961 14662 14971 14714
rect 14971 14662 15017 14714
rect 14721 14660 14777 14662
rect 14801 14660 14857 14662
rect 14881 14660 14937 14662
rect 14961 14660 15017 14662
rect 14721 13626 14777 13628
rect 14801 13626 14857 13628
rect 14881 13626 14937 13628
rect 14961 13626 15017 13628
rect 14721 13574 14767 13626
rect 14767 13574 14777 13626
rect 14801 13574 14831 13626
rect 14831 13574 14843 13626
rect 14843 13574 14857 13626
rect 14881 13574 14895 13626
rect 14895 13574 14907 13626
rect 14907 13574 14937 13626
rect 14961 13574 14971 13626
rect 14971 13574 15017 13626
rect 14721 13572 14777 13574
rect 14801 13572 14857 13574
rect 14881 13572 14937 13574
rect 14961 13572 15017 13574
rect 16687 15258 16743 15260
rect 16767 15258 16823 15260
rect 16847 15258 16903 15260
rect 16927 15258 16983 15260
rect 16687 15206 16733 15258
rect 16733 15206 16743 15258
rect 16767 15206 16797 15258
rect 16797 15206 16809 15258
rect 16809 15206 16823 15258
rect 16847 15206 16861 15258
rect 16861 15206 16873 15258
rect 16873 15206 16903 15258
rect 16927 15206 16937 15258
rect 16937 15206 16983 15258
rect 16687 15204 16743 15206
rect 16767 15204 16823 15206
rect 16847 15204 16903 15206
rect 16927 15204 16983 15206
rect 14721 12538 14777 12540
rect 14801 12538 14857 12540
rect 14881 12538 14937 12540
rect 14961 12538 15017 12540
rect 14721 12486 14767 12538
rect 14767 12486 14777 12538
rect 14801 12486 14831 12538
rect 14831 12486 14843 12538
rect 14843 12486 14857 12538
rect 14881 12486 14895 12538
rect 14895 12486 14907 12538
rect 14907 12486 14937 12538
rect 14961 12486 14971 12538
rect 14971 12486 15017 12538
rect 14721 12484 14777 12486
rect 14801 12484 14857 12486
rect 14881 12484 14937 12486
rect 14961 12484 15017 12486
rect 14721 11450 14777 11452
rect 14801 11450 14857 11452
rect 14881 11450 14937 11452
rect 14961 11450 15017 11452
rect 14721 11398 14767 11450
rect 14767 11398 14777 11450
rect 14801 11398 14831 11450
rect 14831 11398 14843 11450
rect 14843 11398 14857 11450
rect 14881 11398 14895 11450
rect 14895 11398 14907 11450
rect 14907 11398 14937 11450
rect 14961 11398 14971 11450
rect 14971 11398 15017 11450
rect 14721 11396 14777 11398
rect 14801 11396 14857 11398
rect 14881 11396 14937 11398
rect 14961 11396 15017 11398
rect 14721 10362 14777 10364
rect 14801 10362 14857 10364
rect 14881 10362 14937 10364
rect 14961 10362 15017 10364
rect 14721 10310 14767 10362
rect 14767 10310 14777 10362
rect 14801 10310 14831 10362
rect 14831 10310 14843 10362
rect 14843 10310 14857 10362
rect 14881 10310 14895 10362
rect 14895 10310 14907 10362
rect 14907 10310 14937 10362
rect 14961 10310 14971 10362
rect 14971 10310 15017 10362
rect 14721 10308 14777 10310
rect 14801 10308 14857 10310
rect 14881 10308 14937 10310
rect 14961 10308 15017 10310
rect 16687 14170 16743 14172
rect 16767 14170 16823 14172
rect 16847 14170 16903 14172
rect 16927 14170 16983 14172
rect 16687 14118 16733 14170
rect 16733 14118 16743 14170
rect 16767 14118 16797 14170
rect 16797 14118 16809 14170
rect 16809 14118 16823 14170
rect 16847 14118 16861 14170
rect 16861 14118 16873 14170
rect 16873 14118 16903 14170
rect 16927 14118 16937 14170
rect 16937 14118 16983 14170
rect 16687 14116 16743 14118
rect 16767 14116 16823 14118
rect 16847 14116 16903 14118
rect 16927 14116 16983 14118
rect 16687 13082 16743 13084
rect 16767 13082 16823 13084
rect 16847 13082 16903 13084
rect 16927 13082 16983 13084
rect 16687 13030 16733 13082
rect 16733 13030 16743 13082
rect 16767 13030 16797 13082
rect 16797 13030 16809 13082
rect 16809 13030 16823 13082
rect 16847 13030 16861 13082
rect 16861 13030 16873 13082
rect 16873 13030 16903 13082
rect 16927 13030 16937 13082
rect 16937 13030 16983 13082
rect 16687 13028 16743 13030
rect 16767 13028 16823 13030
rect 16847 13028 16903 13030
rect 16927 13028 16983 13030
rect 16687 11994 16743 11996
rect 16767 11994 16823 11996
rect 16847 11994 16903 11996
rect 16927 11994 16983 11996
rect 16687 11942 16733 11994
rect 16733 11942 16743 11994
rect 16767 11942 16797 11994
rect 16797 11942 16809 11994
rect 16809 11942 16823 11994
rect 16847 11942 16861 11994
rect 16861 11942 16873 11994
rect 16873 11942 16903 11994
rect 16927 11942 16937 11994
rect 16937 11942 16983 11994
rect 16687 11940 16743 11942
rect 16767 11940 16823 11942
rect 16847 11940 16903 11942
rect 16927 11940 16983 11942
rect 16687 10906 16743 10908
rect 16767 10906 16823 10908
rect 16847 10906 16903 10908
rect 16927 10906 16983 10908
rect 16687 10854 16733 10906
rect 16733 10854 16743 10906
rect 16767 10854 16797 10906
rect 16797 10854 16809 10906
rect 16809 10854 16823 10906
rect 16847 10854 16861 10906
rect 16861 10854 16873 10906
rect 16873 10854 16903 10906
rect 16927 10854 16937 10906
rect 16937 10854 16983 10906
rect 16687 10852 16743 10854
rect 16767 10852 16823 10854
rect 16847 10852 16903 10854
rect 16927 10852 16983 10854
rect 16687 9818 16743 9820
rect 16767 9818 16823 9820
rect 16847 9818 16903 9820
rect 16927 9818 16983 9820
rect 16687 9766 16733 9818
rect 16733 9766 16743 9818
rect 16767 9766 16797 9818
rect 16797 9766 16809 9818
rect 16809 9766 16823 9818
rect 16847 9766 16861 9818
rect 16861 9766 16873 9818
rect 16873 9766 16903 9818
rect 16927 9766 16937 9818
rect 16937 9766 16983 9818
rect 16687 9764 16743 9766
rect 16767 9764 16823 9766
rect 16847 9764 16903 9766
rect 16927 9764 16983 9766
rect 14721 9274 14777 9276
rect 14801 9274 14857 9276
rect 14881 9274 14937 9276
rect 14961 9274 15017 9276
rect 14721 9222 14767 9274
rect 14767 9222 14777 9274
rect 14801 9222 14831 9274
rect 14831 9222 14843 9274
rect 14843 9222 14857 9274
rect 14881 9222 14895 9274
rect 14895 9222 14907 9274
rect 14907 9222 14937 9274
rect 14961 9222 14971 9274
rect 14971 9222 15017 9274
rect 14721 9220 14777 9222
rect 14801 9220 14857 9222
rect 14881 9220 14937 9222
rect 14961 9220 15017 9222
rect 14721 8186 14777 8188
rect 14801 8186 14857 8188
rect 14881 8186 14937 8188
rect 14961 8186 15017 8188
rect 14721 8134 14767 8186
rect 14767 8134 14777 8186
rect 14801 8134 14831 8186
rect 14831 8134 14843 8186
rect 14843 8134 14857 8186
rect 14881 8134 14895 8186
rect 14895 8134 14907 8186
rect 14907 8134 14937 8186
rect 14961 8134 14971 8186
rect 14971 8134 15017 8186
rect 14721 8132 14777 8134
rect 14801 8132 14857 8134
rect 14881 8132 14937 8134
rect 14961 8132 15017 8134
rect 16687 8730 16743 8732
rect 16767 8730 16823 8732
rect 16847 8730 16903 8732
rect 16927 8730 16983 8732
rect 16687 8678 16733 8730
rect 16733 8678 16743 8730
rect 16767 8678 16797 8730
rect 16797 8678 16809 8730
rect 16809 8678 16823 8730
rect 16847 8678 16861 8730
rect 16861 8678 16873 8730
rect 16873 8678 16903 8730
rect 16927 8678 16937 8730
rect 16937 8678 16983 8730
rect 16687 8676 16743 8678
rect 16767 8676 16823 8678
rect 16847 8676 16903 8678
rect 16927 8676 16983 8678
rect 16687 7642 16743 7644
rect 16767 7642 16823 7644
rect 16847 7642 16903 7644
rect 16927 7642 16983 7644
rect 16687 7590 16733 7642
rect 16733 7590 16743 7642
rect 16767 7590 16797 7642
rect 16797 7590 16809 7642
rect 16809 7590 16823 7642
rect 16847 7590 16861 7642
rect 16861 7590 16873 7642
rect 16873 7590 16903 7642
rect 16927 7590 16937 7642
rect 16937 7590 16983 7642
rect 16687 7588 16743 7590
rect 16767 7588 16823 7590
rect 16847 7588 16903 7590
rect 16927 7588 16983 7590
rect 12754 6554 12810 6556
rect 12834 6554 12890 6556
rect 12914 6554 12970 6556
rect 12994 6554 13050 6556
rect 12754 6502 12800 6554
rect 12800 6502 12810 6554
rect 12834 6502 12864 6554
rect 12864 6502 12876 6554
rect 12876 6502 12890 6554
rect 12914 6502 12928 6554
rect 12928 6502 12940 6554
rect 12940 6502 12970 6554
rect 12994 6502 13004 6554
rect 13004 6502 13050 6554
rect 12754 6500 12810 6502
rect 12834 6500 12890 6502
rect 12914 6500 12970 6502
rect 12994 6500 13050 6502
rect 10788 6010 10844 6012
rect 10868 6010 10924 6012
rect 10948 6010 11004 6012
rect 11028 6010 11084 6012
rect 10788 5958 10834 6010
rect 10834 5958 10844 6010
rect 10868 5958 10898 6010
rect 10898 5958 10910 6010
rect 10910 5958 10924 6010
rect 10948 5958 10962 6010
rect 10962 5958 10974 6010
rect 10974 5958 11004 6010
rect 11028 5958 11038 6010
rect 11038 5958 11084 6010
rect 10788 5956 10844 5958
rect 10868 5956 10924 5958
rect 10948 5956 11004 5958
rect 11028 5956 11084 5958
rect 10788 4922 10844 4924
rect 10868 4922 10924 4924
rect 10948 4922 11004 4924
rect 11028 4922 11084 4924
rect 10788 4870 10834 4922
rect 10834 4870 10844 4922
rect 10868 4870 10898 4922
rect 10898 4870 10910 4922
rect 10910 4870 10924 4922
rect 10948 4870 10962 4922
rect 10962 4870 10974 4922
rect 10974 4870 11004 4922
rect 11028 4870 11038 4922
rect 11038 4870 11084 4922
rect 10788 4868 10844 4870
rect 10868 4868 10924 4870
rect 10948 4868 11004 4870
rect 11028 4868 11084 4870
rect 8821 3290 8877 3292
rect 8901 3290 8957 3292
rect 8981 3290 9037 3292
rect 9061 3290 9117 3292
rect 8821 3238 8867 3290
rect 8867 3238 8877 3290
rect 8901 3238 8931 3290
rect 8931 3238 8943 3290
rect 8943 3238 8957 3290
rect 8981 3238 8995 3290
rect 8995 3238 9007 3290
rect 9007 3238 9037 3290
rect 9061 3238 9071 3290
rect 9071 3238 9117 3290
rect 8821 3236 8877 3238
rect 8901 3236 8957 3238
rect 8981 3236 9037 3238
rect 9061 3236 9117 3238
rect 10788 3834 10844 3836
rect 10868 3834 10924 3836
rect 10948 3834 11004 3836
rect 11028 3834 11084 3836
rect 10788 3782 10834 3834
rect 10834 3782 10844 3834
rect 10868 3782 10898 3834
rect 10898 3782 10910 3834
rect 10910 3782 10924 3834
rect 10948 3782 10962 3834
rect 10962 3782 10974 3834
rect 10974 3782 11004 3834
rect 11028 3782 11038 3834
rect 11038 3782 11084 3834
rect 10788 3780 10844 3782
rect 10868 3780 10924 3782
rect 10948 3780 11004 3782
rect 11028 3780 11084 3782
rect 12754 5466 12810 5468
rect 12834 5466 12890 5468
rect 12914 5466 12970 5468
rect 12994 5466 13050 5468
rect 12754 5414 12800 5466
rect 12800 5414 12810 5466
rect 12834 5414 12864 5466
rect 12864 5414 12876 5466
rect 12876 5414 12890 5466
rect 12914 5414 12928 5466
rect 12928 5414 12940 5466
rect 12940 5414 12970 5466
rect 12994 5414 13004 5466
rect 13004 5414 13050 5466
rect 12754 5412 12810 5414
rect 12834 5412 12890 5414
rect 12914 5412 12970 5414
rect 12994 5412 13050 5414
rect 14721 7098 14777 7100
rect 14801 7098 14857 7100
rect 14881 7098 14937 7100
rect 14961 7098 15017 7100
rect 14721 7046 14767 7098
rect 14767 7046 14777 7098
rect 14801 7046 14831 7098
rect 14831 7046 14843 7098
rect 14843 7046 14857 7098
rect 14881 7046 14895 7098
rect 14895 7046 14907 7098
rect 14907 7046 14937 7098
rect 14961 7046 14971 7098
rect 14971 7046 15017 7098
rect 14721 7044 14777 7046
rect 14801 7044 14857 7046
rect 14881 7044 14937 7046
rect 14961 7044 15017 7046
rect 16687 6554 16743 6556
rect 16767 6554 16823 6556
rect 16847 6554 16903 6556
rect 16927 6554 16983 6556
rect 16687 6502 16733 6554
rect 16733 6502 16743 6554
rect 16767 6502 16797 6554
rect 16797 6502 16809 6554
rect 16809 6502 16823 6554
rect 16847 6502 16861 6554
rect 16861 6502 16873 6554
rect 16873 6502 16903 6554
rect 16927 6502 16937 6554
rect 16937 6502 16983 6554
rect 16687 6500 16743 6502
rect 16767 6500 16823 6502
rect 16847 6500 16903 6502
rect 16927 6500 16983 6502
rect 12754 4378 12810 4380
rect 12834 4378 12890 4380
rect 12914 4378 12970 4380
rect 12994 4378 13050 4380
rect 12754 4326 12800 4378
rect 12800 4326 12810 4378
rect 12834 4326 12864 4378
rect 12864 4326 12876 4378
rect 12876 4326 12890 4378
rect 12914 4326 12928 4378
rect 12928 4326 12940 4378
rect 12940 4326 12970 4378
rect 12994 4326 13004 4378
rect 13004 4326 13050 4378
rect 12754 4324 12810 4326
rect 12834 4324 12890 4326
rect 12914 4324 12970 4326
rect 12994 4324 13050 4326
rect 12754 3290 12810 3292
rect 12834 3290 12890 3292
rect 12914 3290 12970 3292
rect 12994 3290 13050 3292
rect 12754 3238 12800 3290
rect 12800 3238 12810 3290
rect 12834 3238 12864 3290
rect 12864 3238 12876 3290
rect 12876 3238 12890 3290
rect 12914 3238 12928 3290
rect 12928 3238 12940 3290
rect 12940 3238 12970 3290
rect 12994 3238 13004 3290
rect 13004 3238 13050 3290
rect 12754 3236 12810 3238
rect 12834 3236 12890 3238
rect 12914 3236 12970 3238
rect 12994 3236 13050 3238
rect 10788 2746 10844 2748
rect 10868 2746 10924 2748
rect 10948 2746 11004 2748
rect 11028 2746 11084 2748
rect 10788 2694 10834 2746
rect 10834 2694 10844 2746
rect 10868 2694 10898 2746
rect 10898 2694 10910 2746
rect 10910 2694 10924 2746
rect 10948 2694 10962 2746
rect 10962 2694 10974 2746
rect 10974 2694 11004 2746
rect 11028 2694 11038 2746
rect 11038 2694 11084 2746
rect 10788 2692 10844 2694
rect 10868 2692 10924 2694
rect 10948 2692 11004 2694
rect 11028 2692 11084 2694
rect 14721 6010 14777 6012
rect 14801 6010 14857 6012
rect 14881 6010 14937 6012
rect 14961 6010 15017 6012
rect 14721 5958 14767 6010
rect 14767 5958 14777 6010
rect 14801 5958 14831 6010
rect 14831 5958 14843 6010
rect 14843 5958 14857 6010
rect 14881 5958 14895 6010
rect 14895 5958 14907 6010
rect 14907 5958 14937 6010
rect 14961 5958 14971 6010
rect 14971 5958 15017 6010
rect 14721 5956 14777 5958
rect 14801 5956 14857 5958
rect 14881 5956 14937 5958
rect 14961 5956 15017 5958
rect 16687 5466 16743 5468
rect 16767 5466 16823 5468
rect 16847 5466 16903 5468
rect 16927 5466 16983 5468
rect 16687 5414 16733 5466
rect 16733 5414 16743 5466
rect 16767 5414 16797 5466
rect 16797 5414 16809 5466
rect 16809 5414 16823 5466
rect 16847 5414 16861 5466
rect 16861 5414 16873 5466
rect 16873 5414 16903 5466
rect 16927 5414 16937 5466
rect 16937 5414 16983 5466
rect 16687 5412 16743 5414
rect 16767 5412 16823 5414
rect 16847 5412 16903 5414
rect 16927 5412 16983 5414
rect 14721 4922 14777 4924
rect 14801 4922 14857 4924
rect 14881 4922 14937 4924
rect 14961 4922 15017 4924
rect 14721 4870 14767 4922
rect 14767 4870 14777 4922
rect 14801 4870 14831 4922
rect 14831 4870 14843 4922
rect 14843 4870 14857 4922
rect 14881 4870 14895 4922
rect 14895 4870 14907 4922
rect 14907 4870 14937 4922
rect 14961 4870 14971 4922
rect 14971 4870 15017 4922
rect 14721 4868 14777 4870
rect 14801 4868 14857 4870
rect 14881 4868 14937 4870
rect 14961 4868 15017 4870
rect 14721 3834 14777 3836
rect 14801 3834 14857 3836
rect 14881 3834 14937 3836
rect 14961 3834 15017 3836
rect 14721 3782 14767 3834
rect 14767 3782 14777 3834
rect 14801 3782 14831 3834
rect 14831 3782 14843 3834
rect 14843 3782 14857 3834
rect 14881 3782 14895 3834
rect 14895 3782 14907 3834
rect 14907 3782 14937 3834
rect 14961 3782 14971 3834
rect 14971 3782 15017 3834
rect 14721 3780 14777 3782
rect 14801 3780 14857 3782
rect 14881 3780 14937 3782
rect 14961 3780 15017 3782
rect 16687 4378 16743 4380
rect 16767 4378 16823 4380
rect 16847 4378 16903 4380
rect 16927 4378 16983 4380
rect 16687 4326 16733 4378
rect 16733 4326 16743 4378
rect 16767 4326 16797 4378
rect 16797 4326 16809 4378
rect 16809 4326 16823 4378
rect 16847 4326 16861 4378
rect 16861 4326 16873 4378
rect 16873 4326 16903 4378
rect 16927 4326 16937 4378
rect 16937 4326 16983 4378
rect 16687 4324 16743 4326
rect 16767 4324 16823 4326
rect 16847 4324 16903 4326
rect 16927 4324 16983 4326
rect 14721 2746 14777 2748
rect 14801 2746 14857 2748
rect 14881 2746 14937 2748
rect 14961 2746 15017 2748
rect 14721 2694 14767 2746
rect 14767 2694 14777 2746
rect 14801 2694 14831 2746
rect 14831 2694 14843 2746
rect 14843 2694 14857 2746
rect 14881 2694 14895 2746
rect 14895 2694 14907 2746
rect 14907 2694 14937 2746
rect 14961 2694 14971 2746
rect 14971 2694 15017 2746
rect 14721 2692 14777 2694
rect 14801 2692 14857 2694
rect 14881 2692 14937 2694
rect 14961 2692 15017 2694
rect 4888 2202 4944 2204
rect 4968 2202 5024 2204
rect 5048 2202 5104 2204
rect 5128 2202 5184 2204
rect 4888 2150 4934 2202
rect 4934 2150 4944 2202
rect 4968 2150 4998 2202
rect 4998 2150 5010 2202
rect 5010 2150 5024 2202
rect 5048 2150 5062 2202
rect 5062 2150 5074 2202
rect 5074 2150 5104 2202
rect 5128 2150 5138 2202
rect 5138 2150 5184 2202
rect 4888 2148 4944 2150
rect 4968 2148 5024 2150
rect 5048 2148 5104 2150
rect 5128 2148 5184 2150
rect 8821 2202 8877 2204
rect 8901 2202 8957 2204
rect 8981 2202 9037 2204
rect 9061 2202 9117 2204
rect 8821 2150 8867 2202
rect 8867 2150 8877 2202
rect 8901 2150 8931 2202
rect 8931 2150 8943 2202
rect 8943 2150 8957 2202
rect 8981 2150 8995 2202
rect 8995 2150 9007 2202
rect 9007 2150 9037 2202
rect 9061 2150 9071 2202
rect 9071 2150 9117 2202
rect 8821 2148 8877 2150
rect 8901 2148 8957 2150
rect 8981 2148 9037 2150
rect 9061 2148 9117 2150
rect 12754 2202 12810 2204
rect 12834 2202 12890 2204
rect 12914 2202 12970 2204
rect 12994 2202 13050 2204
rect 12754 2150 12800 2202
rect 12800 2150 12810 2202
rect 12834 2150 12864 2202
rect 12864 2150 12876 2202
rect 12876 2150 12890 2202
rect 12914 2150 12928 2202
rect 12928 2150 12940 2202
rect 12940 2150 12970 2202
rect 12994 2150 13004 2202
rect 13004 2150 13050 2202
rect 12754 2148 12810 2150
rect 12834 2148 12890 2150
rect 12914 2148 12970 2150
rect 12994 2148 13050 2150
rect 16687 3290 16743 3292
rect 16767 3290 16823 3292
rect 16847 3290 16903 3292
rect 16927 3290 16983 3292
rect 16687 3238 16733 3290
rect 16733 3238 16743 3290
rect 16767 3238 16797 3290
rect 16797 3238 16809 3290
rect 16809 3238 16823 3290
rect 16847 3238 16861 3290
rect 16861 3238 16873 3290
rect 16873 3238 16903 3290
rect 16927 3238 16937 3290
rect 16937 3238 16983 3290
rect 16687 3236 16743 3238
rect 16767 3236 16823 3238
rect 16847 3236 16903 3238
rect 16927 3236 16983 3238
rect 16687 2202 16743 2204
rect 16767 2202 16823 2204
rect 16847 2202 16903 2204
rect 16927 2202 16983 2204
rect 16687 2150 16733 2202
rect 16733 2150 16743 2202
rect 16767 2150 16797 2202
rect 16797 2150 16809 2202
rect 16809 2150 16823 2202
rect 16847 2150 16861 2202
rect 16861 2150 16873 2202
rect 16873 2150 16903 2202
rect 16927 2150 16937 2202
rect 16937 2150 16983 2202
rect 16687 2148 16743 2150
rect 16767 2148 16823 2150
rect 16847 2148 16903 2150
rect 16927 2148 16983 2150
<< metal3 >>
rect 2912 15808 3228 15809
rect 2912 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3228 15808
rect 2912 15743 3228 15744
rect 6845 15808 7161 15809
rect 6845 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7161 15808
rect 6845 15743 7161 15744
rect 10778 15808 11094 15809
rect 10778 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11094 15808
rect 10778 15743 11094 15744
rect 14711 15808 15027 15809
rect 14711 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15027 15808
rect 14711 15743 15027 15744
rect 4878 15264 5194 15265
rect 4878 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5194 15264
rect 4878 15199 5194 15200
rect 8811 15264 9127 15265
rect 8811 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9127 15264
rect 8811 15199 9127 15200
rect 12744 15264 13060 15265
rect 12744 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13060 15264
rect 12744 15199 13060 15200
rect 16677 15264 16993 15265
rect 16677 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16993 15264
rect 16677 15199 16993 15200
rect 2912 14720 3228 14721
rect 2912 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3228 14720
rect 2912 14655 3228 14656
rect 6845 14720 7161 14721
rect 6845 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7161 14720
rect 6845 14655 7161 14656
rect 10778 14720 11094 14721
rect 10778 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11094 14720
rect 10778 14655 11094 14656
rect 14711 14720 15027 14721
rect 14711 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15027 14720
rect 14711 14655 15027 14656
rect 4878 14176 5194 14177
rect 4878 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5194 14176
rect 4878 14111 5194 14112
rect 8811 14176 9127 14177
rect 8811 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9127 14176
rect 8811 14111 9127 14112
rect 12744 14176 13060 14177
rect 12744 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13060 14176
rect 12744 14111 13060 14112
rect 16677 14176 16993 14177
rect 16677 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16993 14176
rect 16677 14111 16993 14112
rect 2912 13632 3228 13633
rect 2912 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3228 13632
rect 2912 13567 3228 13568
rect 6845 13632 7161 13633
rect 6845 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7161 13632
rect 6845 13567 7161 13568
rect 10778 13632 11094 13633
rect 10778 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11094 13632
rect 10778 13567 11094 13568
rect 14711 13632 15027 13633
rect 14711 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15027 13632
rect 14711 13567 15027 13568
rect 4878 13088 5194 13089
rect 4878 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5194 13088
rect 4878 13023 5194 13024
rect 8811 13088 9127 13089
rect 8811 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9127 13088
rect 8811 13023 9127 13024
rect 12744 13088 13060 13089
rect 12744 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13060 13088
rect 12744 13023 13060 13024
rect 16677 13088 16993 13089
rect 16677 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16993 13088
rect 16677 13023 16993 13024
rect 2912 12544 3228 12545
rect 2912 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3228 12544
rect 2912 12479 3228 12480
rect 6845 12544 7161 12545
rect 6845 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7161 12544
rect 6845 12479 7161 12480
rect 10778 12544 11094 12545
rect 10778 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11094 12544
rect 10778 12479 11094 12480
rect 14711 12544 15027 12545
rect 14711 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15027 12544
rect 14711 12479 15027 12480
rect 4878 12000 5194 12001
rect 4878 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5194 12000
rect 4878 11935 5194 11936
rect 8811 12000 9127 12001
rect 8811 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9127 12000
rect 8811 11935 9127 11936
rect 12744 12000 13060 12001
rect 12744 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13060 12000
rect 12744 11935 13060 11936
rect 16677 12000 16993 12001
rect 16677 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16993 12000
rect 16677 11935 16993 11936
rect 2912 11456 3228 11457
rect 2912 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3228 11456
rect 2912 11391 3228 11392
rect 6845 11456 7161 11457
rect 6845 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7161 11456
rect 6845 11391 7161 11392
rect 10778 11456 11094 11457
rect 10778 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11094 11456
rect 10778 11391 11094 11392
rect 14711 11456 15027 11457
rect 14711 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15027 11456
rect 14711 11391 15027 11392
rect 4878 10912 5194 10913
rect 4878 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5194 10912
rect 4878 10847 5194 10848
rect 8811 10912 9127 10913
rect 8811 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9127 10912
rect 8811 10847 9127 10848
rect 12744 10912 13060 10913
rect 12744 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13060 10912
rect 12744 10847 13060 10848
rect 16677 10912 16993 10913
rect 16677 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16993 10912
rect 16677 10847 16993 10848
rect 2912 10368 3228 10369
rect 2912 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3228 10368
rect 2912 10303 3228 10304
rect 6845 10368 7161 10369
rect 6845 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7161 10368
rect 6845 10303 7161 10304
rect 10778 10368 11094 10369
rect 10778 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11094 10368
rect 10778 10303 11094 10304
rect 14711 10368 15027 10369
rect 14711 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15027 10368
rect 14711 10303 15027 10304
rect 4878 9824 5194 9825
rect 4878 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5194 9824
rect 4878 9759 5194 9760
rect 8811 9824 9127 9825
rect 8811 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9127 9824
rect 8811 9759 9127 9760
rect 12744 9824 13060 9825
rect 12744 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13060 9824
rect 12744 9759 13060 9760
rect 16677 9824 16993 9825
rect 16677 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16993 9824
rect 16677 9759 16993 9760
rect 2912 9280 3228 9281
rect 2912 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3228 9280
rect 2912 9215 3228 9216
rect 6845 9280 7161 9281
rect 6845 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7161 9280
rect 6845 9215 7161 9216
rect 10778 9280 11094 9281
rect 10778 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11094 9280
rect 10778 9215 11094 9216
rect 14711 9280 15027 9281
rect 14711 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15027 9280
rect 14711 9215 15027 9216
rect 4878 8736 5194 8737
rect 4878 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5194 8736
rect 4878 8671 5194 8672
rect 8811 8736 9127 8737
rect 8811 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9127 8736
rect 8811 8671 9127 8672
rect 12744 8736 13060 8737
rect 12744 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13060 8736
rect 12744 8671 13060 8672
rect 16677 8736 16993 8737
rect 16677 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16993 8736
rect 16677 8671 16993 8672
rect 2912 8192 3228 8193
rect 2912 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3228 8192
rect 2912 8127 3228 8128
rect 6845 8192 7161 8193
rect 6845 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7161 8192
rect 6845 8127 7161 8128
rect 10778 8192 11094 8193
rect 10778 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11094 8192
rect 10778 8127 11094 8128
rect 14711 8192 15027 8193
rect 14711 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15027 8192
rect 14711 8127 15027 8128
rect 4878 7648 5194 7649
rect 4878 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5194 7648
rect 4878 7583 5194 7584
rect 8811 7648 9127 7649
rect 8811 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9127 7648
rect 8811 7583 9127 7584
rect 12744 7648 13060 7649
rect 12744 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13060 7648
rect 12744 7583 13060 7584
rect 16677 7648 16993 7649
rect 16677 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16993 7648
rect 16677 7583 16993 7584
rect 2912 7104 3228 7105
rect 2912 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3228 7104
rect 2912 7039 3228 7040
rect 6845 7104 7161 7105
rect 6845 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7161 7104
rect 6845 7039 7161 7040
rect 10778 7104 11094 7105
rect 10778 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11094 7104
rect 10778 7039 11094 7040
rect 14711 7104 15027 7105
rect 14711 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15027 7104
rect 14711 7039 15027 7040
rect 4878 6560 5194 6561
rect 4878 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5194 6560
rect 4878 6495 5194 6496
rect 8811 6560 9127 6561
rect 8811 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9127 6560
rect 8811 6495 9127 6496
rect 12744 6560 13060 6561
rect 12744 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13060 6560
rect 12744 6495 13060 6496
rect 16677 6560 16993 6561
rect 16677 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16993 6560
rect 16677 6495 16993 6496
rect 2912 6016 3228 6017
rect 2912 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3228 6016
rect 2912 5951 3228 5952
rect 6845 6016 7161 6017
rect 6845 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7161 6016
rect 6845 5951 7161 5952
rect 10778 6016 11094 6017
rect 10778 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11094 6016
rect 10778 5951 11094 5952
rect 14711 6016 15027 6017
rect 14711 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15027 6016
rect 14711 5951 15027 5952
rect 4878 5472 5194 5473
rect 4878 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5194 5472
rect 4878 5407 5194 5408
rect 8811 5472 9127 5473
rect 8811 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9127 5472
rect 8811 5407 9127 5408
rect 12744 5472 13060 5473
rect 12744 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13060 5472
rect 12744 5407 13060 5408
rect 16677 5472 16993 5473
rect 16677 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16993 5472
rect 16677 5407 16993 5408
rect 2912 4928 3228 4929
rect 2912 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3228 4928
rect 2912 4863 3228 4864
rect 6845 4928 7161 4929
rect 6845 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7161 4928
rect 6845 4863 7161 4864
rect 10778 4928 11094 4929
rect 10778 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11094 4928
rect 10778 4863 11094 4864
rect 14711 4928 15027 4929
rect 14711 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15027 4928
rect 14711 4863 15027 4864
rect 4878 4384 5194 4385
rect 4878 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5194 4384
rect 4878 4319 5194 4320
rect 8811 4384 9127 4385
rect 8811 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9127 4384
rect 8811 4319 9127 4320
rect 12744 4384 13060 4385
rect 12744 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13060 4384
rect 12744 4319 13060 4320
rect 16677 4384 16993 4385
rect 16677 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16993 4384
rect 16677 4319 16993 4320
rect 2912 3840 3228 3841
rect 2912 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3228 3840
rect 2912 3775 3228 3776
rect 6845 3840 7161 3841
rect 6845 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7161 3840
rect 6845 3775 7161 3776
rect 10778 3840 11094 3841
rect 10778 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11094 3840
rect 10778 3775 11094 3776
rect 14711 3840 15027 3841
rect 14711 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15027 3840
rect 14711 3775 15027 3776
rect 4878 3296 5194 3297
rect 4878 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5194 3296
rect 4878 3231 5194 3232
rect 8811 3296 9127 3297
rect 8811 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9127 3296
rect 8811 3231 9127 3232
rect 12744 3296 13060 3297
rect 12744 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13060 3296
rect 12744 3231 13060 3232
rect 16677 3296 16993 3297
rect 16677 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16993 3296
rect 16677 3231 16993 3232
rect 2912 2752 3228 2753
rect 2912 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3228 2752
rect 2912 2687 3228 2688
rect 6845 2752 7161 2753
rect 6845 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7161 2752
rect 6845 2687 7161 2688
rect 10778 2752 11094 2753
rect 10778 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11094 2752
rect 10778 2687 11094 2688
rect 14711 2752 15027 2753
rect 14711 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15027 2752
rect 14711 2687 15027 2688
rect 4878 2208 5194 2209
rect 4878 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5194 2208
rect 4878 2143 5194 2144
rect 8811 2208 9127 2209
rect 8811 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9127 2208
rect 8811 2143 9127 2144
rect 12744 2208 13060 2209
rect 12744 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13060 2208
rect 12744 2143 13060 2144
rect 16677 2208 16993 2209
rect 16677 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16993 2208
rect 16677 2143 16993 2144
<< via3 >>
rect 2918 15804 2982 15808
rect 2918 15748 2922 15804
rect 2922 15748 2978 15804
rect 2978 15748 2982 15804
rect 2918 15744 2982 15748
rect 2998 15804 3062 15808
rect 2998 15748 3002 15804
rect 3002 15748 3058 15804
rect 3058 15748 3062 15804
rect 2998 15744 3062 15748
rect 3078 15804 3142 15808
rect 3078 15748 3082 15804
rect 3082 15748 3138 15804
rect 3138 15748 3142 15804
rect 3078 15744 3142 15748
rect 3158 15804 3222 15808
rect 3158 15748 3162 15804
rect 3162 15748 3218 15804
rect 3218 15748 3222 15804
rect 3158 15744 3222 15748
rect 6851 15804 6915 15808
rect 6851 15748 6855 15804
rect 6855 15748 6911 15804
rect 6911 15748 6915 15804
rect 6851 15744 6915 15748
rect 6931 15804 6995 15808
rect 6931 15748 6935 15804
rect 6935 15748 6991 15804
rect 6991 15748 6995 15804
rect 6931 15744 6995 15748
rect 7011 15804 7075 15808
rect 7011 15748 7015 15804
rect 7015 15748 7071 15804
rect 7071 15748 7075 15804
rect 7011 15744 7075 15748
rect 7091 15804 7155 15808
rect 7091 15748 7095 15804
rect 7095 15748 7151 15804
rect 7151 15748 7155 15804
rect 7091 15744 7155 15748
rect 10784 15804 10848 15808
rect 10784 15748 10788 15804
rect 10788 15748 10844 15804
rect 10844 15748 10848 15804
rect 10784 15744 10848 15748
rect 10864 15804 10928 15808
rect 10864 15748 10868 15804
rect 10868 15748 10924 15804
rect 10924 15748 10928 15804
rect 10864 15744 10928 15748
rect 10944 15804 11008 15808
rect 10944 15748 10948 15804
rect 10948 15748 11004 15804
rect 11004 15748 11008 15804
rect 10944 15744 11008 15748
rect 11024 15804 11088 15808
rect 11024 15748 11028 15804
rect 11028 15748 11084 15804
rect 11084 15748 11088 15804
rect 11024 15744 11088 15748
rect 14717 15804 14781 15808
rect 14717 15748 14721 15804
rect 14721 15748 14777 15804
rect 14777 15748 14781 15804
rect 14717 15744 14781 15748
rect 14797 15804 14861 15808
rect 14797 15748 14801 15804
rect 14801 15748 14857 15804
rect 14857 15748 14861 15804
rect 14797 15744 14861 15748
rect 14877 15804 14941 15808
rect 14877 15748 14881 15804
rect 14881 15748 14937 15804
rect 14937 15748 14941 15804
rect 14877 15744 14941 15748
rect 14957 15804 15021 15808
rect 14957 15748 14961 15804
rect 14961 15748 15017 15804
rect 15017 15748 15021 15804
rect 14957 15744 15021 15748
rect 4884 15260 4948 15264
rect 4884 15204 4888 15260
rect 4888 15204 4944 15260
rect 4944 15204 4948 15260
rect 4884 15200 4948 15204
rect 4964 15260 5028 15264
rect 4964 15204 4968 15260
rect 4968 15204 5024 15260
rect 5024 15204 5028 15260
rect 4964 15200 5028 15204
rect 5044 15260 5108 15264
rect 5044 15204 5048 15260
rect 5048 15204 5104 15260
rect 5104 15204 5108 15260
rect 5044 15200 5108 15204
rect 5124 15260 5188 15264
rect 5124 15204 5128 15260
rect 5128 15204 5184 15260
rect 5184 15204 5188 15260
rect 5124 15200 5188 15204
rect 8817 15260 8881 15264
rect 8817 15204 8821 15260
rect 8821 15204 8877 15260
rect 8877 15204 8881 15260
rect 8817 15200 8881 15204
rect 8897 15260 8961 15264
rect 8897 15204 8901 15260
rect 8901 15204 8957 15260
rect 8957 15204 8961 15260
rect 8897 15200 8961 15204
rect 8977 15260 9041 15264
rect 8977 15204 8981 15260
rect 8981 15204 9037 15260
rect 9037 15204 9041 15260
rect 8977 15200 9041 15204
rect 9057 15260 9121 15264
rect 9057 15204 9061 15260
rect 9061 15204 9117 15260
rect 9117 15204 9121 15260
rect 9057 15200 9121 15204
rect 12750 15260 12814 15264
rect 12750 15204 12754 15260
rect 12754 15204 12810 15260
rect 12810 15204 12814 15260
rect 12750 15200 12814 15204
rect 12830 15260 12894 15264
rect 12830 15204 12834 15260
rect 12834 15204 12890 15260
rect 12890 15204 12894 15260
rect 12830 15200 12894 15204
rect 12910 15260 12974 15264
rect 12910 15204 12914 15260
rect 12914 15204 12970 15260
rect 12970 15204 12974 15260
rect 12910 15200 12974 15204
rect 12990 15260 13054 15264
rect 12990 15204 12994 15260
rect 12994 15204 13050 15260
rect 13050 15204 13054 15260
rect 12990 15200 13054 15204
rect 16683 15260 16747 15264
rect 16683 15204 16687 15260
rect 16687 15204 16743 15260
rect 16743 15204 16747 15260
rect 16683 15200 16747 15204
rect 16763 15260 16827 15264
rect 16763 15204 16767 15260
rect 16767 15204 16823 15260
rect 16823 15204 16827 15260
rect 16763 15200 16827 15204
rect 16843 15260 16907 15264
rect 16843 15204 16847 15260
rect 16847 15204 16903 15260
rect 16903 15204 16907 15260
rect 16843 15200 16907 15204
rect 16923 15260 16987 15264
rect 16923 15204 16927 15260
rect 16927 15204 16983 15260
rect 16983 15204 16987 15260
rect 16923 15200 16987 15204
rect 2918 14716 2982 14720
rect 2918 14660 2922 14716
rect 2922 14660 2978 14716
rect 2978 14660 2982 14716
rect 2918 14656 2982 14660
rect 2998 14716 3062 14720
rect 2998 14660 3002 14716
rect 3002 14660 3058 14716
rect 3058 14660 3062 14716
rect 2998 14656 3062 14660
rect 3078 14716 3142 14720
rect 3078 14660 3082 14716
rect 3082 14660 3138 14716
rect 3138 14660 3142 14716
rect 3078 14656 3142 14660
rect 3158 14716 3222 14720
rect 3158 14660 3162 14716
rect 3162 14660 3218 14716
rect 3218 14660 3222 14716
rect 3158 14656 3222 14660
rect 6851 14716 6915 14720
rect 6851 14660 6855 14716
rect 6855 14660 6911 14716
rect 6911 14660 6915 14716
rect 6851 14656 6915 14660
rect 6931 14716 6995 14720
rect 6931 14660 6935 14716
rect 6935 14660 6991 14716
rect 6991 14660 6995 14716
rect 6931 14656 6995 14660
rect 7011 14716 7075 14720
rect 7011 14660 7015 14716
rect 7015 14660 7071 14716
rect 7071 14660 7075 14716
rect 7011 14656 7075 14660
rect 7091 14716 7155 14720
rect 7091 14660 7095 14716
rect 7095 14660 7151 14716
rect 7151 14660 7155 14716
rect 7091 14656 7155 14660
rect 10784 14716 10848 14720
rect 10784 14660 10788 14716
rect 10788 14660 10844 14716
rect 10844 14660 10848 14716
rect 10784 14656 10848 14660
rect 10864 14716 10928 14720
rect 10864 14660 10868 14716
rect 10868 14660 10924 14716
rect 10924 14660 10928 14716
rect 10864 14656 10928 14660
rect 10944 14716 11008 14720
rect 10944 14660 10948 14716
rect 10948 14660 11004 14716
rect 11004 14660 11008 14716
rect 10944 14656 11008 14660
rect 11024 14716 11088 14720
rect 11024 14660 11028 14716
rect 11028 14660 11084 14716
rect 11084 14660 11088 14716
rect 11024 14656 11088 14660
rect 14717 14716 14781 14720
rect 14717 14660 14721 14716
rect 14721 14660 14777 14716
rect 14777 14660 14781 14716
rect 14717 14656 14781 14660
rect 14797 14716 14861 14720
rect 14797 14660 14801 14716
rect 14801 14660 14857 14716
rect 14857 14660 14861 14716
rect 14797 14656 14861 14660
rect 14877 14716 14941 14720
rect 14877 14660 14881 14716
rect 14881 14660 14937 14716
rect 14937 14660 14941 14716
rect 14877 14656 14941 14660
rect 14957 14716 15021 14720
rect 14957 14660 14961 14716
rect 14961 14660 15017 14716
rect 15017 14660 15021 14716
rect 14957 14656 15021 14660
rect 4884 14172 4948 14176
rect 4884 14116 4888 14172
rect 4888 14116 4944 14172
rect 4944 14116 4948 14172
rect 4884 14112 4948 14116
rect 4964 14172 5028 14176
rect 4964 14116 4968 14172
rect 4968 14116 5024 14172
rect 5024 14116 5028 14172
rect 4964 14112 5028 14116
rect 5044 14172 5108 14176
rect 5044 14116 5048 14172
rect 5048 14116 5104 14172
rect 5104 14116 5108 14172
rect 5044 14112 5108 14116
rect 5124 14172 5188 14176
rect 5124 14116 5128 14172
rect 5128 14116 5184 14172
rect 5184 14116 5188 14172
rect 5124 14112 5188 14116
rect 8817 14172 8881 14176
rect 8817 14116 8821 14172
rect 8821 14116 8877 14172
rect 8877 14116 8881 14172
rect 8817 14112 8881 14116
rect 8897 14172 8961 14176
rect 8897 14116 8901 14172
rect 8901 14116 8957 14172
rect 8957 14116 8961 14172
rect 8897 14112 8961 14116
rect 8977 14172 9041 14176
rect 8977 14116 8981 14172
rect 8981 14116 9037 14172
rect 9037 14116 9041 14172
rect 8977 14112 9041 14116
rect 9057 14172 9121 14176
rect 9057 14116 9061 14172
rect 9061 14116 9117 14172
rect 9117 14116 9121 14172
rect 9057 14112 9121 14116
rect 12750 14172 12814 14176
rect 12750 14116 12754 14172
rect 12754 14116 12810 14172
rect 12810 14116 12814 14172
rect 12750 14112 12814 14116
rect 12830 14172 12894 14176
rect 12830 14116 12834 14172
rect 12834 14116 12890 14172
rect 12890 14116 12894 14172
rect 12830 14112 12894 14116
rect 12910 14172 12974 14176
rect 12910 14116 12914 14172
rect 12914 14116 12970 14172
rect 12970 14116 12974 14172
rect 12910 14112 12974 14116
rect 12990 14172 13054 14176
rect 12990 14116 12994 14172
rect 12994 14116 13050 14172
rect 13050 14116 13054 14172
rect 12990 14112 13054 14116
rect 16683 14172 16747 14176
rect 16683 14116 16687 14172
rect 16687 14116 16743 14172
rect 16743 14116 16747 14172
rect 16683 14112 16747 14116
rect 16763 14172 16827 14176
rect 16763 14116 16767 14172
rect 16767 14116 16823 14172
rect 16823 14116 16827 14172
rect 16763 14112 16827 14116
rect 16843 14172 16907 14176
rect 16843 14116 16847 14172
rect 16847 14116 16903 14172
rect 16903 14116 16907 14172
rect 16843 14112 16907 14116
rect 16923 14172 16987 14176
rect 16923 14116 16927 14172
rect 16927 14116 16983 14172
rect 16983 14116 16987 14172
rect 16923 14112 16987 14116
rect 2918 13628 2982 13632
rect 2918 13572 2922 13628
rect 2922 13572 2978 13628
rect 2978 13572 2982 13628
rect 2918 13568 2982 13572
rect 2998 13628 3062 13632
rect 2998 13572 3002 13628
rect 3002 13572 3058 13628
rect 3058 13572 3062 13628
rect 2998 13568 3062 13572
rect 3078 13628 3142 13632
rect 3078 13572 3082 13628
rect 3082 13572 3138 13628
rect 3138 13572 3142 13628
rect 3078 13568 3142 13572
rect 3158 13628 3222 13632
rect 3158 13572 3162 13628
rect 3162 13572 3218 13628
rect 3218 13572 3222 13628
rect 3158 13568 3222 13572
rect 6851 13628 6915 13632
rect 6851 13572 6855 13628
rect 6855 13572 6911 13628
rect 6911 13572 6915 13628
rect 6851 13568 6915 13572
rect 6931 13628 6995 13632
rect 6931 13572 6935 13628
rect 6935 13572 6991 13628
rect 6991 13572 6995 13628
rect 6931 13568 6995 13572
rect 7011 13628 7075 13632
rect 7011 13572 7015 13628
rect 7015 13572 7071 13628
rect 7071 13572 7075 13628
rect 7011 13568 7075 13572
rect 7091 13628 7155 13632
rect 7091 13572 7095 13628
rect 7095 13572 7151 13628
rect 7151 13572 7155 13628
rect 7091 13568 7155 13572
rect 10784 13628 10848 13632
rect 10784 13572 10788 13628
rect 10788 13572 10844 13628
rect 10844 13572 10848 13628
rect 10784 13568 10848 13572
rect 10864 13628 10928 13632
rect 10864 13572 10868 13628
rect 10868 13572 10924 13628
rect 10924 13572 10928 13628
rect 10864 13568 10928 13572
rect 10944 13628 11008 13632
rect 10944 13572 10948 13628
rect 10948 13572 11004 13628
rect 11004 13572 11008 13628
rect 10944 13568 11008 13572
rect 11024 13628 11088 13632
rect 11024 13572 11028 13628
rect 11028 13572 11084 13628
rect 11084 13572 11088 13628
rect 11024 13568 11088 13572
rect 14717 13628 14781 13632
rect 14717 13572 14721 13628
rect 14721 13572 14777 13628
rect 14777 13572 14781 13628
rect 14717 13568 14781 13572
rect 14797 13628 14861 13632
rect 14797 13572 14801 13628
rect 14801 13572 14857 13628
rect 14857 13572 14861 13628
rect 14797 13568 14861 13572
rect 14877 13628 14941 13632
rect 14877 13572 14881 13628
rect 14881 13572 14937 13628
rect 14937 13572 14941 13628
rect 14877 13568 14941 13572
rect 14957 13628 15021 13632
rect 14957 13572 14961 13628
rect 14961 13572 15017 13628
rect 15017 13572 15021 13628
rect 14957 13568 15021 13572
rect 4884 13084 4948 13088
rect 4884 13028 4888 13084
rect 4888 13028 4944 13084
rect 4944 13028 4948 13084
rect 4884 13024 4948 13028
rect 4964 13084 5028 13088
rect 4964 13028 4968 13084
rect 4968 13028 5024 13084
rect 5024 13028 5028 13084
rect 4964 13024 5028 13028
rect 5044 13084 5108 13088
rect 5044 13028 5048 13084
rect 5048 13028 5104 13084
rect 5104 13028 5108 13084
rect 5044 13024 5108 13028
rect 5124 13084 5188 13088
rect 5124 13028 5128 13084
rect 5128 13028 5184 13084
rect 5184 13028 5188 13084
rect 5124 13024 5188 13028
rect 8817 13084 8881 13088
rect 8817 13028 8821 13084
rect 8821 13028 8877 13084
rect 8877 13028 8881 13084
rect 8817 13024 8881 13028
rect 8897 13084 8961 13088
rect 8897 13028 8901 13084
rect 8901 13028 8957 13084
rect 8957 13028 8961 13084
rect 8897 13024 8961 13028
rect 8977 13084 9041 13088
rect 8977 13028 8981 13084
rect 8981 13028 9037 13084
rect 9037 13028 9041 13084
rect 8977 13024 9041 13028
rect 9057 13084 9121 13088
rect 9057 13028 9061 13084
rect 9061 13028 9117 13084
rect 9117 13028 9121 13084
rect 9057 13024 9121 13028
rect 12750 13084 12814 13088
rect 12750 13028 12754 13084
rect 12754 13028 12810 13084
rect 12810 13028 12814 13084
rect 12750 13024 12814 13028
rect 12830 13084 12894 13088
rect 12830 13028 12834 13084
rect 12834 13028 12890 13084
rect 12890 13028 12894 13084
rect 12830 13024 12894 13028
rect 12910 13084 12974 13088
rect 12910 13028 12914 13084
rect 12914 13028 12970 13084
rect 12970 13028 12974 13084
rect 12910 13024 12974 13028
rect 12990 13084 13054 13088
rect 12990 13028 12994 13084
rect 12994 13028 13050 13084
rect 13050 13028 13054 13084
rect 12990 13024 13054 13028
rect 16683 13084 16747 13088
rect 16683 13028 16687 13084
rect 16687 13028 16743 13084
rect 16743 13028 16747 13084
rect 16683 13024 16747 13028
rect 16763 13084 16827 13088
rect 16763 13028 16767 13084
rect 16767 13028 16823 13084
rect 16823 13028 16827 13084
rect 16763 13024 16827 13028
rect 16843 13084 16907 13088
rect 16843 13028 16847 13084
rect 16847 13028 16903 13084
rect 16903 13028 16907 13084
rect 16843 13024 16907 13028
rect 16923 13084 16987 13088
rect 16923 13028 16927 13084
rect 16927 13028 16983 13084
rect 16983 13028 16987 13084
rect 16923 13024 16987 13028
rect 2918 12540 2982 12544
rect 2918 12484 2922 12540
rect 2922 12484 2978 12540
rect 2978 12484 2982 12540
rect 2918 12480 2982 12484
rect 2998 12540 3062 12544
rect 2998 12484 3002 12540
rect 3002 12484 3058 12540
rect 3058 12484 3062 12540
rect 2998 12480 3062 12484
rect 3078 12540 3142 12544
rect 3078 12484 3082 12540
rect 3082 12484 3138 12540
rect 3138 12484 3142 12540
rect 3078 12480 3142 12484
rect 3158 12540 3222 12544
rect 3158 12484 3162 12540
rect 3162 12484 3218 12540
rect 3218 12484 3222 12540
rect 3158 12480 3222 12484
rect 6851 12540 6915 12544
rect 6851 12484 6855 12540
rect 6855 12484 6911 12540
rect 6911 12484 6915 12540
rect 6851 12480 6915 12484
rect 6931 12540 6995 12544
rect 6931 12484 6935 12540
rect 6935 12484 6991 12540
rect 6991 12484 6995 12540
rect 6931 12480 6995 12484
rect 7011 12540 7075 12544
rect 7011 12484 7015 12540
rect 7015 12484 7071 12540
rect 7071 12484 7075 12540
rect 7011 12480 7075 12484
rect 7091 12540 7155 12544
rect 7091 12484 7095 12540
rect 7095 12484 7151 12540
rect 7151 12484 7155 12540
rect 7091 12480 7155 12484
rect 10784 12540 10848 12544
rect 10784 12484 10788 12540
rect 10788 12484 10844 12540
rect 10844 12484 10848 12540
rect 10784 12480 10848 12484
rect 10864 12540 10928 12544
rect 10864 12484 10868 12540
rect 10868 12484 10924 12540
rect 10924 12484 10928 12540
rect 10864 12480 10928 12484
rect 10944 12540 11008 12544
rect 10944 12484 10948 12540
rect 10948 12484 11004 12540
rect 11004 12484 11008 12540
rect 10944 12480 11008 12484
rect 11024 12540 11088 12544
rect 11024 12484 11028 12540
rect 11028 12484 11084 12540
rect 11084 12484 11088 12540
rect 11024 12480 11088 12484
rect 14717 12540 14781 12544
rect 14717 12484 14721 12540
rect 14721 12484 14777 12540
rect 14777 12484 14781 12540
rect 14717 12480 14781 12484
rect 14797 12540 14861 12544
rect 14797 12484 14801 12540
rect 14801 12484 14857 12540
rect 14857 12484 14861 12540
rect 14797 12480 14861 12484
rect 14877 12540 14941 12544
rect 14877 12484 14881 12540
rect 14881 12484 14937 12540
rect 14937 12484 14941 12540
rect 14877 12480 14941 12484
rect 14957 12540 15021 12544
rect 14957 12484 14961 12540
rect 14961 12484 15017 12540
rect 15017 12484 15021 12540
rect 14957 12480 15021 12484
rect 4884 11996 4948 12000
rect 4884 11940 4888 11996
rect 4888 11940 4944 11996
rect 4944 11940 4948 11996
rect 4884 11936 4948 11940
rect 4964 11996 5028 12000
rect 4964 11940 4968 11996
rect 4968 11940 5024 11996
rect 5024 11940 5028 11996
rect 4964 11936 5028 11940
rect 5044 11996 5108 12000
rect 5044 11940 5048 11996
rect 5048 11940 5104 11996
rect 5104 11940 5108 11996
rect 5044 11936 5108 11940
rect 5124 11996 5188 12000
rect 5124 11940 5128 11996
rect 5128 11940 5184 11996
rect 5184 11940 5188 11996
rect 5124 11936 5188 11940
rect 8817 11996 8881 12000
rect 8817 11940 8821 11996
rect 8821 11940 8877 11996
rect 8877 11940 8881 11996
rect 8817 11936 8881 11940
rect 8897 11996 8961 12000
rect 8897 11940 8901 11996
rect 8901 11940 8957 11996
rect 8957 11940 8961 11996
rect 8897 11936 8961 11940
rect 8977 11996 9041 12000
rect 8977 11940 8981 11996
rect 8981 11940 9037 11996
rect 9037 11940 9041 11996
rect 8977 11936 9041 11940
rect 9057 11996 9121 12000
rect 9057 11940 9061 11996
rect 9061 11940 9117 11996
rect 9117 11940 9121 11996
rect 9057 11936 9121 11940
rect 12750 11996 12814 12000
rect 12750 11940 12754 11996
rect 12754 11940 12810 11996
rect 12810 11940 12814 11996
rect 12750 11936 12814 11940
rect 12830 11996 12894 12000
rect 12830 11940 12834 11996
rect 12834 11940 12890 11996
rect 12890 11940 12894 11996
rect 12830 11936 12894 11940
rect 12910 11996 12974 12000
rect 12910 11940 12914 11996
rect 12914 11940 12970 11996
rect 12970 11940 12974 11996
rect 12910 11936 12974 11940
rect 12990 11996 13054 12000
rect 12990 11940 12994 11996
rect 12994 11940 13050 11996
rect 13050 11940 13054 11996
rect 12990 11936 13054 11940
rect 16683 11996 16747 12000
rect 16683 11940 16687 11996
rect 16687 11940 16743 11996
rect 16743 11940 16747 11996
rect 16683 11936 16747 11940
rect 16763 11996 16827 12000
rect 16763 11940 16767 11996
rect 16767 11940 16823 11996
rect 16823 11940 16827 11996
rect 16763 11936 16827 11940
rect 16843 11996 16907 12000
rect 16843 11940 16847 11996
rect 16847 11940 16903 11996
rect 16903 11940 16907 11996
rect 16843 11936 16907 11940
rect 16923 11996 16987 12000
rect 16923 11940 16927 11996
rect 16927 11940 16983 11996
rect 16983 11940 16987 11996
rect 16923 11936 16987 11940
rect 2918 11452 2982 11456
rect 2918 11396 2922 11452
rect 2922 11396 2978 11452
rect 2978 11396 2982 11452
rect 2918 11392 2982 11396
rect 2998 11452 3062 11456
rect 2998 11396 3002 11452
rect 3002 11396 3058 11452
rect 3058 11396 3062 11452
rect 2998 11392 3062 11396
rect 3078 11452 3142 11456
rect 3078 11396 3082 11452
rect 3082 11396 3138 11452
rect 3138 11396 3142 11452
rect 3078 11392 3142 11396
rect 3158 11452 3222 11456
rect 3158 11396 3162 11452
rect 3162 11396 3218 11452
rect 3218 11396 3222 11452
rect 3158 11392 3222 11396
rect 6851 11452 6915 11456
rect 6851 11396 6855 11452
rect 6855 11396 6911 11452
rect 6911 11396 6915 11452
rect 6851 11392 6915 11396
rect 6931 11452 6995 11456
rect 6931 11396 6935 11452
rect 6935 11396 6991 11452
rect 6991 11396 6995 11452
rect 6931 11392 6995 11396
rect 7011 11452 7075 11456
rect 7011 11396 7015 11452
rect 7015 11396 7071 11452
rect 7071 11396 7075 11452
rect 7011 11392 7075 11396
rect 7091 11452 7155 11456
rect 7091 11396 7095 11452
rect 7095 11396 7151 11452
rect 7151 11396 7155 11452
rect 7091 11392 7155 11396
rect 10784 11452 10848 11456
rect 10784 11396 10788 11452
rect 10788 11396 10844 11452
rect 10844 11396 10848 11452
rect 10784 11392 10848 11396
rect 10864 11452 10928 11456
rect 10864 11396 10868 11452
rect 10868 11396 10924 11452
rect 10924 11396 10928 11452
rect 10864 11392 10928 11396
rect 10944 11452 11008 11456
rect 10944 11396 10948 11452
rect 10948 11396 11004 11452
rect 11004 11396 11008 11452
rect 10944 11392 11008 11396
rect 11024 11452 11088 11456
rect 11024 11396 11028 11452
rect 11028 11396 11084 11452
rect 11084 11396 11088 11452
rect 11024 11392 11088 11396
rect 14717 11452 14781 11456
rect 14717 11396 14721 11452
rect 14721 11396 14777 11452
rect 14777 11396 14781 11452
rect 14717 11392 14781 11396
rect 14797 11452 14861 11456
rect 14797 11396 14801 11452
rect 14801 11396 14857 11452
rect 14857 11396 14861 11452
rect 14797 11392 14861 11396
rect 14877 11452 14941 11456
rect 14877 11396 14881 11452
rect 14881 11396 14937 11452
rect 14937 11396 14941 11452
rect 14877 11392 14941 11396
rect 14957 11452 15021 11456
rect 14957 11396 14961 11452
rect 14961 11396 15017 11452
rect 15017 11396 15021 11452
rect 14957 11392 15021 11396
rect 4884 10908 4948 10912
rect 4884 10852 4888 10908
rect 4888 10852 4944 10908
rect 4944 10852 4948 10908
rect 4884 10848 4948 10852
rect 4964 10908 5028 10912
rect 4964 10852 4968 10908
rect 4968 10852 5024 10908
rect 5024 10852 5028 10908
rect 4964 10848 5028 10852
rect 5044 10908 5108 10912
rect 5044 10852 5048 10908
rect 5048 10852 5104 10908
rect 5104 10852 5108 10908
rect 5044 10848 5108 10852
rect 5124 10908 5188 10912
rect 5124 10852 5128 10908
rect 5128 10852 5184 10908
rect 5184 10852 5188 10908
rect 5124 10848 5188 10852
rect 8817 10908 8881 10912
rect 8817 10852 8821 10908
rect 8821 10852 8877 10908
rect 8877 10852 8881 10908
rect 8817 10848 8881 10852
rect 8897 10908 8961 10912
rect 8897 10852 8901 10908
rect 8901 10852 8957 10908
rect 8957 10852 8961 10908
rect 8897 10848 8961 10852
rect 8977 10908 9041 10912
rect 8977 10852 8981 10908
rect 8981 10852 9037 10908
rect 9037 10852 9041 10908
rect 8977 10848 9041 10852
rect 9057 10908 9121 10912
rect 9057 10852 9061 10908
rect 9061 10852 9117 10908
rect 9117 10852 9121 10908
rect 9057 10848 9121 10852
rect 12750 10908 12814 10912
rect 12750 10852 12754 10908
rect 12754 10852 12810 10908
rect 12810 10852 12814 10908
rect 12750 10848 12814 10852
rect 12830 10908 12894 10912
rect 12830 10852 12834 10908
rect 12834 10852 12890 10908
rect 12890 10852 12894 10908
rect 12830 10848 12894 10852
rect 12910 10908 12974 10912
rect 12910 10852 12914 10908
rect 12914 10852 12970 10908
rect 12970 10852 12974 10908
rect 12910 10848 12974 10852
rect 12990 10908 13054 10912
rect 12990 10852 12994 10908
rect 12994 10852 13050 10908
rect 13050 10852 13054 10908
rect 12990 10848 13054 10852
rect 16683 10908 16747 10912
rect 16683 10852 16687 10908
rect 16687 10852 16743 10908
rect 16743 10852 16747 10908
rect 16683 10848 16747 10852
rect 16763 10908 16827 10912
rect 16763 10852 16767 10908
rect 16767 10852 16823 10908
rect 16823 10852 16827 10908
rect 16763 10848 16827 10852
rect 16843 10908 16907 10912
rect 16843 10852 16847 10908
rect 16847 10852 16903 10908
rect 16903 10852 16907 10908
rect 16843 10848 16907 10852
rect 16923 10908 16987 10912
rect 16923 10852 16927 10908
rect 16927 10852 16983 10908
rect 16983 10852 16987 10908
rect 16923 10848 16987 10852
rect 2918 10364 2982 10368
rect 2918 10308 2922 10364
rect 2922 10308 2978 10364
rect 2978 10308 2982 10364
rect 2918 10304 2982 10308
rect 2998 10364 3062 10368
rect 2998 10308 3002 10364
rect 3002 10308 3058 10364
rect 3058 10308 3062 10364
rect 2998 10304 3062 10308
rect 3078 10364 3142 10368
rect 3078 10308 3082 10364
rect 3082 10308 3138 10364
rect 3138 10308 3142 10364
rect 3078 10304 3142 10308
rect 3158 10364 3222 10368
rect 3158 10308 3162 10364
rect 3162 10308 3218 10364
rect 3218 10308 3222 10364
rect 3158 10304 3222 10308
rect 6851 10364 6915 10368
rect 6851 10308 6855 10364
rect 6855 10308 6911 10364
rect 6911 10308 6915 10364
rect 6851 10304 6915 10308
rect 6931 10364 6995 10368
rect 6931 10308 6935 10364
rect 6935 10308 6991 10364
rect 6991 10308 6995 10364
rect 6931 10304 6995 10308
rect 7011 10364 7075 10368
rect 7011 10308 7015 10364
rect 7015 10308 7071 10364
rect 7071 10308 7075 10364
rect 7011 10304 7075 10308
rect 7091 10364 7155 10368
rect 7091 10308 7095 10364
rect 7095 10308 7151 10364
rect 7151 10308 7155 10364
rect 7091 10304 7155 10308
rect 10784 10364 10848 10368
rect 10784 10308 10788 10364
rect 10788 10308 10844 10364
rect 10844 10308 10848 10364
rect 10784 10304 10848 10308
rect 10864 10364 10928 10368
rect 10864 10308 10868 10364
rect 10868 10308 10924 10364
rect 10924 10308 10928 10364
rect 10864 10304 10928 10308
rect 10944 10364 11008 10368
rect 10944 10308 10948 10364
rect 10948 10308 11004 10364
rect 11004 10308 11008 10364
rect 10944 10304 11008 10308
rect 11024 10364 11088 10368
rect 11024 10308 11028 10364
rect 11028 10308 11084 10364
rect 11084 10308 11088 10364
rect 11024 10304 11088 10308
rect 14717 10364 14781 10368
rect 14717 10308 14721 10364
rect 14721 10308 14777 10364
rect 14777 10308 14781 10364
rect 14717 10304 14781 10308
rect 14797 10364 14861 10368
rect 14797 10308 14801 10364
rect 14801 10308 14857 10364
rect 14857 10308 14861 10364
rect 14797 10304 14861 10308
rect 14877 10364 14941 10368
rect 14877 10308 14881 10364
rect 14881 10308 14937 10364
rect 14937 10308 14941 10364
rect 14877 10304 14941 10308
rect 14957 10364 15021 10368
rect 14957 10308 14961 10364
rect 14961 10308 15017 10364
rect 15017 10308 15021 10364
rect 14957 10304 15021 10308
rect 4884 9820 4948 9824
rect 4884 9764 4888 9820
rect 4888 9764 4944 9820
rect 4944 9764 4948 9820
rect 4884 9760 4948 9764
rect 4964 9820 5028 9824
rect 4964 9764 4968 9820
rect 4968 9764 5024 9820
rect 5024 9764 5028 9820
rect 4964 9760 5028 9764
rect 5044 9820 5108 9824
rect 5044 9764 5048 9820
rect 5048 9764 5104 9820
rect 5104 9764 5108 9820
rect 5044 9760 5108 9764
rect 5124 9820 5188 9824
rect 5124 9764 5128 9820
rect 5128 9764 5184 9820
rect 5184 9764 5188 9820
rect 5124 9760 5188 9764
rect 8817 9820 8881 9824
rect 8817 9764 8821 9820
rect 8821 9764 8877 9820
rect 8877 9764 8881 9820
rect 8817 9760 8881 9764
rect 8897 9820 8961 9824
rect 8897 9764 8901 9820
rect 8901 9764 8957 9820
rect 8957 9764 8961 9820
rect 8897 9760 8961 9764
rect 8977 9820 9041 9824
rect 8977 9764 8981 9820
rect 8981 9764 9037 9820
rect 9037 9764 9041 9820
rect 8977 9760 9041 9764
rect 9057 9820 9121 9824
rect 9057 9764 9061 9820
rect 9061 9764 9117 9820
rect 9117 9764 9121 9820
rect 9057 9760 9121 9764
rect 12750 9820 12814 9824
rect 12750 9764 12754 9820
rect 12754 9764 12810 9820
rect 12810 9764 12814 9820
rect 12750 9760 12814 9764
rect 12830 9820 12894 9824
rect 12830 9764 12834 9820
rect 12834 9764 12890 9820
rect 12890 9764 12894 9820
rect 12830 9760 12894 9764
rect 12910 9820 12974 9824
rect 12910 9764 12914 9820
rect 12914 9764 12970 9820
rect 12970 9764 12974 9820
rect 12910 9760 12974 9764
rect 12990 9820 13054 9824
rect 12990 9764 12994 9820
rect 12994 9764 13050 9820
rect 13050 9764 13054 9820
rect 12990 9760 13054 9764
rect 16683 9820 16747 9824
rect 16683 9764 16687 9820
rect 16687 9764 16743 9820
rect 16743 9764 16747 9820
rect 16683 9760 16747 9764
rect 16763 9820 16827 9824
rect 16763 9764 16767 9820
rect 16767 9764 16823 9820
rect 16823 9764 16827 9820
rect 16763 9760 16827 9764
rect 16843 9820 16907 9824
rect 16843 9764 16847 9820
rect 16847 9764 16903 9820
rect 16903 9764 16907 9820
rect 16843 9760 16907 9764
rect 16923 9820 16987 9824
rect 16923 9764 16927 9820
rect 16927 9764 16983 9820
rect 16983 9764 16987 9820
rect 16923 9760 16987 9764
rect 2918 9276 2982 9280
rect 2918 9220 2922 9276
rect 2922 9220 2978 9276
rect 2978 9220 2982 9276
rect 2918 9216 2982 9220
rect 2998 9276 3062 9280
rect 2998 9220 3002 9276
rect 3002 9220 3058 9276
rect 3058 9220 3062 9276
rect 2998 9216 3062 9220
rect 3078 9276 3142 9280
rect 3078 9220 3082 9276
rect 3082 9220 3138 9276
rect 3138 9220 3142 9276
rect 3078 9216 3142 9220
rect 3158 9276 3222 9280
rect 3158 9220 3162 9276
rect 3162 9220 3218 9276
rect 3218 9220 3222 9276
rect 3158 9216 3222 9220
rect 6851 9276 6915 9280
rect 6851 9220 6855 9276
rect 6855 9220 6911 9276
rect 6911 9220 6915 9276
rect 6851 9216 6915 9220
rect 6931 9276 6995 9280
rect 6931 9220 6935 9276
rect 6935 9220 6991 9276
rect 6991 9220 6995 9276
rect 6931 9216 6995 9220
rect 7011 9276 7075 9280
rect 7011 9220 7015 9276
rect 7015 9220 7071 9276
rect 7071 9220 7075 9276
rect 7011 9216 7075 9220
rect 7091 9276 7155 9280
rect 7091 9220 7095 9276
rect 7095 9220 7151 9276
rect 7151 9220 7155 9276
rect 7091 9216 7155 9220
rect 10784 9276 10848 9280
rect 10784 9220 10788 9276
rect 10788 9220 10844 9276
rect 10844 9220 10848 9276
rect 10784 9216 10848 9220
rect 10864 9276 10928 9280
rect 10864 9220 10868 9276
rect 10868 9220 10924 9276
rect 10924 9220 10928 9276
rect 10864 9216 10928 9220
rect 10944 9276 11008 9280
rect 10944 9220 10948 9276
rect 10948 9220 11004 9276
rect 11004 9220 11008 9276
rect 10944 9216 11008 9220
rect 11024 9276 11088 9280
rect 11024 9220 11028 9276
rect 11028 9220 11084 9276
rect 11084 9220 11088 9276
rect 11024 9216 11088 9220
rect 14717 9276 14781 9280
rect 14717 9220 14721 9276
rect 14721 9220 14777 9276
rect 14777 9220 14781 9276
rect 14717 9216 14781 9220
rect 14797 9276 14861 9280
rect 14797 9220 14801 9276
rect 14801 9220 14857 9276
rect 14857 9220 14861 9276
rect 14797 9216 14861 9220
rect 14877 9276 14941 9280
rect 14877 9220 14881 9276
rect 14881 9220 14937 9276
rect 14937 9220 14941 9276
rect 14877 9216 14941 9220
rect 14957 9276 15021 9280
rect 14957 9220 14961 9276
rect 14961 9220 15017 9276
rect 15017 9220 15021 9276
rect 14957 9216 15021 9220
rect 4884 8732 4948 8736
rect 4884 8676 4888 8732
rect 4888 8676 4944 8732
rect 4944 8676 4948 8732
rect 4884 8672 4948 8676
rect 4964 8732 5028 8736
rect 4964 8676 4968 8732
rect 4968 8676 5024 8732
rect 5024 8676 5028 8732
rect 4964 8672 5028 8676
rect 5044 8732 5108 8736
rect 5044 8676 5048 8732
rect 5048 8676 5104 8732
rect 5104 8676 5108 8732
rect 5044 8672 5108 8676
rect 5124 8732 5188 8736
rect 5124 8676 5128 8732
rect 5128 8676 5184 8732
rect 5184 8676 5188 8732
rect 5124 8672 5188 8676
rect 8817 8732 8881 8736
rect 8817 8676 8821 8732
rect 8821 8676 8877 8732
rect 8877 8676 8881 8732
rect 8817 8672 8881 8676
rect 8897 8732 8961 8736
rect 8897 8676 8901 8732
rect 8901 8676 8957 8732
rect 8957 8676 8961 8732
rect 8897 8672 8961 8676
rect 8977 8732 9041 8736
rect 8977 8676 8981 8732
rect 8981 8676 9037 8732
rect 9037 8676 9041 8732
rect 8977 8672 9041 8676
rect 9057 8732 9121 8736
rect 9057 8676 9061 8732
rect 9061 8676 9117 8732
rect 9117 8676 9121 8732
rect 9057 8672 9121 8676
rect 12750 8732 12814 8736
rect 12750 8676 12754 8732
rect 12754 8676 12810 8732
rect 12810 8676 12814 8732
rect 12750 8672 12814 8676
rect 12830 8732 12894 8736
rect 12830 8676 12834 8732
rect 12834 8676 12890 8732
rect 12890 8676 12894 8732
rect 12830 8672 12894 8676
rect 12910 8732 12974 8736
rect 12910 8676 12914 8732
rect 12914 8676 12970 8732
rect 12970 8676 12974 8732
rect 12910 8672 12974 8676
rect 12990 8732 13054 8736
rect 12990 8676 12994 8732
rect 12994 8676 13050 8732
rect 13050 8676 13054 8732
rect 12990 8672 13054 8676
rect 16683 8732 16747 8736
rect 16683 8676 16687 8732
rect 16687 8676 16743 8732
rect 16743 8676 16747 8732
rect 16683 8672 16747 8676
rect 16763 8732 16827 8736
rect 16763 8676 16767 8732
rect 16767 8676 16823 8732
rect 16823 8676 16827 8732
rect 16763 8672 16827 8676
rect 16843 8732 16907 8736
rect 16843 8676 16847 8732
rect 16847 8676 16903 8732
rect 16903 8676 16907 8732
rect 16843 8672 16907 8676
rect 16923 8732 16987 8736
rect 16923 8676 16927 8732
rect 16927 8676 16983 8732
rect 16983 8676 16987 8732
rect 16923 8672 16987 8676
rect 2918 8188 2982 8192
rect 2918 8132 2922 8188
rect 2922 8132 2978 8188
rect 2978 8132 2982 8188
rect 2918 8128 2982 8132
rect 2998 8188 3062 8192
rect 2998 8132 3002 8188
rect 3002 8132 3058 8188
rect 3058 8132 3062 8188
rect 2998 8128 3062 8132
rect 3078 8188 3142 8192
rect 3078 8132 3082 8188
rect 3082 8132 3138 8188
rect 3138 8132 3142 8188
rect 3078 8128 3142 8132
rect 3158 8188 3222 8192
rect 3158 8132 3162 8188
rect 3162 8132 3218 8188
rect 3218 8132 3222 8188
rect 3158 8128 3222 8132
rect 6851 8188 6915 8192
rect 6851 8132 6855 8188
rect 6855 8132 6911 8188
rect 6911 8132 6915 8188
rect 6851 8128 6915 8132
rect 6931 8188 6995 8192
rect 6931 8132 6935 8188
rect 6935 8132 6991 8188
rect 6991 8132 6995 8188
rect 6931 8128 6995 8132
rect 7011 8188 7075 8192
rect 7011 8132 7015 8188
rect 7015 8132 7071 8188
rect 7071 8132 7075 8188
rect 7011 8128 7075 8132
rect 7091 8188 7155 8192
rect 7091 8132 7095 8188
rect 7095 8132 7151 8188
rect 7151 8132 7155 8188
rect 7091 8128 7155 8132
rect 10784 8188 10848 8192
rect 10784 8132 10788 8188
rect 10788 8132 10844 8188
rect 10844 8132 10848 8188
rect 10784 8128 10848 8132
rect 10864 8188 10928 8192
rect 10864 8132 10868 8188
rect 10868 8132 10924 8188
rect 10924 8132 10928 8188
rect 10864 8128 10928 8132
rect 10944 8188 11008 8192
rect 10944 8132 10948 8188
rect 10948 8132 11004 8188
rect 11004 8132 11008 8188
rect 10944 8128 11008 8132
rect 11024 8188 11088 8192
rect 11024 8132 11028 8188
rect 11028 8132 11084 8188
rect 11084 8132 11088 8188
rect 11024 8128 11088 8132
rect 14717 8188 14781 8192
rect 14717 8132 14721 8188
rect 14721 8132 14777 8188
rect 14777 8132 14781 8188
rect 14717 8128 14781 8132
rect 14797 8188 14861 8192
rect 14797 8132 14801 8188
rect 14801 8132 14857 8188
rect 14857 8132 14861 8188
rect 14797 8128 14861 8132
rect 14877 8188 14941 8192
rect 14877 8132 14881 8188
rect 14881 8132 14937 8188
rect 14937 8132 14941 8188
rect 14877 8128 14941 8132
rect 14957 8188 15021 8192
rect 14957 8132 14961 8188
rect 14961 8132 15017 8188
rect 15017 8132 15021 8188
rect 14957 8128 15021 8132
rect 4884 7644 4948 7648
rect 4884 7588 4888 7644
rect 4888 7588 4944 7644
rect 4944 7588 4948 7644
rect 4884 7584 4948 7588
rect 4964 7644 5028 7648
rect 4964 7588 4968 7644
rect 4968 7588 5024 7644
rect 5024 7588 5028 7644
rect 4964 7584 5028 7588
rect 5044 7644 5108 7648
rect 5044 7588 5048 7644
rect 5048 7588 5104 7644
rect 5104 7588 5108 7644
rect 5044 7584 5108 7588
rect 5124 7644 5188 7648
rect 5124 7588 5128 7644
rect 5128 7588 5184 7644
rect 5184 7588 5188 7644
rect 5124 7584 5188 7588
rect 8817 7644 8881 7648
rect 8817 7588 8821 7644
rect 8821 7588 8877 7644
rect 8877 7588 8881 7644
rect 8817 7584 8881 7588
rect 8897 7644 8961 7648
rect 8897 7588 8901 7644
rect 8901 7588 8957 7644
rect 8957 7588 8961 7644
rect 8897 7584 8961 7588
rect 8977 7644 9041 7648
rect 8977 7588 8981 7644
rect 8981 7588 9037 7644
rect 9037 7588 9041 7644
rect 8977 7584 9041 7588
rect 9057 7644 9121 7648
rect 9057 7588 9061 7644
rect 9061 7588 9117 7644
rect 9117 7588 9121 7644
rect 9057 7584 9121 7588
rect 12750 7644 12814 7648
rect 12750 7588 12754 7644
rect 12754 7588 12810 7644
rect 12810 7588 12814 7644
rect 12750 7584 12814 7588
rect 12830 7644 12894 7648
rect 12830 7588 12834 7644
rect 12834 7588 12890 7644
rect 12890 7588 12894 7644
rect 12830 7584 12894 7588
rect 12910 7644 12974 7648
rect 12910 7588 12914 7644
rect 12914 7588 12970 7644
rect 12970 7588 12974 7644
rect 12910 7584 12974 7588
rect 12990 7644 13054 7648
rect 12990 7588 12994 7644
rect 12994 7588 13050 7644
rect 13050 7588 13054 7644
rect 12990 7584 13054 7588
rect 16683 7644 16747 7648
rect 16683 7588 16687 7644
rect 16687 7588 16743 7644
rect 16743 7588 16747 7644
rect 16683 7584 16747 7588
rect 16763 7644 16827 7648
rect 16763 7588 16767 7644
rect 16767 7588 16823 7644
rect 16823 7588 16827 7644
rect 16763 7584 16827 7588
rect 16843 7644 16907 7648
rect 16843 7588 16847 7644
rect 16847 7588 16903 7644
rect 16903 7588 16907 7644
rect 16843 7584 16907 7588
rect 16923 7644 16987 7648
rect 16923 7588 16927 7644
rect 16927 7588 16983 7644
rect 16983 7588 16987 7644
rect 16923 7584 16987 7588
rect 2918 7100 2982 7104
rect 2918 7044 2922 7100
rect 2922 7044 2978 7100
rect 2978 7044 2982 7100
rect 2918 7040 2982 7044
rect 2998 7100 3062 7104
rect 2998 7044 3002 7100
rect 3002 7044 3058 7100
rect 3058 7044 3062 7100
rect 2998 7040 3062 7044
rect 3078 7100 3142 7104
rect 3078 7044 3082 7100
rect 3082 7044 3138 7100
rect 3138 7044 3142 7100
rect 3078 7040 3142 7044
rect 3158 7100 3222 7104
rect 3158 7044 3162 7100
rect 3162 7044 3218 7100
rect 3218 7044 3222 7100
rect 3158 7040 3222 7044
rect 6851 7100 6915 7104
rect 6851 7044 6855 7100
rect 6855 7044 6911 7100
rect 6911 7044 6915 7100
rect 6851 7040 6915 7044
rect 6931 7100 6995 7104
rect 6931 7044 6935 7100
rect 6935 7044 6991 7100
rect 6991 7044 6995 7100
rect 6931 7040 6995 7044
rect 7011 7100 7075 7104
rect 7011 7044 7015 7100
rect 7015 7044 7071 7100
rect 7071 7044 7075 7100
rect 7011 7040 7075 7044
rect 7091 7100 7155 7104
rect 7091 7044 7095 7100
rect 7095 7044 7151 7100
rect 7151 7044 7155 7100
rect 7091 7040 7155 7044
rect 10784 7100 10848 7104
rect 10784 7044 10788 7100
rect 10788 7044 10844 7100
rect 10844 7044 10848 7100
rect 10784 7040 10848 7044
rect 10864 7100 10928 7104
rect 10864 7044 10868 7100
rect 10868 7044 10924 7100
rect 10924 7044 10928 7100
rect 10864 7040 10928 7044
rect 10944 7100 11008 7104
rect 10944 7044 10948 7100
rect 10948 7044 11004 7100
rect 11004 7044 11008 7100
rect 10944 7040 11008 7044
rect 11024 7100 11088 7104
rect 11024 7044 11028 7100
rect 11028 7044 11084 7100
rect 11084 7044 11088 7100
rect 11024 7040 11088 7044
rect 14717 7100 14781 7104
rect 14717 7044 14721 7100
rect 14721 7044 14777 7100
rect 14777 7044 14781 7100
rect 14717 7040 14781 7044
rect 14797 7100 14861 7104
rect 14797 7044 14801 7100
rect 14801 7044 14857 7100
rect 14857 7044 14861 7100
rect 14797 7040 14861 7044
rect 14877 7100 14941 7104
rect 14877 7044 14881 7100
rect 14881 7044 14937 7100
rect 14937 7044 14941 7100
rect 14877 7040 14941 7044
rect 14957 7100 15021 7104
rect 14957 7044 14961 7100
rect 14961 7044 15017 7100
rect 15017 7044 15021 7100
rect 14957 7040 15021 7044
rect 4884 6556 4948 6560
rect 4884 6500 4888 6556
rect 4888 6500 4944 6556
rect 4944 6500 4948 6556
rect 4884 6496 4948 6500
rect 4964 6556 5028 6560
rect 4964 6500 4968 6556
rect 4968 6500 5024 6556
rect 5024 6500 5028 6556
rect 4964 6496 5028 6500
rect 5044 6556 5108 6560
rect 5044 6500 5048 6556
rect 5048 6500 5104 6556
rect 5104 6500 5108 6556
rect 5044 6496 5108 6500
rect 5124 6556 5188 6560
rect 5124 6500 5128 6556
rect 5128 6500 5184 6556
rect 5184 6500 5188 6556
rect 5124 6496 5188 6500
rect 8817 6556 8881 6560
rect 8817 6500 8821 6556
rect 8821 6500 8877 6556
rect 8877 6500 8881 6556
rect 8817 6496 8881 6500
rect 8897 6556 8961 6560
rect 8897 6500 8901 6556
rect 8901 6500 8957 6556
rect 8957 6500 8961 6556
rect 8897 6496 8961 6500
rect 8977 6556 9041 6560
rect 8977 6500 8981 6556
rect 8981 6500 9037 6556
rect 9037 6500 9041 6556
rect 8977 6496 9041 6500
rect 9057 6556 9121 6560
rect 9057 6500 9061 6556
rect 9061 6500 9117 6556
rect 9117 6500 9121 6556
rect 9057 6496 9121 6500
rect 12750 6556 12814 6560
rect 12750 6500 12754 6556
rect 12754 6500 12810 6556
rect 12810 6500 12814 6556
rect 12750 6496 12814 6500
rect 12830 6556 12894 6560
rect 12830 6500 12834 6556
rect 12834 6500 12890 6556
rect 12890 6500 12894 6556
rect 12830 6496 12894 6500
rect 12910 6556 12974 6560
rect 12910 6500 12914 6556
rect 12914 6500 12970 6556
rect 12970 6500 12974 6556
rect 12910 6496 12974 6500
rect 12990 6556 13054 6560
rect 12990 6500 12994 6556
rect 12994 6500 13050 6556
rect 13050 6500 13054 6556
rect 12990 6496 13054 6500
rect 16683 6556 16747 6560
rect 16683 6500 16687 6556
rect 16687 6500 16743 6556
rect 16743 6500 16747 6556
rect 16683 6496 16747 6500
rect 16763 6556 16827 6560
rect 16763 6500 16767 6556
rect 16767 6500 16823 6556
rect 16823 6500 16827 6556
rect 16763 6496 16827 6500
rect 16843 6556 16907 6560
rect 16843 6500 16847 6556
rect 16847 6500 16903 6556
rect 16903 6500 16907 6556
rect 16843 6496 16907 6500
rect 16923 6556 16987 6560
rect 16923 6500 16927 6556
rect 16927 6500 16983 6556
rect 16983 6500 16987 6556
rect 16923 6496 16987 6500
rect 2918 6012 2982 6016
rect 2918 5956 2922 6012
rect 2922 5956 2978 6012
rect 2978 5956 2982 6012
rect 2918 5952 2982 5956
rect 2998 6012 3062 6016
rect 2998 5956 3002 6012
rect 3002 5956 3058 6012
rect 3058 5956 3062 6012
rect 2998 5952 3062 5956
rect 3078 6012 3142 6016
rect 3078 5956 3082 6012
rect 3082 5956 3138 6012
rect 3138 5956 3142 6012
rect 3078 5952 3142 5956
rect 3158 6012 3222 6016
rect 3158 5956 3162 6012
rect 3162 5956 3218 6012
rect 3218 5956 3222 6012
rect 3158 5952 3222 5956
rect 6851 6012 6915 6016
rect 6851 5956 6855 6012
rect 6855 5956 6911 6012
rect 6911 5956 6915 6012
rect 6851 5952 6915 5956
rect 6931 6012 6995 6016
rect 6931 5956 6935 6012
rect 6935 5956 6991 6012
rect 6991 5956 6995 6012
rect 6931 5952 6995 5956
rect 7011 6012 7075 6016
rect 7011 5956 7015 6012
rect 7015 5956 7071 6012
rect 7071 5956 7075 6012
rect 7011 5952 7075 5956
rect 7091 6012 7155 6016
rect 7091 5956 7095 6012
rect 7095 5956 7151 6012
rect 7151 5956 7155 6012
rect 7091 5952 7155 5956
rect 10784 6012 10848 6016
rect 10784 5956 10788 6012
rect 10788 5956 10844 6012
rect 10844 5956 10848 6012
rect 10784 5952 10848 5956
rect 10864 6012 10928 6016
rect 10864 5956 10868 6012
rect 10868 5956 10924 6012
rect 10924 5956 10928 6012
rect 10864 5952 10928 5956
rect 10944 6012 11008 6016
rect 10944 5956 10948 6012
rect 10948 5956 11004 6012
rect 11004 5956 11008 6012
rect 10944 5952 11008 5956
rect 11024 6012 11088 6016
rect 11024 5956 11028 6012
rect 11028 5956 11084 6012
rect 11084 5956 11088 6012
rect 11024 5952 11088 5956
rect 14717 6012 14781 6016
rect 14717 5956 14721 6012
rect 14721 5956 14777 6012
rect 14777 5956 14781 6012
rect 14717 5952 14781 5956
rect 14797 6012 14861 6016
rect 14797 5956 14801 6012
rect 14801 5956 14857 6012
rect 14857 5956 14861 6012
rect 14797 5952 14861 5956
rect 14877 6012 14941 6016
rect 14877 5956 14881 6012
rect 14881 5956 14937 6012
rect 14937 5956 14941 6012
rect 14877 5952 14941 5956
rect 14957 6012 15021 6016
rect 14957 5956 14961 6012
rect 14961 5956 15017 6012
rect 15017 5956 15021 6012
rect 14957 5952 15021 5956
rect 4884 5468 4948 5472
rect 4884 5412 4888 5468
rect 4888 5412 4944 5468
rect 4944 5412 4948 5468
rect 4884 5408 4948 5412
rect 4964 5468 5028 5472
rect 4964 5412 4968 5468
rect 4968 5412 5024 5468
rect 5024 5412 5028 5468
rect 4964 5408 5028 5412
rect 5044 5468 5108 5472
rect 5044 5412 5048 5468
rect 5048 5412 5104 5468
rect 5104 5412 5108 5468
rect 5044 5408 5108 5412
rect 5124 5468 5188 5472
rect 5124 5412 5128 5468
rect 5128 5412 5184 5468
rect 5184 5412 5188 5468
rect 5124 5408 5188 5412
rect 8817 5468 8881 5472
rect 8817 5412 8821 5468
rect 8821 5412 8877 5468
rect 8877 5412 8881 5468
rect 8817 5408 8881 5412
rect 8897 5468 8961 5472
rect 8897 5412 8901 5468
rect 8901 5412 8957 5468
rect 8957 5412 8961 5468
rect 8897 5408 8961 5412
rect 8977 5468 9041 5472
rect 8977 5412 8981 5468
rect 8981 5412 9037 5468
rect 9037 5412 9041 5468
rect 8977 5408 9041 5412
rect 9057 5468 9121 5472
rect 9057 5412 9061 5468
rect 9061 5412 9117 5468
rect 9117 5412 9121 5468
rect 9057 5408 9121 5412
rect 12750 5468 12814 5472
rect 12750 5412 12754 5468
rect 12754 5412 12810 5468
rect 12810 5412 12814 5468
rect 12750 5408 12814 5412
rect 12830 5468 12894 5472
rect 12830 5412 12834 5468
rect 12834 5412 12890 5468
rect 12890 5412 12894 5468
rect 12830 5408 12894 5412
rect 12910 5468 12974 5472
rect 12910 5412 12914 5468
rect 12914 5412 12970 5468
rect 12970 5412 12974 5468
rect 12910 5408 12974 5412
rect 12990 5468 13054 5472
rect 12990 5412 12994 5468
rect 12994 5412 13050 5468
rect 13050 5412 13054 5468
rect 12990 5408 13054 5412
rect 16683 5468 16747 5472
rect 16683 5412 16687 5468
rect 16687 5412 16743 5468
rect 16743 5412 16747 5468
rect 16683 5408 16747 5412
rect 16763 5468 16827 5472
rect 16763 5412 16767 5468
rect 16767 5412 16823 5468
rect 16823 5412 16827 5468
rect 16763 5408 16827 5412
rect 16843 5468 16907 5472
rect 16843 5412 16847 5468
rect 16847 5412 16903 5468
rect 16903 5412 16907 5468
rect 16843 5408 16907 5412
rect 16923 5468 16987 5472
rect 16923 5412 16927 5468
rect 16927 5412 16983 5468
rect 16983 5412 16987 5468
rect 16923 5408 16987 5412
rect 2918 4924 2982 4928
rect 2918 4868 2922 4924
rect 2922 4868 2978 4924
rect 2978 4868 2982 4924
rect 2918 4864 2982 4868
rect 2998 4924 3062 4928
rect 2998 4868 3002 4924
rect 3002 4868 3058 4924
rect 3058 4868 3062 4924
rect 2998 4864 3062 4868
rect 3078 4924 3142 4928
rect 3078 4868 3082 4924
rect 3082 4868 3138 4924
rect 3138 4868 3142 4924
rect 3078 4864 3142 4868
rect 3158 4924 3222 4928
rect 3158 4868 3162 4924
rect 3162 4868 3218 4924
rect 3218 4868 3222 4924
rect 3158 4864 3222 4868
rect 6851 4924 6915 4928
rect 6851 4868 6855 4924
rect 6855 4868 6911 4924
rect 6911 4868 6915 4924
rect 6851 4864 6915 4868
rect 6931 4924 6995 4928
rect 6931 4868 6935 4924
rect 6935 4868 6991 4924
rect 6991 4868 6995 4924
rect 6931 4864 6995 4868
rect 7011 4924 7075 4928
rect 7011 4868 7015 4924
rect 7015 4868 7071 4924
rect 7071 4868 7075 4924
rect 7011 4864 7075 4868
rect 7091 4924 7155 4928
rect 7091 4868 7095 4924
rect 7095 4868 7151 4924
rect 7151 4868 7155 4924
rect 7091 4864 7155 4868
rect 10784 4924 10848 4928
rect 10784 4868 10788 4924
rect 10788 4868 10844 4924
rect 10844 4868 10848 4924
rect 10784 4864 10848 4868
rect 10864 4924 10928 4928
rect 10864 4868 10868 4924
rect 10868 4868 10924 4924
rect 10924 4868 10928 4924
rect 10864 4864 10928 4868
rect 10944 4924 11008 4928
rect 10944 4868 10948 4924
rect 10948 4868 11004 4924
rect 11004 4868 11008 4924
rect 10944 4864 11008 4868
rect 11024 4924 11088 4928
rect 11024 4868 11028 4924
rect 11028 4868 11084 4924
rect 11084 4868 11088 4924
rect 11024 4864 11088 4868
rect 14717 4924 14781 4928
rect 14717 4868 14721 4924
rect 14721 4868 14777 4924
rect 14777 4868 14781 4924
rect 14717 4864 14781 4868
rect 14797 4924 14861 4928
rect 14797 4868 14801 4924
rect 14801 4868 14857 4924
rect 14857 4868 14861 4924
rect 14797 4864 14861 4868
rect 14877 4924 14941 4928
rect 14877 4868 14881 4924
rect 14881 4868 14937 4924
rect 14937 4868 14941 4924
rect 14877 4864 14941 4868
rect 14957 4924 15021 4928
rect 14957 4868 14961 4924
rect 14961 4868 15017 4924
rect 15017 4868 15021 4924
rect 14957 4864 15021 4868
rect 4884 4380 4948 4384
rect 4884 4324 4888 4380
rect 4888 4324 4944 4380
rect 4944 4324 4948 4380
rect 4884 4320 4948 4324
rect 4964 4380 5028 4384
rect 4964 4324 4968 4380
rect 4968 4324 5024 4380
rect 5024 4324 5028 4380
rect 4964 4320 5028 4324
rect 5044 4380 5108 4384
rect 5044 4324 5048 4380
rect 5048 4324 5104 4380
rect 5104 4324 5108 4380
rect 5044 4320 5108 4324
rect 5124 4380 5188 4384
rect 5124 4324 5128 4380
rect 5128 4324 5184 4380
rect 5184 4324 5188 4380
rect 5124 4320 5188 4324
rect 8817 4380 8881 4384
rect 8817 4324 8821 4380
rect 8821 4324 8877 4380
rect 8877 4324 8881 4380
rect 8817 4320 8881 4324
rect 8897 4380 8961 4384
rect 8897 4324 8901 4380
rect 8901 4324 8957 4380
rect 8957 4324 8961 4380
rect 8897 4320 8961 4324
rect 8977 4380 9041 4384
rect 8977 4324 8981 4380
rect 8981 4324 9037 4380
rect 9037 4324 9041 4380
rect 8977 4320 9041 4324
rect 9057 4380 9121 4384
rect 9057 4324 9061 4380
rect 9061 4324 9117 4380
rect 9117 4324 9121 4380
rect 9057 4320 9121 4324
rect 12750 4380 12814 4384
rect 12750 4324 12754 4380
rect 12754 4324 12810 4380
rect 12810 4324 12814 4380
rect 12750 4320 12814 4324
rect 12830 4380 12894 4384
rect 12830 4324 12834 4380
rect 12834 4324 12890 4380
rect 12890 4324 12894 4380
rect 12830 4320 12894 4324
rect 12910 4380 12974 4384
rect 12910 4324 12914 4380
rect 12914 4324 12970 4380
rect 12970 4324 12974 4380
rect 12910 4320 12974 4324
rect 12990 4380 13054 4384
rect 12990 4324 12994 4380
rect 12994 4324 13050 4380
rect 13050 4324 13054 4380
rect 12990 4320 13054 4324
rect 16683 4380 16747 4384
rect 16683 4324 16687 4380
rect 16687 4324 16743 4380
rect 16743 4324 16747 4380
rect 16683 4320 16747 4324
rect 16763 4380 16827 4384
rect 16763 4324 16767 4380
rect 16767 4324 16823 4380
rect 16823 4324 16827 4380
rect 16763 4320 16827 4324
rect 16843 4380 16907 4384
rect 16843 4324 16847 4380
rect 16847 4324 16903 4380
rect 16903 4324 16907 4380
rect 16843 4320 16907 4324
rect 16923 4380 16987 4384
rect 16923 4324 16927 4380
rect 16927 4324 16983 4380
rect 16983 4324 16987 4380
rect 16923 4320 16987 4324
rect 2918 3836 2982 3840
rect 2918 3780 2922 3836
rect 2922 3780 2978 3836
rect 2978 3780 2982 3836
rect 2918 3776 2982 3780
rect 2998 3836 3062 3840
rect 2998 3780 3002 3836
rect 3002 3780 3058 3836
rect 3058 3780 3062 3836
rect 2998 3776 3062 3780
rect 3078 3836 3142 3840
rect 3078 3780 3082 3836
rect 3082 3780 3138 3836
rect 3138 3780 3142 3836
rect 3078 3776 3142 3780
rect 3158 3836 3222 3840
rect 3158 3780 3162 3836
rect 3162 3780 3218 3836
rect 3218 3780 3222 3836
rect 3158 3776 3222 3780
rect 6851 3836 6915 3840
rect 6851 3780 6855 3836
rect 6855 3780 6911 3836
rect 6911 3780 6915 3836
rect 6851 3776 6915 3780
rect 6931 3836 6995 3840
rect 6931 3780 6935 3836
rect 6935 3780 6991 3836
rect 6991 3780 6995 3836
rect 6931 3776 6995 3780
rect 7011 3836 7075 3840
rect 7011 3780 7015 3836
rect 7015 3780 7071 3836
rect 7071 3780 7075 3836
rect 7011 3776 7075 3780
rect 7091 3836 7155 3840
rect 7091 3780 7095 3836
rect 7095 3780 7151 3836
rect 7151 3780 7155 3836
rect 7091 3776 7155 3780
rect 10784 3836 10848 3840
rect 10784 3780 10788 3836
rect 10788 3780 10844 3836
rect 10844 3780 10848 3836
rect 10784 3776 10848 3780
rect 10864 3836 10928 3840
rect 10864 3780 10868 3836
rect 10868 3780 10924 3836
rect 10924 3780 10928 3836
rect 10864 3776 10928 3780
rect 10944 3836 11008 3840
rect 10944 3780 10948 3836
rect 10948 3780 11004 3836
rect 11004 3780 11008 3836
rect 10944 3776 11008 3780
rect 11024 3836 11088 3840
rect 11024 3780 11028 3836
rect 11028 3780 11084 3836
rect 11084 3780 11088 3836
rect 11024 3776 11088 3780
rect 14717 3836 14781 3840
rect 14717 3780 14721 3836
rect 14721 3780 14777 3836
rect 14777 3780 14781 3836
rect 14717 3776 14781 3780
rect 14797 3836 14861 3840
rect 14797 3780 14801 3836
rect 14801 3780 14857 3836
rect 14857 3780 14861 3836
rect 14797 3776 14861 3780
rect 14877 3836 14941 3840
rect 14877 3780 14881 3836
rect 14881 3780 14937 3836
rect 14937 3780 14941 3836
rect 14877 3776 14941 3780
rect 14957 3836 15021 3840
rect 14957 3780 14961 3836
rect 14961 3780 15017 3836
rect 15017 3780 15021 3836
rect 14957 3776 15021 3780
rect 4884 3292 4948 3296
rect 4884 3236 4888 3292
rect 4888 3236 4944 3292
rect 4944 3236 4948 3292
rect 4884 3232 4948 3236
rect 4964 3292 5028 3296
rect 4964 3236 4968 3292
rect 4968 3236 5024 3292
rect 5024 3236 5028 3292
rect 4964 3232 5028 3236
rect 5044 3292 5108 3296
rect 5044 3236 5048 3292
rect 5048 3236 5104 3292
rect 5104 3236 5108 3292
rect 5044 3232 5108 3236
rect 5124 3292 5188 3296
rect 5124 3236 5128 3292
rect 5128 3236 5184 3292
rect 5184 3236 5188 3292
rect 5124 3232 5188 3236
rect 8817 3292 8881 3296
rect 8817 3236 8821 3292
rect 8821 3236 8877 3292
rect 8877 3236 8881 3292
rect 8817 3232 8881 3236
rect 8897 3292 8961 3296
rect 8897 3236 8901 3292
rect 8901 3236 8957 3292
rect 8957 3236 8961 3292
rect 8897 3232 8961 3236
rect 8977 3292 9041 3296
rect 8977 3236 8981 3292
rect 8981 3236 9037 3292
rect 9037 3236 9041 3292
rect 8977 3232 9041 3236
rect 9057 3292 9121 3296
rect 9057 3236 9061 3292
rect 9061 3236 9117 3292
rect 9117 3236 9121 3292
rect 9057 3232 9121 3236
rect 12750 3292 12814 3296
rect 12750 3236 12754 3292
rect 12754 3236 12810 3292
rect 12810 3236 12814 3292
rect 12750 3232 12814 3236
rect 12830 3292 12894 3296
rect 12830 3236 12834 3292
rect 12834 3236 12890 3292
rect 12890 3236 12894 3292
rect 12830 3232 12894 3236
rect 12910 3292 12974 3296
rect 12910 3236 12914 3292
rect 12914 3236 12970 3292
rect 12970 3236 12974 3292
rect 12910 3232 12974 3236
rect 12990 3292 13054 3296
rect 12990 3236 12994 3292
rect 12994 3236 13050 3292
rect 13050 3236 13054 3292
rect 12990 3232 13054 3236
rect 16683 3292 16747 3296
rect 16683 3236 16687 3292
rect 16687 3236 16743 3292
rect 16743 3236 16747 3292
rect 16683 3232 16747 3236
rect 16763 3292 16827 3296
rect 16763 3236 16767 3292
rect 16767 3236 16823 3292
rect 16823 3236 16827 3292
rect 16763 3232 16827 3236
rect 16843 3292 16907 3296
rect 16843 3236 16847 3292
rect 16847 3236 16903 3292
rect 16903 3236 16907 3292
rect 16843 3232 16907 3236
rect 16923 3292 16987 3296
rect 16923 3236 16927 3292
rect 16927 3236 16983 3292
rect 16983 3236 16987 3292
rect 16923 3232 16987 3236
rect 2918 2748 2982 2752
rect 2918 2692 2922 2748
rect 2922 2692 2978 2748
rect 2978 2692 2982 2748
rect 2918 2688 2982 2692
rect 2998 2748 3062 2752
rect 2998 2692 3002 2748
rect 3002 2692 3058 2748
rect 3058 2692 3062 2748
rect 2998 2688 3062 2692
rect 3078 2748 3142 2752
rect 3078 2692 3082 2748
rect 3082 2692 3138 2748
rect 3138 2692 3142 2748
rect 3078 2688 3142 2692
rect 3158 2748 3222 2752
rect 3158 2692 3162 2748
rect 3162 2692 3218 2748
rect 3218 2692 3222 2748
rect 3158 2688 3222 2692
rect 6851 2748 6915 2752
rect 6851 2692 6855 2748
rect 6855 2692 6911 2748
rect 6911 2692 6915 2748
rect 6851 2688 6915 2692
rect 6931 2748 6995 2752
rect 6931 2692 6935 2748
rect 6935 2692 6991 2748
rect 6991 2692 6995 2748
rect 6931 2688 6995 2692
rect 7011 2748 7075 2752
rect 7011 2692 7015 2748
rect 7015 2692 7071 2748
rect 7071 2692 7075 2748
rect 7011 2688 7075 2692
rect 7091 2748 7155 2752
rect 7091 2692 7095 2748
rect 7095 2692 7151 2748
rect 7151 2692 7155 2748
rect 7091 2688 7155 2692
rect 10784 2748 10848 2752
rect 10784 2692 10788 2748
rect 10788 2692 10844 2748
rect 10844 2692 10848 2748
rect 10784 2688 10848 2692
rect 10864 2748 10928 2752
rect 10864 2692 10868 2748
rect 10868 2692 10924 2748
rect 10924 2692 10928 2748
rect 10864 2688 10928 2692
rect 10944 2748 11008 2752
rect 10944 2692 10948 2748
rect 10948 2692 11004 2748
rect 11004 2692 11008 2748
rect 10944 2688 11008 2692
rect 11024 2748 11088 2752
rect 11024 2692 11028 2748
rect 11028 2692 11084 2748
rect 11084 2692 11088 2748
rect 11024 2688 11088 2692
rect 14717 2748 14781 2752
rect 14717 2692 14721 2748
rect 14721 2692 14777 2748
rect 14777 2692 14781 2748
rect 14717 2688 14781 2692
rect 14797 2748 14861 2752
rect 14797 2692 14801 2748
rect 14801 2692 14857 2748
rect 14857 2692 14861 2748
rect 14797 2688 14861 2692
rect 14877 2748 14941 2752
rect 14877 2692 14881 2748
rect 14881 2692 14937 2748
rect 14937 2692 14941 2748
rect 14877 2688 14941 2692
rect 14957 2748 15021 2752
rect 14957 2692 14961 2748
rect 14961 2692 15017 2748
rect 15017 2692 15021 2748
rect 14957 2688 15021 2692
rect 4884 2204 4948 2208
rect 4884 2148 4888 2204
rect 4888 2148 4944 2204
rect 4944 2148 4948 2204
rect 4884 2144 4948 2148
rect 4964 2204 5028 2208
rect 4964 2148 4968 2204
rect 4968 2148 5024 2204
rect 5024 2148 5028 2204
rect 4964 2144 5028 2148
rect 5044 2204 5108 2208
rect 5044 2148 5048 2204
rect 5048 2148 5104 2204
rect 5104 2148 5108 2204
rect 5044 2144 5108 2148
rect 5124 2204 5188 2208
rect 5124 2148 5128 2204
rect 5128 2148 5184 2204
rect 5184 2148 5188 2204
rect 5124 2144 5188 2148
rect 8817 2204 8881 2208
rect 8817 2148 8821 2204
rect 8821 2148 8877 2204
rect 8877 2148 8881 2204
rect 8817 2144 8881 2148
rect 8897 2204 8961 2208
rect 8897 2148 8901 2204
rect 8901 2148 8957 2204
rect 8957 2148 8961 2204
rect 8897 2144 8961 2148
rect 8977 2204 9041 2208
rect 8977 2148 8981 2204
rect 8981 2148 9037 2204
rect 9037 2148 9041 2204
rect 8977 2144 9041 2148
rect 9057 2204 9121 2208
rect 9057 2148 9061 2204
rect 9061 2148 9117 2204
rect 9117 2148 9121 2204
rect 9057 2144 9121 2148
rect 12750 2204 12814 2208
rect 12750 2148 12754 2204
rect 12754 2148 12810 2204
rect 12810 2148 12814 2204
rect 12750 2144 12814 2148
rect 12830 2204 12894 2208
rect 12830 2148 12834 2204
rect 12834 2148 12890 2204
rect 12890 2148 12894 2204
rect 12830 2144 12894 2148
rect 12910 2204 12974 2208
rect 12910 2148 12914 2204
rect 12914 2148 12970 2204
rect 12970 2148 12974 2204
rect 12910 2144 12974 2148
rect 12990 2204 13054 2208
rect 12990 2148 12994 2204
rect 12994 2148 13050 2204
rect 13050 2148 13054 2204
rect 12990 2144 13054 2148
rect 16683 2204 16747 2208
rect 16683 2148 16687 2204
rect 16687 2148 16743 2204
rect 16743 2148 16747 2204
rect 16683 2144 16747 2148
rect 16763 2204 16827 2208
rect 16763 2148 16767 2204
rect 16767 2148 16823 2204
rect 16823 2148 16827 2204
rect 16763 2144 16827 2148
rect 16843 2204 16907 2208
rect 16843 2148 16847 2204
rect 16847 2148 16903 2204
rect 16903 2148 16907 2204
rect 16843 2144 16907 2148
rect 16923 2204 16987 2208
rect 16923 2148 16927 2204
rect 16927 2148 16983 2204
rect 16983 2148 16987 2204
rect 16923 2144 16987 2148
<< metal4 >>
rect 2910 15808 3230 15824
rect 2910 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3230 15808
rect 2910 14720 3230 15744
rect 2910 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3230 14720
rect 2910 13632 3230 14656
rect 2910 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3230 13632
rect 2910 12544 3230 13568
rect 2910 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3230 12544
rect 2910 11456 3230 12480
rect 2910 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3230 11456
rect 2910 10368 3230 11392
rect 2910 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3230 10368
rect 2910 9280 3230 10304
rect 2910 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3230 9280
rect 2910 8192 3230 9216
rect 2910 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3230 8192
rect 2910 7104 3230 8128
rect 2910 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3230 7104
rect 2910 6016 3230 7040
rect 2910 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3230 6016
rect 2910 4928 3230 5952
rect 2910 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3230 4928
rect 2910 3840 3230 4864
rect 2910 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3230 3840
rect 2910 2752 3230 3776
rect 2910 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3230 2752
rect 2910 2128 3230 2688
rect 4876 15264 5196 15824
rect 4876 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5196 15264
rect 4876 14176 5196 15200
rect 4876 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5196 14176
rect 4876 13088 5196 14112
rect 4876 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5196 13088
rect 4876 12000 5196 13024
rect 4876 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5196 12000
rect 4876 10912 5196 11936
rect 4876 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5196 10912
rect 4876 9824 5196 10848
rect 4876 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5196 9824
rect 4876 8736 5196 9760
rect 4876 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5196 8736
rect 4876 7648 5196 8672
rect 4876 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5196 7648
rect 4876 6560 5196 7584
rect 4876 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5196 6560
rect 4876 5472 5196 6496
rect 4876 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5196 5472
rect 4876 4384 5196 5408
rect 4876 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5196 4384
rect 4876 3296 5196 4320
rect 4876 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5196 3296
rect 4876 2208 5196 3232
rect 4876 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5196 2208
rect 4876 2128 5196 2144
rect 6843 15808 7163 15824
rect 6843 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7163 15808
rect 6843 14720 7163 15744
rect 6843 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7163 14720
rect 6843 13632 7163 14656
rect 6843 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7163 13632
rect 6843 12544 7163 13568
rect 6843 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7163 12544
rect 6843 11456 7163 12480
rect 6843 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7163 11456
rect 6843 10368 7163 11392
rect 6843 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7163 10368
rect 6843 9280 7163 10304
rect 6843 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7163 9280
rect 6843 8192 7163 9216
rect 6843 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7163 8192
rect 6843 7104 7163 8128
rect 6843 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7163 7104
rect 6843 6016 7163 7040
rect 6843 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7163 6016
rect 6843 4928 7163 5952
rect 6843 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7163 4928
rect 6843 3840 7163 4864
rect 6843 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7163 3840
rect 6843 2752 7163 3776
rect 6843 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7163 2752
rect 6843 2128 7163 2688
rect 8809 15264 9129 15824
rect 8809 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9129 15264
rect 8809 14176 9129 15200
rect 8809 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9129 14176
rect 8809 13088 9129 14112
rect 8809 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9129 13088
rect 8809 12000 9129 13024
rect 8809 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9129 12000
rect 8809 10912 9129 11936
rect 8809 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9129 10912
rect 8809 9824 9129 10848
rect 8809 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9129 9824
rect 8809 8736 9129 9760
rect 8809 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9129 8736
rect 8809 7648 9129 8672
rect 8809 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9129 7648
rect 8809 6560 9129 7584
rect 8809 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9129 6560
rect 8809 5472 9129 6496
rect 8809 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9129 5472
rect 8809 4384 9129 5408
rect 8809 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9129 4384
rect 8809 3296 9129 4320
rect 8809 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9129 3296
rect 8809 2208 9129 3232
rect 8809 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9129 2208
rect 8809 2128 9129 2144
rect 10776 15808 11096 15824
rect 10776 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11096 15808
rect 10776 14720 11096 15744
rect 10776 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11096 14720
rect 10776 13632 11096 14656
rect 10776 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11096 13632
rect 10776 12544 11096 13568
rect 10776 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11096 12544
rect 10776 11456 11096 12480
rect 10776 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11096 11456
rect 10776 10368 11096 11392
rect 10776 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11096 10368
rect 10776 9280 11096 10304
rect 10776 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11096 9280
rect 10776 8192 11096 9216
rect 10776 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11096 8192
rect 10776 7104 11096 8128
rect 10776 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11096 7104
rect 10776 6016 11096 7040
rect 10776 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11096 6016
rect 10776 4928 11096 5952
rect 10776 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11096 4928
rect 10776 3840 11096 4864
rect 10776 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11096 3840
rect 10776 2752 11096 3776
rect 10776 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11096 2752
rect 10776 2128 11096 2688
rect 12742 15264 13062 15824
rect 12742 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13062 15264
rect 12742 14176 13062 15200
rect 12742 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13062 14176
rect 12742 13088 13062 14112
rect 12742 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13062 13088
rect 12742 12000 13062 13024
rect 12742 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13062 12000
rect 12742 10912 13062 11936
rect 12742 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13062 10912
rect 12742 9824 13062 10848
rect 12742 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13062 9824
rect 12742 8736 13062 9760
rect 12742 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13062 8736
rect 12742 7648 13062 8672
rect 12742 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13062 7648
rect 12742 6560 13062 7584
rect 12742 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13062 6560
rect 12742 5472 13062 6496
rect 12742 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13062 5472
rect 12742 4384 13062 5408
rect 12742 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13062 4384
rect 12742 3296 13062 4320
rect 12742 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13062 3296
rect 12742 2208 13062 3232
rect 12742 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13062 2208
rect 12742 2128 13062 2144
rect 14709 15808 15029 15824
rect 14709 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15029 15808
rect 14709 14720 15029 15744
rect 14709 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15029 14720
rect 14709 13632 15029 14656
rect 14709 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15029 13632
rect 14709 12544 15029 13568
rect 14709 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15029 12544
rect 14709 11456 15029 12480
rect 14709 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15029 11456
rect 14709 10368 15029 11392
rect 14709 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15029 10368
rect 14709 9280 15029 10304
rect 14709 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15029 9280
rect 14709 8192 15029 9216
rect 14709 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15029 8192
rect 14709 7104 15029 8128
rect 14709 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15029 7104
rect 14709 6016 15029 7040
rect 14709 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15029 6016
rect 14709 4928 15029 5952
rect 14709 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15029 4928
rect 14709 3840 15029 4864
rect 14709 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15029 3840
rect 14709 2752 15029 3776
rect 14709 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15029 2752
rect 14709 2128 15029 2688
rect 16675 15264 16995 15824
rect 16675 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16995 15264
rect 16675 14176 16995 15200
rect 16675 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16995 14176
rect 16675 13088 16995 14112
rect 16675 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16995 13088
rect 16675 12000 16995 13024
rect 16675 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16995 12000
rect 16675 10912 16995 11936
rect 16675 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16995 10912
rect 16675 9824 16995 10848
rect 16675 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16995 9824
rect 16675 8736 16995 9760
rect 16675 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16995 8736
rect 16675 7648 16995 8672
rect 16675 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16995 7648
rect 16675 6560 16995 7584
rect 16675 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16995 6560
rect 16675 5472 16995 6496
rect 16675 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16995 5472
rect 16675 4384 16995 5408
rect 16675 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16995 4384
rect 16675 3296 16995 4320
rect 16675 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16995 3296
rect 16675 2208 16995 3232
rect 16675 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16995 2208
rect 16675 2128 16995 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1676037725
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1676037725
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_74
timestamp 1676037725
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1676037725
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1676037725
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1676037725
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_16
timestamp 1676037725
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1676037725
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1676037725
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1676037725
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1676037725
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1676037725
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1676037725
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1676037725
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_94
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1676037725
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1676037725
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1676037725
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_50
timestamp 1676037725
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1676037725
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1676037725
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1676037725
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_92
timestamp 1676037725
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_104
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp 1676037725
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_132
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_157
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_166
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1676037725
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_31
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1676037725
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_98
timestamp 1676037725
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_92
timestamp 1676037725
transform 1 0 9568 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_104
timestamp 1676037725
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_116
timestamp 1676037725
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_128
timestamp 1676037725
transform 1 0 12880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_148
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_160
timestamp 1676037725
transform 1 0 15824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 1676037725
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1676037725
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1676037725
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1676037725
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1676037725
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_72
timestamp 1676037725
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1676037725
transform 1 0 11960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1676037725
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1676037725
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1676037725
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1676037725
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1676037725
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1676037725
transform 1 0 7360 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1676037725
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1676037725
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1676037725
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1676037725
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1676037725
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1676037725
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1676037725
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1676037725
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_50
timestamp 1676037725
transform 1 0 5704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1676037725
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_118
timestamp 1676037725
transform 1 0 11960 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_130
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_145
timestamp 1676037725
transform 1 0 14444 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_34
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_42
timestamp 1676037725
transform 1 0 4968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_75
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_92
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_17
timestamp 1676037725
transform 1 0 2668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1676037725
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1676037725
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1676037725
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 1676037725
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_84
timestamp 1676037725
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_148
timestamp 1676037725
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1676037725
transform 1 0 6256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_146
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1676037725
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1676037725
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_67
timestamp 1676037725
transform 1 0 7268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1676037725
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1676037725
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_102
timestamp 1676037725
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_126
timestamp 1676037725
transform 1 0 12696 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_154
timestamp 1676037725
transform 1 0 15272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1676037725
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1676037725
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1676037725
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1676037725
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_117
timestamp 1676037725
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_25
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_37
timestamp 1676037725
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1676037725
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_80
timestamp 1676037725
transform 1 0 8464 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_101
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_152
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1676037725
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1676037725
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1676037725
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1676037725
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1676037725
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_20
timestamp 1676037725
transform 1 0 2944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1676037725
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1676037725
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_78
timestamp 1676037725
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_118
timestamp 1676037725
transform 1 0 11960 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_130
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1676037725
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_17
timestamp 1676037725
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1676037725
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_36
timestamp 1676037725
transform 1 0 4416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1676037725
transform 1 0 5520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_118
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_64
timestamp 1676037725
transform 1 0 6992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_70
timestamp 1676037725
transform 1 0 7544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_92
timestamp 1676037725
transform 1 0 9568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_98
timestamp 1676037725
transform 1 0 10120 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1676037725
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1676037725
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_36
timestamp 1676037725
transform 1 0 4416 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_48
timestamp 1676037725
transform 1 0 5520 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_70
timestamp 1676037725
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_92
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 1676037725
transform 1 0 10120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1676037725
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1676037725
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_62
timestamp 1676037725
transform 1 0 6808 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_74
timestamp 1676037725
transform 1 0 7912 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_86
timestamp 1676037725
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1676037725
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1676037725
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_34
timestamp 1676037725
transform 1 0 4232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_46
timestamp 1676037725
transform 1 0 5336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_54
timestamp 1676037725
transform 1 0 6072 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1676037725
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1676037725
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_113
timestamp 1676037725
transform 1 0 11500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1676037725
transform 1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1676037725
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1676037725
transform -1 0 6072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1676037725
transform -1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1676037725
transform -1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1676037725
transform -1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1676037725
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1676037725
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1676037725
transform -1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1676037725
transform -1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1676037725
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1676037725
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1676037725
transform -1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1676037725
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1676037725
transform 1 0 2668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1676037725
transform -1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1676037725
transform -1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1676037725
transform -1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1676037725
transform -1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1676037725
transform 1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1676037725
transform -1 0 10488 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1676037725
transform 1 0 14996 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1676037725
transform -1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1676037725
transform -1 0 15180 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1676037725
transform -1 0 10212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1676037725
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1676037725
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125__1
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _127__10
timestamp 1676037725
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _129_
timestamp 1676037725
transform -1 0 3496 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _130_
timestamp 1676037725
transform -1 0 9292 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _131_
timestamp 1676037725
transform -1 0 4416 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _132_
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 1676037725
transform 1 0 14720 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _136_
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _138_
timestamp 1676037725
transform -1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12144 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _142_
timestamp 1676037725
transform 1 0 7912 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _144_
timestamp 1676037725
transform -1 0 7636 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  _146_
timestamp 1676037725
transform 1 0 4600 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4968 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8096 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_4  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1676037725
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _156_
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _159_
timestamp 1676037725
transform -1 0 4692 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3864 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1676037725
transform -1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1676037725
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _168_
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5152 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6348 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _171_
timestamp 1676037725
transform -1 0 7268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _172_
timestamp 1676037725
transform -1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _173__11
timestamp 1676037725
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__12
timestamp 1676037725
transform -1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175__13
timestamp 1676037725
transform -1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _176_
timestamp 1676037725
transform 1 0 9108 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _177_
timestamp 1676037725
transform -1 0 9568 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _178_
timestamp 1676037725
transform -1 0 3496 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _179_
timestamp 1676037725
transform -1 0 3404 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _180_
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _181_
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _182_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _183_
timestamp 1676037725
transform -1 0 3404 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _184__14
timestamp 1676037725
transform -1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185__15
timestamp 1676037725
transform -1 0 15824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186__16
timestamp 1676037725
transform -1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187__17
timestamp 1676037725
transform -1 0 15824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188__18
timestamp 1676037725
transform -1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189__19
timestamp 1676037725
transform -1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190__20
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191__21
timestamp 1676037725
transform -1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192__22
timestamp 1676037725
transform -1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193__2
timestamp 1676037725
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194__3
timestamp 1676037725
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195__4
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196__5
timestamp 1676037725
transform -1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197__23
timestamp 1676037725
transform -1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1676037725
transform -1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1676037725
transform 1 0 12420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1676037725
transform 1 0 15824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1676037725
transform 1 0 15364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1676037725
transform -1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1676037725
transform -1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1676037725
transform -1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1676037725
transform -1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207__6
timestamp 1676037725
transform -1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208__7
timestamp 1676037725
transform -1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _209_
timestamp 1676037725
transform -1 0 4508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1676037725
transform -1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1676037725
transform -1 0 2668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1676037725
transform -1 0 9752 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1676037725
transform -1 0 6072 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1676037725
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1676037725
transform -1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216__8
timestamp 1676037725
transform -1 0 4232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217__9
timestamp 1676037725
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1676037725
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1676037725
transform -1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1676037725
transform -1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _221_
timestamp 1676037725
transform -1 0 4416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1676037725
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1676037725
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1676037725
transform -1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _225_
timestamp 1676037725
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1676037725
transform 1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1676037725
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1676037725
transform -1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230__24
timestamp 1676037725
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1676037725
transform -1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _237_
timestamp 1676037725
transform 1 0 10580 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _238_
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _239_
timestamp 1676037725
transform -1 0 16376 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _240_
timestamp 1676037725
transform -1 0 16376 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _241_
timestamp 1676037725
transform 1 0 9844 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _242_
timestamp 1676037725
transform -1 0 16376 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _243_
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _244_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _245_
timestamp 1676037725
transform -1 0 12328 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_4  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5244 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _249_
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _250_
timestamp 1676037725
transform 1 0 2208 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _251_
timestamp 1676037725
transform -1 0 9568 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _252_
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _253_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _254_
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _255_
timestamp 1676037725
transform -1 0 4968 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _256_
timestamp 1676037725
transform 1 0 6900 0 1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfrtp_4  _257_
timestamp 1676037725
transform 1 0 1840 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _258_
timestamp 1676037725
transform 1 0 2208 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _259_
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _260_
timestamp 1676037725
transform 1 0 2392 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _261_
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _262_
timestamp 1676037725
transform 1 0 8188 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _263_
timestamp 1676037725
transform 1 0 9016 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _264_
timestamp 1676037725
transform 1 0 6716 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _265_
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _266_
timestamp 1676037725
transform -1 0 12696 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _267_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _268_
timestamp 1676037725
transform -1 0 16376 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _269_
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11132 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1676037725
transform 1 0 8924 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform -1 0 9016 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f__068_
timestamp 1676037725
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f__068_
timestamp 1676037725
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f__068_
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f__068_
timestamp 1676037725
transform 1 0 9384 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output3
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1676037725
transform 1 0 15824 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform -1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 12236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 15640 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 4434 17200 4490 18000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_out[10]
port 2 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 io_out[11]
port 3 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 io_out[1]
port 4 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 io_out[2]
port 5 nsew signal tristate
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 io_out[3]
port 6 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_out[4]
port 7 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 io_out[5]
port 8 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_out[6]
port 9 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_out[7]
port 10 nsew signal tristate
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 io_out[8]
port 11 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[9]
port 12 nsew signal tristate
flabel metal2 s 13450 17200 13506 18000 0 FreeSans 224 90 0 0 rst
port 13 nsew signal input
flabel metal4 s 2910 2128 3230 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 6843 2128 7163 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 10776 2128 11096 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 14709 2128 15029 15824 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 4876 2128 5196 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 8809 2128 9129 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 12742 2128 13062 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 16675 2128 16995 15824 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
