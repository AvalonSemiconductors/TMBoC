magic
tech sky130B
magscale 1 2
timestamp 1680605653
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 382 1776 68816 67584
<< metal2 >>
rect 3238 0 3294 800
rect 9586 0 9642 800
rect 15934 0 15990 800
rect 22282 0 22338 800
rect 28630 0 28686 800
rect 34978 0 35034 800
rect 41326 0 41382 800
rect 47674 0 47730 800
rect 54022 0 54078 800
rect 60370 0 60426 800
rect 66718 0 66774 800
<< obsm2 >>
rect 386 856 68244 67969
rect 386 734 3182 856
rect 3350 734 9530 856
rect 9698 734 15878 856
rect 16046 734 22226 856
rect 22394 734 28574 856
rect 28742 734 34922 856
rect 35090 734 41270 856
rect 41438 734 47618 856
rect 47786 734 53966 856
rect 54134 734 60314 856
rect 60482 734 66662 856
rect 66830 734 68244 856
<< metal3 >>
rect 0 67872 800 67992
rect 0 65424 800 65544
rect 0 62976 800 63096
rect 0 60528 800 60648
rect 0 58080 800 58200
rect 0 55632 800 55752
rect 0 53184 800 53304
rect 0 50736 800 50856
rect 0 48288 800 48408
rect 0 45840 800 45960
rect 0 43392 800 43512
rect 0 40944 800 41064
rect 0 38496 800 38616
rect 0 36048 800 36168
rect 0 33600 800 33720
rect 0 31152 800 31272
rect 0 28704 800 28824
rect 0 26256 800 26376
rect 0 23808 800 23928
rect 0 21360 800 21480
rect 0 18912 800 19032
rect 0 16464 800 16584
rect 0 14016 800 14136
rect 0 11568 800 11688
rect 0 9120 800 9240
rect 0 6672 800 6792
rect 0 4224 800 4344
rect 0 1776 800 1896
<< obsm3 >>
rect 880 67792 66227 67965
rect 381 65624 66227 67792
rect 880 65344 66227 65624
rect 381 63176 66227 65344
rect 880 62896 66227 63176
rect 381 60728 66227 62896
rect 880 60448 66227 60728
rect 381 58280 66227 60448
rect 880 58000 66227 58280
rect 381 55832 66227 58000
rect 880 55552 66227 55832
rect 381 53384 66227 55552
rect 880 53104 66227 53384
rect 381 50936 66227 53104
rect 880 50656 66227 50936
rect 381 48488 66227 50656
rect 880 48208 66227 48488
rect 381 46040 66227 48208
rect 880 45760 66227 46040
rect 381 43592 66227 45760
rect 880 43312 66227 43592
rect 381 41144 66227 43312
rect 880 40864 66227 41144
rect 381 38696 66227 40864
rect 880 38416 66227 38696
rect 381 36248 66227 38416
rect 880 35968 66227 36248
rect 381 33800 66227 35968
rect 880 33520 66227 33800
rect 381 31352 66227 33520
rect 880 31072 66227 31352
rect 381 28904 66227 31072
rect 880 28624 66227 28904
rect 381 26456 66227 28624
rect 880 26176 66227 26456
rect 381 24008 66227 26176
rect 880 23728 66227 24008
rect 381 21560 66227 23728
rect 880 21280 66227 21560
rect 381 19112 66227 21280
rect 880 18832 66227 19112
rect 381 16664 66227 18832
rect 880 16384 66227 16664
rect 381 14216 66227 16384
rect 880 13936 66227 14216
rect 381 11768 66227 13936
rect 880 11488 66227 11768
rect 381 9320 66227 11488
rect 880 9040 66227 9320
rect 381 6872 66227 9040
rect 880 6592 66227 6872
rect 381 4424 66227 6592
rect 880 4144 66227 4424
rect 381 1976 66227 4144
rect 880 1803 66227 1976
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 611 3163 4128 67013
rect 4608 3163 19488 67013
rect 19968 3163 34848 67013
rect 35328 3163 50208 67013
rect 50688 3163 56613 67013
<< labels >>
rlabel metal2 s 60370 0 60426 800 6 clk
port 1 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 io_in[8]
port 10 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_oeb
port 11 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_out[0]
port 12 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 io_out[10]
port 13 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 io_out[11]
port 14 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 io_out[12]
port 15 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 io_out[13]
port 16 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[14]
port 17 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_out[15]
port 18 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_out[16]
port 19 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_out[17]
port 20 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_out[18]
port 21 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_out[19]
port 22 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[1]
port 23 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 io_out[20]
port 24 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 io_out[21]
port 25 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_out[22]
port 26 nsew signal output
rlabel metal3 s 0 58080 800 58200 6 io_out[23]
port 27 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 io_out[24]
port 28 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 io_out[25]
port 29 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 io_out[26]
port 30 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_out[2]
port 31 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_out[3]
port 32 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[4]
port 33 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_out[5]
port 34 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 io_out[6]
port 35 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 io_out[7]
port 36 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[8]
port 37 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_out[9]
port 38 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 rst
port 39 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16772784
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS2650/runs/23_04_04_12_29/results/signoff/wrapped_as2650.magic.gds
string GDS_START 1393080
<< end >>

