// This is the unpowered netlist.
module wrapped_as2650 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [7:0] io_in;
 output [26:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.sense ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \lfsr[0] ;
 wire \lfsr[10] ;
 wire \lfsr[11] ;
 wire \lfsr[12] ;
 wire \lfsr[13] ;
 wire \lfsr[14] ;
 wire \lfsr[15] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \lfsr[8] ;
 wire \lfsr[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _3407_ (.A(io_out[21]),
    .Y(io_oeb));
 sky130_fd_sc_hd__buf_4 _3408_ (.A(net1),
    .X(_3028_));
 sky130_fd_sc_hd__buf_4 _3409_ (.A(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__clkbuf_4 _3410_ (.A(\as2650.addr_buff[0] ),
    .X(_3030_));
 sky130_fd_sc_hd__or4_1 _3411_ (.A(\as2650.cycle[7] ),
    .B(\as2650.cycle[6] ),
    .C(\as2650.cycle[5] ),
    .D(\as2650.cycle[4] ),
    .X(_3031_));
 sky130_fd_sc_hd__clkbuf_4 _3412_ (.A(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__clkbuf_2 _3413_ (.A(\as2650.cycle[3] ),
    .X(_3033_));
 sky130_fd_sc_hd__clkbuf_2 _3414_ (.A(\as2650.cycle[2] ),
    .X(_3034_));
 sky130_fd_sc_hd__inv_2 _3415_ (.A(\as2650.cycle[0] ),
    .Y(_3035_));
 sky130_fd_sc_hd__or4_2 _3416_ (.A(_3033_),
    .B(_3034_),
    .C(\as2650.cycle[1] ),
    .D(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__nor2_2 _3417_ (.A(_3032_),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__buf_2 _3418_ (.A(\as2650.ins_reg[4] ),
    .X(_3038_));
 sky130_fd_sc_hd__buf_4 _3419_ (.A(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__buf_4 _3420_ (.A(\as2650.cycle[1] ),
    .X(_3040_));
 sky130_fd_sc_hd__or3b_1 _3421_ (.A(_3034_),
    .B(_3032_),
    .C_N(_3033_),
    .X(_3041_));
 sky130_fd_sc_hd__or2_1 _3422_ (.A(_3040_),
    .B(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__nor2_1 _3423_ (.A(_3039_),
    .B(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__or3_1 _3424_ (.A(_3033_),
    .B(_3034_),
    .C(_3032_),
    .X(_3044_));
 sky130_fd_sc_hd__buf_4 _3425_ (.A(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__buf_4 _3426_ (.A(\as2650.cycle[0] ),
    .X(_3046_));
 sky130_fd_sc_hd__or2_4 _3427_ (.A(\as2650.cycle[1] ),
    .B(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__or2_1 _3428_ (.A(_3045_),
    .B(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__clkinv_4 _3429_ (.A(\as2650.ins_reg[4] ),
    .Y(_3049_));
 sky130_fd_sc_hd__or4b_4 _3430_ (.A(\as2650.cycle[3] ),
    .B(_3035_),
    .C(\as2650.cycle[2] ),
    .D_N(\as2650.cycle[1] ),
    .X(_3050_));
 sky130_fd_sc_hd__nor2_4 _3431_ (.A(_3032_),
    .B(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__nand2_1 _3432_ (.A(_3049_),
    .B(_3051_),
    .Y(_3052_));
 sky130_fd_sc_hd__nand2_1 _3433_ (.A(_3048_),
    .B(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__or3_1 _3434_ (.A(_3037_),
    .B(_3043_),
    .C(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__or2_1 _3435_ (.A(\as2650.halted ),
    .B(net9),
    .X(_3055_));
 sky130_fd_sc_hd__buf_4 _3436_ (.A(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__or3b_2 _3437_ (.A(_3047_),
    .B(_3033_),
    .C_N(_3034_),
    .X(_3057_));
 sky130_fd_sc_hd__clkinv_2 _3438_ (.A(\as2650.cycle[7] ),
    .Y(_3058_));
 sky130_fd_sc_hd__or3_1 _3439_ (.A(_3033_),
    .B(_3034_),
    .C(_3047_),
    .X(_3059_));
 sky130_fd_sc_hd__or4_4 _3440_ (.A(_3058_),
    .B(\as2650.cycle[5] ),
    .C(\as2650.cycle[4] ),
    .D(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__nor2_2 _3441_ (.A(\as2650.cycle[6] ),
    .B(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__nor2_4 _3442_ (.A(_3045_),
    .B(_3047_),
    .Y(_3062_));
 sky130_fd_sc_hd__nor2_1 _3443_ (.A(_3039_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__nand2_1 _3444_ (.A(_3061_),
    .B(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__clkbuf_4 _3445_ (.A(\as2650.ins_reg[2] ),
    .X(_3065_));
 sky130_fd_sc_hd__nand2_2 _3446_ (.A(\as2650.ins_reg[3] ),
    .B(_3038_),
    .Y(_3066_));
 sky130_fd_sc_hd__buf_4 _3447_ (.A(\as2650.ins_reg[6] ),
    .X(_3067_));
 sky130_fd_sc_hd__buf_4 _3448_ (.A(\as2650.ins_reg[7] ),
    .X(_3068_));
 sky130_fd_sc_hd__nand2b_4 _3449_ (.A_N(_3067_),
    .B(_3068_),
    .Y(_3069_));
 sky130_fd_sc_hd__clkbuf_4 _3450_ (.A(\as2650.ins_reg[0] ),
    .X(_3070_));
 sky130_fd_sc_hd__clkbuf_4 _3451_ (.A(\as2650.ins_reg[1] ),
    .X(_3071_));
 sky130_fd_sc_hd__nand2_2 _3452_ (.A(_3070_),
    .B(_3071_),
    .Y(_3072_));
 sky130_fd_sc_hd__clkbuf_4 _3453_ (.A(_3072_),
    .X(_3073_));
 sky130_fd_sc_hd__or3_2 _3454_ (.A(_3066_),
    .B(_3069_),
    .C(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__or2_1 _3455_ (.A(_3065_),
    .B(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__buf_4 _3456_ (.A(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__nand2_2 _3457_ (.A(\as2650.cycle[1] ),
    .B(_3035_),
    .Y(_3077_));
 sky130_fd_sc_hd__or2_1 _3458_ (.A(_3045_),
    .B(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__buf_4 _3459_ (.A(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__buf_4 _3460_ (.A(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__buf_4 _3461_ (.A(_3065_),
    .X(_3081_));
 sky130_fd_sc_hd__or2_1 _3462_ (.A(_3032_),
    .B(_3050_),
    .X(_3082_));
 sky130_fd_sc_hd__buf_2 _3463_ (.A(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__or2_1 _3464_ (.A(_3081_),
    .B(_3083_),
    .X(_3084_));
 sky130_fd_sc_hd__clkbuf_4 _3465_ (.A(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__a31o_1 _3466_ (.A1(_3076_),
    .A2(_3080_),
    .A3(_3085_),
    .B1(_3066_),
    .X(_3086_));
 sky130_fd_sc_hd__nand3_1 _3467_ (.A(_3057_),
    .B(_3064_),
    .C(_3086_),
    .Y(_3087_));
 sky130_fd_sc_hd__or3b_2 _3468_ (.A(\as2650.cycle[5] ),
    .B(\as2650.cycle[4] ),
    .C_N(\as2650.cycle[6] ),
    .X(_3088_));
 sky130_fd_sc_hd__nor2_1 _3469_ (.A(_3036_),
    .B(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__nand2_4 _3470_ (.A(\as2650.cycle[7] ),
    .B(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__clkbuf_4 _3471_ (.A(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__nor2_1 _3472_ (.A(_3088_),
    .B(_3059_),
    .Y(_3092_));
 sky130_fd_sc_hd__nand2_1 _3473_ (.A(_3058_),
    .B(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_3090_),
    .B(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__nor2_1 _3475_ (.A(_3040_),
    .B(_3041_),
    .Y(_3095_));
 sky130_fd_sc_hd__or2_1 _3476_ (.A(_3032_),
    .B(_3057_),
    .X(_3096_));
 sky130_fd_sc_hd__buf_4 _3477_ (.A(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__nand2_2 _3478_ (.A(_3083_),
    .B(_3097_),
    .Y(_3098_));
 sky130_fd_sc_hd__or3b_1 _3479_ (.A(_3095_),
    .B(_3098_),
    .C_N(_3060_),
    .X(_3099_));
 sky130_fd_sc_hd__or2_1 _3480_ (.A(_3094_),
    .B(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_4 _3481_ (.A(_3039_),
    .X(_3101_));
 sky130_fd_sc_hd__nor2_4 _3482_ (.A(_3045_),
    .B(_3077_),
    .Y(_3102_));
 sky130_fd_sc_hd__nor2_4 _3483_ (.A(_3101_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__inv_2 _3484_ (.A(\as2650.ins_reg[3] ),
    .Y(_3104_));
 sky130_fd_sc_hd__nor2_1 _3485_ (.A(_3104_),
    .B(_3049_),
    .Y(_3105_));
 sky130_fd_sc_hd__and2b_1 _3486_ (.A_N(_3067_),
    .B(_3068_),
    .X(_3106_));
 sky130_fd_sc_hd__buf_4 _3487_ (.A(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__and2_1 _3488_ (.A(_3070_),
    .B(\as2650.ins_reg[1] ),
    .X(_3108_));
 sky130_fd_sc_hd__clkbuf_4 _3489_ (.A(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__and3_2 _3490_ (.A(_3105_),
    .B(_3107_),
    .C(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__and2_1 _3491_ (.A(_3065_),
    .B(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__nor2_1 _3492_ (.A(_3047_),
    .B(_3041_),
    .Y(_3112_));
 sky130_fd_sc_hd__nand2_1 _3493_ (.A(_3083_),
    .B(_3111_),
    .Y(_3113_));
 sky130_fd_sc_hd__or3b_4 _3494_ (.A(_3032_),
    .B(_3033_),
    .C_N(_3034_),
    .X(_3114_));
 sky130_fd_sc_hd__nor2_1 _3495_ (.A(_3040_),
    .B(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__o32a_1 _3496_ (.A1(_3111_),
    .A2(_3112_),
    .A3(_3098_),
    .B1(_3113_),
    .B2(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__nor2_2 _3497_ (.A(_3081_),
    .B(_3074_),
    .Y(_3117_));
 sky130_fd_sc_hd__nor3_2 _3498_ (.A(_3033_),
    .B(_3034_),
    .C(_3032_),
    .Y(_3118_));
 sky130_fd_sc_hd__nand2_4 _3499_ (.A(_3040_),
    .B(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__nor2_4 _3500_ (.A(_3046_),
    .B(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__buf_4 _3501_ (.A(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__or3_1 _3502_ (.A(_3116_),
    .B(_3117_),
    .C(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__clkbuf_4 _3503_ (.A(_3105_),
    .X(_3123_));
 sky130_fd_sc_hd__a32o_1 _3504_ (.A1(_3091_),
    .A2(_3100_),
    .A3(_3103_),
    .B1(_3122_),
    .B2(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__or4b_1 _3505_ (.A(_3054_),
    .B(_3056_),
    .C(_3087_),
    .D_N(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__buf_2 _3506_ (.A(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(_3029_),
    .A1(_3030_),
    .S(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(_3127_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _3509_ (.A(net2),
    .X(_3128_));
 sky130_fd_sc_hd__buf_4 _3510_ (.A(_3128_),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(_3129_),
    .A1(\as2650.addr_buff[1] ),
    .S(_3126_),
    .X(_3130_));
 sky130_fd_sc_hd__clkbuf_1 _3512_ (.A(_3130_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_4 _3513_ (.A(net3),
    .X(_3131_));
 sky130_fd_sc_hd__buf_4 _3514_ (.A(_3131_),
    .X(_3132_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(_3132_),
    .A1(\as2650.addr_buff[2] ),
    .S(_3126_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_1 _3516_ (.A(_3133_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _3517_ (.A(net4),
    .X(_3134_));
 sky130_fd_sc_hd__buf_4 _3518_ (.A(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(_3135_),
    .A1(\as2650.addr_buff[3] ),
    .S(_3126_),
    .X(_3136_));
 sky130_fd_sc_hd__clkbuf_1 _3520_ (.A(_3136_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_4 _3521_ (.A(net5),
    .X(_3137_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(_3137_),
    .A1(\as2650.addr_buff[4] ),
    .S(_3126_),
    .X(_3138_));
 sky130_fd_sc_hd__clkbuf_1 _3523_ (.A(_3138_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _3524_ (.A(net6),
    .X(_3139_));
 sky130_fd_sc_hd__buf_6 _3525_ (.A(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(_3140_),
    .A1(\as2650.addr_buff[5] ),
    .S(_3126_),
    .X(_3141_));
 sky130_fd_sc_hd__clkbuf_1 _3527_ (.A(_3141_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_4 _3528_ (.A(net7),
    .X(_3142_));
 sky130_fd_sc_hd__buf_4 _3529_ (.A(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__buf_6 _3530_ (.A(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(_3144_),
    .A1(\as2650.addr_buff[6] ),
    .S(_3126_),
    .X(_3145_));
 sky130_fd_sc_hd__clkbuf_1 _3532_ (.A(_3145_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _3533_ (.A(net8),
    .X(_3146_));
 sky130_fd_sc_hd__buf_6 _3534_ (.A(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_4 _3535_ (.A(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__buf_4 _3536_ (.A(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__buf_6 _3537_ (.A(_3149_),
    .X(_3150_));
 sky130_fd_sc_hd__buf_4 _3538_ (.A(\as2650.addr_buff[7] ),
    .X(_3151_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(_3150_),
    .A1(_3151_),
    .S(_3126_),
    .X(_3152_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_3152_),
    .X(_0007_));
 sky130_fd_sc_hd__clkinv_2 _3541_ (.A(net9),
    .Y(_3153_));
 sky130_fd_sc_hd__clkbuf_4 _3542_ (.A(_3153_),
    .X(_3154_));
 sky130_fd_sc_hd__clkbuf_4 _3543_ (.A(_3035_),
    .X(_3155_));
 sky130_fd_sc_hd__and2_1 _3544_ (.A(\as2650.cycle[1] ),
    .B(_3118_),
    .X(_3156_));
 sky130_fd_sc_hd__nand2_1 _3545_ (.A(_3155_),
    .B(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__clkbuf_4 _3546_ (.A(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__buf_4 _3548_ (.A(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__clkbuf_4 _3549_ (.A(\as2650.psl[4] ),
    .X(_3161_));
 sky130_fd_sc_hd__buf_4 _3550_ (.A(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__buf_4 _3551_ (.A(_3162_),
    .X(_3163_));
 sky130_fd_sc_hd__or2_1 _3552_ (.A(_3163_),
    .B(_3056_),
    .X(_3164_));
 sky130_fd_sc_hd__buf_4 _3553_ (.A(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__nor2_1 _3554_ (.A(_3070_),
    .B(_3071_),
    .Y(_3166_));
 sky130_fd_sc_hd__buf_4 _3555_ (.A(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__nor2_4 _3556_ (.A(\as2650.ins_reg[2] ),
    .B(\as2650.ins_reg[3] ),
    .Y(_3168_));
 sky130_fd_sc_hd__nand2_2 _3557_ (.A(_3167_),
    .B(_3168_),
    .Y(_3169_));
 sky130_fd_sc_hd__nor2_4 _3558_ (.A(_3067_),
    .B(_3068_),
    .Y(_3170_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(_3038_),
    .B(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__or2_1 _3560_ (.A(\as2650.ins_reg[5] ),
    .B(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__clkbuf_4 _3561_ (.A(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__or2_2 _3562_ (.A(_3169_),
    .B(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__or2_2 _3563_ (.A(\as2650.ins_reg[2] ),
    .B(\as2650.ins_reg[3] ),
    .X(_3175_));
 sky130_fd_sc_hd__buf_4 _3564_ (.A(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__or3_2 _3565_ (.A(_3049_),
    .B(\as2650.ins_reg[5] ),
    .C(_3069_),
    .X(_3177_));
 sky130_fd_sc_hd__clkbuf_4 _3566_ (.A(_3070_),
    .X(_3178_));
 sky130_fd_sc_hd__inv_2 _3567_ (.A(_3071_),
    .Y(_3179_));
 sky130_fd_sc_hd__nand2_2 _3568_ (.A(_3178_),
    .B(_3179_),
    .Y(_3180_));
 sky130_fd_sc_hd__or3_4 _3569_ (.A(_3176_),
    .B(_3177_),
    .C(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__and2_1 _3570_ (.A(_3174_),
    .B(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__or3_2 _3571_ (.A(_3160_),
    .B(_3165_),
    .C(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__inv_2 _3572_ (.A(_3163_),
    .Y(_3184_));
 sky130_fd_sc_hd__or2_2 _3573_ (.A(_3070_),
    .B(\as2650.ins_reg[1] ),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_4 _3574_ (.A(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__nand2_1 _3575_ (.A(_3184_),
    .B(_3186_),
    .Y(_3187_));
 sky130_fd_sc_hd__or2_2 _3576_ (.A(_3056_),
    .B(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__inv_2 _3577_ (.A(\as2650.ins_reg[5] ),
    .Y(_3189_));
 sky130_fd_sc_hd__and3_1 _3578_ (.A(\as2650.ins_reg[4] ),
    .B(_3067_),
    .C(_3068_),
    .X(_3190_));
 sky130_fd_sc_hd__nand2_1 _3579_ (.A(_3189_),
    .B(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__or2_1 _3580_ (.A(_3065_),
    .B(_3191_),
    .X(_3192_));
 sky130_fd_sc_hd__nand2_2 _3581_ (.A(_3104_),
    .B(_3120_),
    .Y(_3193_));
 sky130_fd_sc_hd__or3_1 _3582_ (.A(_3188_),
    .B(_3192_),
    .C(_3193_),
    .X(_3194_));
 sky130_fd_sc_hd__buf_2 _3583_ (.A(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__nand2_2 _3584_ (.A(\as2650.ins_reg[4] ),
    .B(\as2650.ins_reg[5] ),
    .Y(_3196_));
 sky130_fd_sc_hd__or2_4 _3585_ (.A(\as2650.ins_reg[2] ),
    .B(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__nor2_2 _3586_ (.A(_3068_),
    .B(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__nand2_1 _3587_ (.A(_3104_),
    .B(_3198_),
    .Y(_3199_));
 sky130_fd_sc_hd__or2_2 _3588_ (.A(_3083_),
    .B(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__or2_1 _3589_ (.A(_3188_),
    .B(_3200_),
    .X(_3201_));
 sky130_fd_sc_hd__buf_4 _3590_ (.A(_3168_),
    .X(_3202_));
 sky130_fd_sc_hd__nand2_2 _3591_ (.A(\as2650.ins_reg[6] ),
    .B(\as2650.ins_reg[7] ),
    .Y(_3203_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(\as2650.ins_reg[5] ),
    .B(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__buf_4 _3593_ (.A(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__nor2_1 _3594_ (.A(_3039_),
    .B(_3205_),
    .Y(_3206_));
 sky130_fd_sc_hd__nand2_1 _3595_ (.A(_3202_),
    .B(_3206_),
    .Y(_3207_));
 sky130_fd_sc_hd__or4_2 _3596_ (.A(_3158_),
    .B(_3167_),
    .C(_3207_),
    .D(_3165_),
    .X(_3208_));
 sky130_fd_sc_hd__or2_1 _3597_ (.A(_3038_),
    .B(_3055_),
    .X(_3209_));
 sky130_fd_sc_hd__nor2_2 _3598_ (.A(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_3210_));
 sky130_fd_sc_hd__or2_1 _3599_ (.A(\as2650.addr_buff[7] ),
    .B(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__buf_2 _3600_ (.A(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__or4_2 _3601_ (.A(_3090_),
    .B(_3187_),
    .C(_3209_),
    .D(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__nand2_2 _3602_ (.A(_3058_),
    .B(_3089_),
    .Y(_3214_));
 sky130_fd_sc_hd__nor2_1 _3603_ (.A(_3038_),
    .B(_3055_),
    .Y(_3215_));
 sky130_fd_sc_hd__or2_2 _3604_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .X(_3216_));
 sky130_fd_sc_hd__nand2_1 _3605_ (.A(_3215_),
    .B(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__or3_1 _3606_ (.A(_3187_),
    .B(_3214_),
    .C(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__and4_1 _3607_ (.A(_3201_),
    .B(_3208_),
    .C(_3213_),
    .D(_3218_),
    .X(_3219_));
 sky130_fd_sc_hd__nor2b_4 _3608_ (.A(_3068_),
    .B_N(\as2650.ins_reg[6] ),
    .Y(_3220_));
 sky130_fd_sc_hd__nand2_4 _3609_ (.A(_3189_),
    .B(_3220_),
    .Y(_3221_));
 sky130_fd_sc_hd__or3_1 _3610_ (.A(\as2650.ins_reg[2] ),
    .B(_3049_),
    .C(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__or3_2 _3611_ (.A(\as2650.ins_reg[3] ),
    .B(_3157_),
    .C(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__or2_1 _3612_ (.A(_3188_),
    .B(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__clkbuf_2 _3613_ (.A(_3224_),
    .X(_3225_));
 sky130_fd_sc_hd__nand2_2 _3614_ (.A(_3039_),
    .B(_3067_),
    .Y(_3226_));
 sky130_fd_sc_hd__buf_4 _3615_ (.A(\as2650.ins_reg[3] ),
    .X(_3227_));
 sky130_fd_sc_hd__nand2_4 _3616_ (.A(_3227_),
    .B(_3120_),
    .Y(_3228_));
 sky130_fd_sc_hd__nor2_2 _3617_ (.A(_3189_),
    .B(_3203_),
    .Y(_3229_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_3186_),
    .B(_3176_),
    .Y(_3230_));
 sky130_fd_sc_hd__or2_1 _3619_ (.A(_3229_),
    .B(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__or4_1 _3620_ (.A(_3101_),
    .B(_3097_),
    .C(_3216_),
    .D(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__o32a_1 _3621_ (.A1(_3188_),
    .A2(_3226_),
    .A3(_3228_),
    .B1(_3232_),
    .B2(_3165_),
    .X(_3233_));
 sky130_fd_sc_hd__and4_4 _3622_ (.A(_3195_),
    .B(_3219_),
    .C(_3225_),
    .D(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__or2_2 _3623_ (.A(_3071_),
    .B(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__nand3_4 _3624_ (.A(_3154_),
    .B(_3183_),
    .C(_3235_),
    .Y(_3236_));
 sky130_fd_sc_hd__clkinv_2 _3625_ (.A(_3235_),
    .Y(_3237_));
 sky130_fd_sc_hd__or3_4 _3626_ (.A(_3187_),
    .B(_3214_),
    .C(_3217_),
    .X(_3238_));
 sky130_fd_sc_hd__mux2_4 _3627_ (.A0(\as2650.r123[2][0] ),
    .A1(\as2650.r123_2[2][0] ),
    .S(_3161_),
    .X(_3239_));
 sky130_fd_sc_hd__and2_2 _3628_ (.A(_3109_),
    .B(_3239_),
    .X(_3240_));
 sky130_fd_sc_hd__mux4_2 _3629_ (.A0(\as2650.r123[1][0] ),
    .A1(\as2650.r123[0][0] ),
    .A2(\as2650.r123_2[1][0] ),
    .A3(\as2650.r123_2[0][0] ),
    .S0(_3070_),
    .S1(_3161_),
    .X(_3241_));
 sky130_fd_sc_hd__nor3b_2 _3630_ (.A(_3070_),
    .B(_3071_),
    .C_N(\as2650.r0[0] ),
    .Y(_3242_));
 sky130_fd_sc_hd__a31o_2 _3631_ (.A1(_3073_),
    .A2(_3185_),
    .A3(_3241_),
    .B1(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__nor2_8 _3632_ (.A(_3240_),
    .B(_3243_),
    .Y(_3244_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(\as2650.idx_ctrl[1] ),
    .Y(_3245_));
 sky130_fd_sc_hd__nand2_2 _3634_ (.A(_3245_),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_3246_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(\as2650.idx_ctrl[0] ),
    .Y(_3247_));
 sky130_fd_sc_hd__nand2_4 _3636_ (.A(\as2650.idx_ctrl[1] ),
    .B(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__nand2_4 _3637_ (.A(_3246_),
    .B(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__xnor2_4 _3638_ (.A(_3244_),
    .B(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__or2_2 _3639_ (.A(_3036_),
    .B(_3088_),
    .X(_3251_));
 sky130_fd_sc_hd__nor2_4 _3640_ (.A(_3058_),
    .B(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__nor2_1 _3641_ (.A(_3163_),
    .B(_3167_),
    .Y(_3253_));
 sky130_fd_sc_hd__nor2_4 _3642_ (.A(_3151_),
    .B(_3210_),
    .Y(_3254_));
 sky130_fd_sc_hd__and4_1 _3643_ (.A(_3252_),
    .B(_3253_),
    .C(_3215_),
    .D(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__buf_2 _3644_ (.A(_3255_),
    .X(_3256_));
 sky130_fd_sc_hd__nand2b_4 _3645_ (.A_N(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_3257_));
 sky130_fd_sc_hd__nand2b_4 _3646_ (.A_N(\as2650.addr_buff[5] ),
    .B(\as2650.addr_buff[6] ),
    .Y(_3258_));
 sky130_fd_sc_hd__nand2_4 _3647_ (.A(_3257_),
    .B(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__xnor2_4 _3648_ (.A(_3244_),
    .B(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__buf_2 _3649_ (.A(\as2650.r0[0] ),
    .X(_3261_));
 sky130_fd_sc_hd__buf_4 _3650_ (.A(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__or2_1 _3651_ (.A(_3176_),
    .B(_3191_),
    .X(_3263_));
 sky130_fd_sc_hd__nor3_1 _3652_ (.A(_3159_),
    .B(_3188_),
    .C(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(\as2650.r123[2][7] ),
    .A1(\as2650.r123_2[2][7] ),
    .S(_3163_),
    .X(_3265_));
 sky130_fd_sc_hd__a22o_1 _3654_ (.A1(\as2650.r0[7] ),
    .A2(_3167_),
    .B1(_3265_),
    .B2(_3109_),
    .X(_3266_));
 sky130_fd_sc_hd__mux4_1 _3655_ (.A0(\as2650.r123[1][7] ),
    .A1(\as2650.r123[0][7] ),
    .A2(\as2650.r123_2[1][7] ),
    .A3(\as2650.r123_2[0][7] ),
    .S0(_3178_),
    .S1(_3163_),
    .X(_3267_));
 sky130_fd_sc_hd__and3_1 _3656_ (.A(_3073_),
    .B(_3186_),
    .C(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__or2_1 _3657_ (.A(_3266_),
    .B(_3268_),
    .X(_3269_));
 sky130_fd_sc_hd__buf_2 _3658_ (.A(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_4 _3659_ (.A(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__or2b_1 _3660_ (.A(\as2650.carry ),
    .B_N(\as2650.psl[3] ),
    .X(_3272_));
 sky130_fd_sc_hd__o21a_1 _3661_ (.A1(\as2650.psl[3] ),
    .A2(_3271_),
    .B1(_3272_),
    .X(_3273_));
 sky130_fd_sc_hd__mux4_1 _3662_ (.A0(\as2650.r123[1][1] ),
    .A1(\as2650.r123[0][1] ),
    .A2(\as2650.r123_2[1][1] ),
    .A3(\as2650.r123_2[0][1] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(\as2650.psl[4] ),
    .X(_3274_));
 sky130_fd_sc_hd__and3_1 _3663_ (.A(_3072_),
    .B(_3185_),
    .C(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__mux2_4 _3664_ (.A0(\as2650.r123[2][1] ),
    .A1(\as2650.r123_2[2][1] ),
    .S(\as2650.psl[4] ),
    .X(_3276_));
 sky130_fd_sc_hd__a22o_1 _3665_ (.A1(\as2650.r0[1] ),
    .A2(_3166_),
    .B1(_3276_),
    .B2(_3108_),
    .X(_3277_));
 sky130_fd_sc_hd__or2_4 _3666_ (.A(_3275_),
    .B(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__buf_4 _3667_ (.A(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__buf_4 _3668_ (.A(_3279_),
    .X(_3280_));
 sky130_fd_sc_hd__nor2_1 _3669_ (.A(_3188_),
    .B(_3200_),
    .Y(_3281_));
 sky130_fd_sc_hd__buf_2 _3670_ (.A(_3281_),
    .X(_3282_));
 sky130_fd_sc_hd__nor2_2 _3671_ (.A(_3188_),
    .B(_3223_),
    .Y(_3283_));
 sky130_fd_sc_hd__nand2_1 _3672_ (.A(_3109_),
    .B(_3239_),
    .Y(_3284_));
 sky130_fd_sc_hd__a31oi_4 _3673_ (.A1(_3072_),
    .A2(_3185_),
    .A3(_3241_),
    .B1(_3242_),
    .Y(_3285_));
 sky130_fd_sc_hd__nand2_4 _3674_ (.A(_3284_),
    .B(_3285_),
    .Y(_3286_));
 sky130_fd_sc_hd__buf_4 _3675_ (.A(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__xnor2_2 _3676_ (.A(_3190_),
    .B(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__nor2_1 _3677_ (.A(_3282_),
    .B(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__a211o_1 _3678_ (.A1(_3028_),
    .A2(_3282_),
    .B1(_3283_),
    .C1(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__o211a_1 _3679_ (.A1(_3225_),
    .A2(_3280_),
    .B1(_3290_),
    .C1(_3195_),
    .X(_3291_));
 sky130_fd_sc_hd__buf_4 _3680_ (.A(_3176_),
    .X(_3292_));
 sky130_fd_sc_hd__or2_1 _3681_ (.A(_3038_),
    .B(_3205_),
    .X(_3293_));
 sky130_fd_sc_hd__nor2_1 _3682_ (.A(_3292_),
    .B(_3293_),
    .Y(_3294_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(_3079_),
    .B(_3165_),
    .Y(_3295_));
 sky130_fd_sc_hd__and3_2 _3684_ (.A(_3186_),
    .B(_3294_),
    .C(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__a211o_1 _3685_ (.A1(_3264_),
    .A2(_3273_),
    .B1(_3291_),
    .C1(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__o211a_1 _3686_ (.A1(_3262_),
    .A2(_3208_),
    .B1(_3213_),
    .C1(_3297_),
    .X(_3298_));
 sky130_fd_sc_hd__nor2_1 _3687_ (.A(\as2650.cycle[7] ),
    .B(_3251_),
    .Y(_3299_));
 sky130_fd_sc_hd__nor2_2 _3688_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_3300_));
 sky130_fd_sc_hd__nor2_1 _3689_ (.A(_3209_),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__and3_2 _3690_ (.A(_3253_),
    .B(_3299_),
    .C(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__a211o_1 _3691_ (.A1(_3256_),
    .A2(_3260_),
    .B1(_3298_),
    .C1(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__o21a_1 _3692_ (.A1(_3238_),
    .A2(_3250_),
    .B1(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__or2_1 _3693_ (.A(\as2650.holding_reg[0] ),
    .B(_3168_),
    .X(_3305_));
 sky130_fd_sc_hd__o31a_2 _3694_ (.A1(_3175_),
    .A2(_3240_),
    .A3(_3243_),
    .B1(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__nor2_1 _3695_ (.A(\as2650.holding_reg[0] ),
    .B(_3175_),
    .Y(_3307_));
 sky130_fd_sc_hd__a31o_2 _3696_ (.A1(_3175_),
    .A2(_3284_),
    .A3(_3285_),
    .B1(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__xor2_4 _3697_ (.A(_3306_),
    .B(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__inv_2 _3698_ (.A(_3309_),
    .Y(_3310_));
 sky130_fd_sc_hd__nand2_1 _3699_ (.A(\as2650.psl[3] ),
    .B(\as2650.carry ),
    .Y(_3311_));
 sky130_fd_sc_hd__nor2_2 _3700_ (.A(\as2650.ins_reg[5] ),
    .B(_3069_),
    .Y(_3312_));
 sky130_fd_sc_hd__o21ai_1 _3701_ (.A1(_3311_),
    .A2(_3309_),
    .B1(_3312_),
    .Y(_3313_));
 sky130_fd_sc_hd__a21oi_1 _3702_ (.A1(_3311_),
    .A2(_3309_),
    .B1(_3313_),
    .Y(_3314_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_3272_),
    .B(_3309_),
    .Y(_3315_));
 sky130_fd_sc_hd__o2111a_1 _3704_ (.A1(_3272_),
    .A2(_3309_),
    .B1(_3315_),
    .C1(_3107_),
    .D1(\as2650.ins_reg[5] ),
    .X(_3316_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(_3308_),
    .Y(_3317_));
 sky130_fd_sc_hd__nand2b_2 _3706_ (.A_N(\as2650.ins_reg[7] ),
    .B(\as2650.ins_reg[6] ),
    .Y(_3318_));
 sky130_fd_sc_hd__nor2_4 _3707_ (.A(\as2650.ins_reg[5] ),
    .B(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__a221o_1 _3708_ (.A1(_3069_),
    .A2(_3306_),
    .B1(_3317_),
    .B2(_3220_),
    .C1(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__and2_1 _3709_ (.A(\as2650.holding_reg[0] ),
    .B(_3287_),
    .X(_3321_));
 sky130_fd_sc_hd__o32a_1 _3710_ (.A1(_3314_),
    .A2(_3316_),
    .A3(_3320_),
    .B1(_3321_),
    .B2(_3221_),
    .X(_3322_));
 sky130_fd_sc_hd__buf_4 _3711_ (.A(\as2650.ins_reg[5] ),
    .X(_3323_));
 sky130_fd_sc_hd__nand2_4 _3712_ (.A(_3323_),
    .B(_3170_),
    .Y(_3324_));
 sky130_fd_sc_hd__mux2_2 _3713_ (.A0(_3310_),
    .A1(_3322_),
    .S(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__or2_2 _3714_ (.A(_3114_),
    .B(_3047_),
    .X(_3326_));
 sky130_fd_sc_hd__or4_2 _3715_ (.A(_3038_),
    .B(_3326_),
    .C(_3216_),
    .D(_3231_),
    .X(_3327_));
 sky130_fd_sc_hd__nor2_2 _3716_ (.A(_3165_),
    .B(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__mux2_2 _3717_ (.A0(_3304_),
    .A1(_3325_),
    .S(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__buf_4 _3718_ (.A(_3160_),
    .X(_3330_));
 sky130_fd_sc_hd__buf_2 _3719_ (.A(_3174_),
    .X(_3331_));
 sky130_fd_sc_hd__or3_2 _3720_ (.A(_3330_),
    .B(_3165_),
    .C(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__nor2_2 _3721_ (.A(\as2650.psu[0] ),
    .B(\as2650.psu[1] ),
    .Y(_3333_));
 sky130_fd_sc_hd__nor2_8 _3722_ (.A(\as2650.psu[2] ),
    .B(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__clkbuf_4 _3723_ (.A(_3333_),
    .X(_3335_));
 sky130_fd_sc_hd__nand2_4 _3724_ (.A(\as2650.psu[2] ),
    .B(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__nor2b_4 _3725_ (.A(_3334_),
    .B_N(_3336_),
    .Y(_3337_));
 sky130_fd_sc_hd__buf_4 _3726_ (.A(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__buf_6 _3727_ (.A(\as2650.psu[0] ),
    .X(_3339_));
 sky130_fd_sc_hd__or2_1 _3728_ (.A(_3339_),
    .B(\as2650.psu[1] ),
    .X(_3340_));
 sky130_fd_sc_hd__clkbuf_4 _3729_ (.A(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__clkbuf_4 _3730_ (.A(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__buf_4 _3731_ (.A(\as2650.psu[1] ),
    .X(_3343_));
 sky130_fd_sc_hd__nand2_2 _3732_ (.A(_3339_),
    .B(_3343_),
    .Y(_3344_));
 sky130_fd_sc_hd__clkbuf_4 _3733_ (.A(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__clkbuf_4 _3734_ (.A(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__o22a_1 _3735_ (.A1(\as2650.stack[7][8] ),
    .A2(_3342_),
    .B1(_3346_),
    .B2(\as2650.stack[6][8] ),
    .X(_3347_));
 sky130_fd_sc_hd__inv_2 _3736_ (.A(\as2650.psu[0] ),
    .Y(_3348_));
 sky130_fd_sc_hd__or2_1 _3737_ (.A(_3348_),
    .B(\as2650.psu[1] ),
    .X(_3349_));
 sky130_fd_sc_hd__clkbuf_4 _3738_ (.A(_3349_),
    .X(_3350_));
 sky130_fd_sc_hd__buf_4 _3739_ (.A(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_4 _3740_ (.A(_3351_),
    .X(_3352_));
 sky130_fd_sc_hd__nand2_1 _3741_ (.A(_3348_),
    .B(\as2650.psu[1] ),
    .Y(_3353_));
 sky130_fd_sc_hd__clkbuf_4 _3742_ (.A(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_4 _3743_ (.A(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__o22a_1 _3744_ (.A1(\as2650.stack[4][8] ),
    .A2(_3352_),
    .B1(_3355_),
    .B2(\as2650.stack[5][8] ),
    .X(_3356_));
 sky130_fd_sc_hd__and3_1 _3745_ (.A(\as2650.psu[2] ),
    .B(\as2650.stack[3][8] ),
    .C(_3335_),
    .X(_3357_));
 sky130_fd_sc_hd__o22a_1 _3746_ (.A1(\as2650.stack[0][8] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[1][8] ),
    .X(_3358_));
 sky130_fd_sc_hd__o221a_1 _3747_ (.A1(_3334_),
    .A2(_3357_),
    .B1(_3346_),
    .B2(\as2650.stack[2][8] ),
    .C1(_3358_),
    .X(_3359_));
 sky130_fd_sc_hd__a31o_2 _3748_ (.A1(_3338_),
    .A2(_3347_),
    .A3(_3356_),
    .B1(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__inv_2 _3749_ (.A(_3262_),
    .Y(_3361_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_3361_),
    .B(_3332_),
    .Y(_3362_));
 sky130_fd_sc_hd__or2_4 _3751_ (.A(_3169_),
    .B(_3177_),
    .X(_3363_));
 sky130_fd_sc_hd__or3_1 _3752_ (.A(_3160_),
    .B(_3165_),
    .C(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__nand2_2 _3753_ (.A(_3183_),
    .B(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__o211a_1 _3754_ (.A1(_3332_),
    .A2(_3360_),
    .B1(_3362_),
    .C1(_3365_),
    .X(_3366_));
 sky130_fd_sc_hd__and3_2 _3755_ (.A(_3153_),
    .B(_3183_),
    .C(_3235_),
    .X(_3367_));
 sky130_fd_sc_hd__a211o_1 _3756_ (.A1(_3237_),
    .A2(_3329_),
    .B1(_3366_),
    .C1(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__o21a_1 _3757_ (.A1(\as2650.r123[0][0] ),
    .A2(_3236_),
    .B1(_3368_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _3758_ (.A(\as2650.holding_reg[1] ),
    .B(_3279_),
    .X(_3369_));
 sky130_fd_sc_hd__nor2_1 _3759_ (.A(\as2650.holding_reg[1] ),
    .B(_3279_),
    .Y(_3370_));
 sky130_fd_sc_hd__nor2_2 _3760_ (.A(_3369_),
    .B(_3370_),
    .Y(_3371_));
 sky130_fd_sc_hd__o2bb2a_1 _3761_ (.A1_N(_3272_),
    .A2_N(_3309_),
    .B1(_3321_),
    .B2(_3308_),
    .X(_3372_));
 sky130_fd_sc_hd__or2_1 _3762_ (.A(_3371_),
    .B(_3372_),
    .X(_3373_));
 sky130_fd_sc_hd__nand2_1 _3763_ (.A(_3371_),
    .B(_3372_),
    .Y(_3374_));
 sky130_fd_sc_hd__nand2_2 _3764_ (.A(_3323_),
    .B(_3107_),
    .Y(_3375_));
 sky130_fd_sc_hd__a21o_1 _3765_ (.A1(_3373_),
    .A2(_3374_),
    .B1(_3375_),
    .X(_3376_));
 sky130_fd_sc_hd__nand2_1 _3766_ (.A(_3323_),
    .B(_3220_),
    .Y(_3377_));
 sky130_fd_sc_hd__nand2_2 _3767_ (.A(_3189_),
    .B(_3107_),
    .Y(_3378_));
 sky130_fd_sc_hd__o21bai_1 _3768_ (.A1(_3311_),
    .A2(_3309_),
    .B1_N(_3321_),
    .Y(_3379_));
 sky130_fd_sc_hd__xor2_1 _3769_ (.A(_3371_),
    .B(_3379_),
    .X(_3380_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(\as2650.holding_reg[1] ),
    .A1(_3279_),
    .S(_3168_),
    .X(_3381_));
 sky130_fd_sc_hd__o22a_1 _3771_ (.A1(_3378_),
    .A2(_3380_),
    .B1(_3381_),
    .B2(_3107_),
    .X(_3382_));
 sky130_fd_sc_hd__a21oi_1 _3772_ (.A1(_3323_),
    .A2(_3370_),
    .B1(_3318_),
    .Y(_3383_));
 sky130_fd_sc_hd__a31o_1 _3773_ (.A1(_3376_),
    .A2(_3377_),
    .A3(_3382_),
    .B1(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__o21a_1 _3774_ (.A1(_3221_),
    .A2(_3369_),
    .B1(_3384_),
    .X(_3385_));
 sky130_fd_sc_hd__or2_1 _3775_ (.A(\as2650.holding_reg[1] ),
    .B(_3175_),
    .X(_3386_));
 sky130_fd_sc_hd__o21ai_2 _3776_ (.A1(_3168_),
    .A2(_3279_),
    .B1(_3386_),
    .Y(_3387_));
 sky130_fd_sc_hd__or2_1 _3777_ (.A(_3324_),
    .B(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__xnor2_2 _3778_ (.A(_3385_),
    .B(_3388_),
    .Y(_3389_));
 sky130_fd_sc_hd__buf_2 _3779_ (.A(\as2650.r0[1] ),
    .X(_3390_));
 sky130_fd_sc_hd__buf_4 _3780_ (.A(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__mux2_2 _3781_ (.A0(\as2650.r123[2][2] ),
    .A1(\as2650.r123_2[2][2] ),
    .S(_3162_),
    .X(_3392_));
 sky130_fd_sc_hd__mux4_1 _3782_ (.A0(\as2650.r123[1][2] ),
    .A1(\as2650.r123[0][2] ),
    .A2(\as2650.r123_2[1][2] ),
    .A3(\as2650.r123_2[0][2] ),
    .S0(_3070_),
    .S1(_3161_),
    .X(_3393_));
 sky130_fd_sc_hd__and3_1 _3783_ (.A(_3072_),
    .B(_3185_),
    .C(_3393_),
    .X(_3394_));
 sky130_fd_sc_hd__a221o_4 _3784_ (.A1(\as2650.r0[2] ),
    .A2(_3167_),
    .B1(_3392_),
    .B2(_3109_),
    .C1(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__buf_4 _3785_ (.A(_3395_),
    .X(_3396_));
 sky130_fd_sc_hd__buf_4 _3786_ (.A(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__nor2_4 _3787_ (.A(_3049_),
    .B(_3205_),
    .Y(_3398_));
 sky130_fd_sc_hd__nor2_4 _3788_ (.A(_3203_),
    .B(_3196_),
    .Y(_3399_));
 sky130_fd_sc_hd__mux2_1 _3789_ (.A0(_3398_),
    .A1(_3399_),
    .S(_3244_),
    .X(_3400_));
 sky130_fd_sc_hd__xor2_4 _3790_ (.A(_3279_),
    .B(_3400_),
    .X(_3401_));
 sky130_fd_sc_hd__or2_1 _3791_ (.A(_3281_),
    .B(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__o211a_1 _3792_ (.A1(_3128_),
    .A2(_3201_),
    .B1(_3225_),
    .C1(_3402_),
    .X(_3403_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(_3194_),
    .Y(_3404_));
 sky130_fd_sc_hd__a211o_1 _3794_ (.A1(_3283_),
    .A2(_3397_),
    .B1(_3403_),
    .C1(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__o211a_1 _3795_ (.A1(_3195_),
    .A2(_3287_),
    .B1(_3405_),
    .C1(_3208_),
    .X(_3406_));
 sky130_fd_sc_hd__a21o_1 _3796_ (.A1(_3391_),
    .A2(_3296_),
    .B1(_3406_),
    .X(_0300_));
 sky130_fd_sc_hd__xnor2_4 _3797_ (.A(_3286_),
    .B(_3278_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21bo_1 _3798_ (.A1(_3287_),
    .A2(_3257_),
    .B1_N(_3258_),
    .X(_0302_));
 sky130_fd_sc_hd__xnor2_4 _3799_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__mux2_1 _3800_ (.A0(_0300_),
    .A1(_0303_),
    .S(_3256_),
    .X(_0304_));
 sky130_fd_sc_hd__nor2_1 _3801_ (.A(\as2650.idx_ctrl[1] ),
    .B(_3247_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21a_1 _3802_ (.A1(_3244_),
    .A2(_0305_),
    .B1(_3248_),
    .X(_0306_));
 sky130_fd_sc_hd__xor2_4 _3803_ (.A(_0301_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _3804_ (.A(_3165_),
    .B(_3327_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_2 _3805_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o21a_1 _3806_ (.A1(_3238_),
    .A2(_0307_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__o21ai_1 _3807_ (.A1(_3302_),
    .A2(_0304_),
    .B1(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__a21bo_2 _3808_ (.A1(_3328_),
    .A2(_3389_),
    .B1_N(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_4 _3809_ (.A(_3169_),
    .B(_3173_),
    .Y(_0313_));
 sky130_fd_sc_hd__buf_2 _3810_ (.A(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__mux4_2 _3811_ (.A0(\as2650.stack[7][9] ),
    .A1(\as2650.stack[4][9] ),
    .A2(\as2650.stack[5][9] ),
    .A3(\as2650.stack[6][9] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_0315_));
 sky130_fd_sc_hd__buf_4 _3812_ (.A(_3346_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_4 _3813_ (.A(\as2650.psu[2] ),
    .X(_0317_));
 sky130_fd_sc_hd__and3_1 _3814_ (.A(_0317_),
    .B(\as2650.stack[3][9] ),
    .C(_3335_),
    .X(_0318_));
 sky130_fd_sc_hd__o22a_1 _3815_ (.A1(\as2650.stack[0][9] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[1][9] ),
    .X(_0319_));
 sky130_fd_sc_hd__o221a_1 _3816_ (.A1(\as2650.stack[2][9] ),
    .A2(_0316_),
    .B1(_0318_),
    .B2(_3334_),
    .C1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__a21oi_4 _3817_ (.A1(_3338_),
    .A2(_0315_),
    .B1(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _3818_ (.A(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__o221a_1 _3819_ (.A1(_3391_),
    .A2(_0314_),
    .B1(_3332_),
    .B2(_0322_),
    .C1(_3365_),
    .X(_0323_));
 sky130_fd_sc_hd__a211o_1 _3820_ (.A1(_3237_),
    .A2(_0312_),
    .B1(_0323_),
    .C1(_3367_),
    .X(_0324_));
 sky130_fd_sc_hd__o21a_1 _3821_ (.A1(\as2650.r123[0][1] ),
    .A2(_3236_),
    .B1(_0324_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _3822_ (.A(\as2650.r0[2] ),
    .X(_0325_));
 sky130_fd_sc_hd__buf_4 _3823_ (.A(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__mux4_1 _3824_ (.A0(\as2650.stack[7][10] ),
    .A1(\as2650.stack[4][10] ),
    .A2(\as2650.stack[5][10] ),
    .A3(\as2650.stack[6][10] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _3825_ (.A(_0317_),
    .B(\as2650.stack[3][10] ),
    .C(_3335_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _3826_ (.A(_3355_),
    .X(_0329_));
 sky130_fd_sc_hd__o22a_1 _3827_ (.A1(\as2650.stack[0][10] ),
    .A2(_3352_),
    .B1(_0329_),
    .B2(\as2650.stack[1][10] ),
    .X(_0330_));
 sky130_fd_sc_hd__o221a_1 _3828_ (.A1(\as2650.stack[2][10] ),
    .A2(_0316_),
    .B1(_0328_),
    .B2(_3334_),
    .C1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__a21o_2 _3829_ (.A1(_3338_),
    .A2(_0327_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__o221a_1 _3830_ (.A1(_0326_),
    .A2(_0313_),
    .B1(_3332_),
    .B2(_0332_),
    .C1(_3365_),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _3831_ (.A(_3367_),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__o22a_2 _3832_ (.A1(_3240_),
    .A2(_3243_),
    .B1(_3275_),
    .B2(_3277_),
    .X(_0335_));
 sky130_fd_sc_hd__xor2_1 _3833_ (.A(_3395_),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nor3_1 _3834_ (.A(_3287_),
    .B(_3279_),
    .C(_3395_),
    .Y(_0337_));
 sky130_fd_sc_hd__o21a_1 _3835_ (.A1(_3286_),
    .A2(_3279_),
    .B1(_3395_),
    .X(_0338_));
 sky130_fd_sc_hd__or3_1 _3836_ (.A(_3248_),
    .B(_0337_),
    .C(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__o221a_2 _3837_ (.A1(_3249_),
    .A2(_3396_),
    .B1(_0336_),
    .B2(_3246_),
    .C1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__o32a_1 _3838_ (.A1(_3258_),
    .A2(_0337_),
    .A3(_0338_),
    .B1(_0336_),
    .B2(_3257_),
    .X(_0341_));
 sky130_fd_sc_hd__o21a_2 _3839_ (.A1(_3259_),
    .A2(_3396_),
    .B1(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _3840_ (.A(_3287_),
    .B(_3279_),
    .Y(_0343_));
 sky130_fd_sc_hd__a22o_1 _3841_ (.A1(_3398_),
    .A2(_0335_),
    .B1(_0343_),
    .B2(_3399_),
    .X(_0344_));
 sky130_fd_sc_hd__xnor2_4 _3842_ (.A(_3396_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _3843_ (.A(_3282_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a211o_1 _3844_ (.A1(_3131_),
    .A2(_3282_),
    .B1(_3283_),
    .C1(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_4 _3845_ (.A(\as2650.r0[3] ),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_2 _3846_ (.A0(\as2650.r123[2][3] ),
    .A1(\as2650.r123_2[2][3] ),
    .S(_3162_),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _3847_ (.A0(\as2650.r123[1][3] ),
    .A1(\as2650.r123[0][3] ),
    .A2(\as2650.r123_2[1][3] ),
    .A3(\as2650.r123_2[0][3] ),
    .S0(_3070_),
    .S1(_3161_),
    .X(_0350_));
 sky130_fd_sc_hd__and3_1 _3848_ (.A(_3072_),
    .B(_3185_),
    .C(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_4 _3849_ (.A1(_0348_),
    .A2(_3167_),
    .B1(_0349_),
    .B2(_3109_),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_4 _3850_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_4 _3851_ (.A(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _3852_ (.A(_3225_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_1 _3853_ (.A(_3176_),
    .B(_3191_),
    .Y(_0356_));
 sky130_fd_sc_hd__and3_1 _3854_ (.A(_3186_),
    .B(_0356_),
    .C(_3295_),
    .X(_0357_));
 sky130_fd_sc_hd__a32o_1 _3855_ (.A1(_3195_),
    .A2(_0347_),
    .A3(_0355_),
    .B1(_0357_),
    .B2(_3280_),
    .X(_0358_));
 sky130_fd_sc_hd__o221a_1 _3856_ (.A1(_0326_),
    .A2(_3208_),
    .B1(_3296_),
    .B2(_0358_),
    .C1(_3213_),
    .X(_0359_));
 sky130_fd_sc_hd__a211o_1 _3857_ (.A1(_3256_),
    .A2(_0342_),
    .B1(_0359_),
    .C1(_3302_),
    .X(_0360_));
 sky130_fd_sc_hd__o21a_1 _3858_ (.A1(_3238_),
    .A2(_0340_),
    .B1(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _3859_ (.A(\as2650.holding_reg[2] ),
    .B(_3396_),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_1 _3860_ (.A(\as2650.holding_reg[2] ),
    .B(_3396_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_2 _3861_ (.A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _3862_ (.A(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__and2_2 _3863_ (.A(_3323_),
    .B(_3170_),
    .X(_0366_));
 sky130_fd_sc_hd__o22ai_2 _3864_ (.A1(_3371_),
    .A2(_3372_),
    .B1(_3387_),
    .B2(_3369_),
    .Y(_0367_));
 sky130_fd_sc_hd__xnor2_1 _3865_ (.A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__a21oi_1 _3866_ (.A1(_3371_),
    .A2(_3379_),
    .B1(_3369_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_1 _3867_ (.A(_0364_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__mux2_1 _3868_ (.A0(\as2650.holding_reg[2] ),
    .A1(_3396_),
    .S(_3168_),
    .X(_0371_));
 sky130_fd_sc_hd__o221a_1 _3869_ (.A1(_3378_),
    .A2(_0370_),
    .B1(_0371_),
    .B2(_3107_),
    .C1(_3377_),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_1 _3870_ (.A1(_3375_),
    .A2(_0368_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__o211a_1 _3871_ (.A1(_3377_),
    .A2(_0363_),
    .B1(_0373_),
    .C1(_3221_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _3872_ (.A(_3221_),
    .B(_0362_),
    .Y(_0375_));
 sky130_fd_sc_hd__or3_1 _3873_ (.A(_0366_),
    .B(_0374_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o21ai_2 _3874_ (.A1(_3324_),
    .A2(_0365_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__mux2_2 _3875_ (.A0(_0361_),
    .A1(_0377_),
    .S(_3328_),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _3876_ (.A(_3237_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _3877_ (.A1(\as2650.r123[0][2] ),
    .A2(_3236_),
    .B1(_0334_),
    .B2(_0379_),
    .X(_0010_));
 sky130_fd_sc_hd__nand2_1 _3878_ (.A(\as2650.holding_reg[3] ),
    .B(_0353_),
    .Y(_0380_));
 sky130_fd_sc_hd__or2_1 _3879_ (.A(\as2650.holding_reg[3] ),
    .B(_0353_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_0380_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_2 _3881_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _3882_ (.A(\as2650.holding_reg[3] ),
    .B(_0353_),
    .X(_0384_));
 sky130_fd_sc_hd__o2bb2a_1 _3883_ (.A1_N(_0365_),
    .A2_N(_0367_),
    .B1(_0371_),
    .B2(_0363_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _3884_ (.A(_0383_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a21oi_1 _3885_ (.A1(_0383_),
    .A2(_0385_),
    .B1(_3375_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _3886_ (.A(_0363_),
    .B(_0369_),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_1 _3887_ (.A(_0362_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__xnor2_1 _3888_ (.A(_0383_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__mux2_1 _3889_ (.A0(\as2650.holding_reg[3] ),
    .A1(_0353_),
    .S(_3176_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3890_ (.A0(\as2650.holding_reg[3] ),
    .A1(_0353_),
    .S(_3202_),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _3891_ (.A1(_3220_),
    .A2(_0391_),
    .B1(_0392_),
    .B2(_3069_),
    .C1(_3319_),
    .X(_0393_));
 sky130_fd_sc_hd__a21o_1 _3892_ (.A1(_3312_),
    .A2(_0390_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a21o_1 _3893_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__o211a_1 _3894_ (.A1(_3221_),
    .A2(_0384_),
    .B1(_0395_),
    .C1(_3324_),
    .X(_0396_));
 sky130_fd_sc_hd__a21oi_4 _3895_ (.A1(_0366_),
    .A2(_0383_),
    .B1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _3896_ (.A(_3396_),
    .B(_0335_),
    .Y(_0398_));
 sky130_fd_sc_hd__xnor2_1 _3897_ (.A(_0398_),
    .B(_0352_),
    .Y(_0399_));
 sky130_fd_sc_hd__nor4_4 _3898_ (.A(_3286_),
    .B(_3278_),
    .C(_3395_),
    .D(_0352_),
    .Y(_0400_));
 sky130_fd_sc_hd__o31a_1 _3899_ (.A1(_3286_),
    .A2(_3279_),
    .A3(_3395_),
    .B1(_0352_),
    .X(_0401_));
 sky130_fd_sc_hd__or3_1 _3900_ (.A(_3248_),
    .B(_0400_),
    .C(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__o221a_2 _3901_ (.A1(_3249_),
    .A2(_0353_),
    .B1(_0399_),
    .B2(_3246_),
    .C1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _3902_ (.A(_3398_),
    .B(_3396_),
    .C(_0335_),
    .X(_0404_));
 sky130_fd_sc_hd__a21oi_2 _3903_ (.A1(_3399_),
    .A2(_0337_),
    .B1(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__xnor2_4 _3904_ (.A(_0353_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__or2_1 _3905_ (.A(_3281_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__o211a_1 _3906_ (.A1(_3135_),
    .A2(_3201_),
    .B1(_3225_),
    .C1(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_2 _3907_ (.A0(\as2650.r123[2][4] ),
    .A1(\as2650.r123_2[2][4] ),
    .S(\as2650.psl[4] ),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _3908_ (.A1(\as2650.r0[4] ),
    .A2(_3166_),
    .B1(_0409_),
    .B2(_3108_),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _3909_ (.A0(\as2650.r123[1][4] ),
    .A1(\as2650.r123[0][4] ),
    .A2(\as2650.r123_2[1][4] ),
    .A3(\as2650.r123_2[0][4] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_3161_),
    .X(_0411_));
 sky130_fd_sc_hd__and3_1 _3910_ (.A(_3072_),
    .B(_3185_),
    .C(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_2 _3911_ (.A(_0410_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__buf_6 _3912_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__o21ai_1 _3913_ (.A1(_3225_),
    .A2(_0414_),
    .B1(_3195_),
    .Y(_0415_));
 sky130_fd_sc_hd__o22a_1 _3914_ (.A1(_3195_),
    .A2(_3397_),
    .B1(_0408_),
    .B2(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__buf_4 _3915_ (.A(_0348_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(_0416_),
    .A1(_0417_),
    .S(_3296_),
    .X(_0418_));
 sky130_fd_sc_hd__or3_1 _3917_ (.A(_3258_),
    .B(_0400_),
    .C(_0401_),
    .X(_0419_));
 sky130_fd_sc_hd__o221a_2 _3918_ (.A1(_3259_),
    .A2(_0353_),
    .B1(_0399_),
    .B2(_3257_),
    .C1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(_0418_),
    .A1(_0420_),
    .S(_3256_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(_0403_),
    .A1(_0421_),
    .S(_3238_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_0309_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__o21ai_4 _3922_ (.A1(_0309_),
    .A2(_0397_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2b_4 _3923_ (.A_N(_3334_),
    .B(_3336_),
    .Y(_0425_));
 sky130_fd_sc_hd__o22a_1 _3924_ (.A1(\as2650.stack[3][11] ),
    .A2(_3342_),
    .B1(_3355_),
    .B2(\as2650.stack[1][11] ),
    .X(_0426_));
 sky130_fd_sc_hd__o221a_1 _3925_ (.A1(\as2650.stack[0][11] ),
    .A2(_3352_),
    .B1(_0316_),
    .B2(\as2650.stack[2][11] ),
    .C1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__o221a_1 _3926_ (.A1(\as2650.stack[4][11] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[5][11] ),
    .C1(_3338_),
    .X(_0428_));
 sky130_fd_sc_hd__o221a_1 _3927_ (.A1(\as2650.stack[7][11] ),
    .A2(_3342_),
    .B1(_0316_),
    .B2(\as2650.stack[6][11] ),
    .C1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a21oi_4 _3928_ (.A1(_0425_),
    .A2(_0427_),
    .B1(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _3929_ (.A(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__o221a_1 _3930_ (.A1(_0417_),
    .A2(_0314_),
    .B1(_3332_),
    .B2(_0431_),
    .C1(_3365_),
    .X(_0432_));
 sky130_fd_sc_hd__a211o_1 _3931_ (.A1(_3237_),
    .A2(_0424_),
    .B1(_0432_),
    .C1(_3367_),
    .X(_0433_));
 sky130_fd_sc_hd__o21a_1 _3932_ (.A1(\as2650.r123[0][3] ),
    .A2(_3236_),
    .B1(_0433_),
    .X(_0011_));
 sky130_fd_sc_hd__inv_2 _3933_ (.A(\as2650.holding_reg[4] ),
    .Y(_0434_));
 sky130_fd_sc_hd__mux2_1 _3934_ (.A0(_0434_),
    .A1(_0414_),
    .S(_3176_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_2 _3935_ (.A(_3324_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(_0434_),
    .B(_0414_),
    .Y(_0437_));
 sky130_fd_sc_hd__or2_1 _3937_ (.A(_0410_),
    .B(_0412_),
    .X(_0438_));
 sky130_fd_sc_hd__buf_4 _3938_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_1 _3939_ (.A(\as2650.holding_reg[4] ),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_2 _3940_ (.A(_0437_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__o31a_1 _3941_ (.A1(_0362_),
    .A2(_0384_),
    .A3(_0388_),
    .B1(_0381_),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21a_1 _3943_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_3312_),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_0380_),
    .B(_0391_),
    .Y(_0445_));
 sky130_fd_sc_hd__a31o_1 _3945_ (.A1(_0386_),
    .A2(_0441_),
    .A3(_0445_),
    .B1(_3375_),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _3946_ (.A1(_0386_),
    .A2(_0445_),
    .B1(_0441_),
    .X(_0447_));
 sky130_fd_sc_hd__and2b_1 _3947_ (.A_N(_0446_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__inv_2 _3948_ (.A(_0435_),
    .Y(_0449_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\as2650.holding_reg[4] ),
    .A1(_0439_),
    .S(_3202_),
    .X(_0450_));
 sky130_fd_sc_hd__a221o_1 _3950_ (.A1(_3220_),
    .A2(_0449_),
    .B1(_0450_),
    .B2(_3069_),
    .C1(_3319_),
    .X(_0451_));
 sky130_fd_sc_hd__a211o_1 _3951_ (.A1(_0443_),
    .A2(_0444_),
    .B1(_0448_),
    .C1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_2 _3952_ (.A1(_3221_),
    .A2(_0437_),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__xnor2_4 _3953_ (.A(_0436_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__mux2_2 _3954_ (.A0(\as2650.r123[2][5] ),
    .A1(\as2650.r123_2[2][5] ),
    .S(_3162_),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _3955_ (.A1(\as2650.r0[5] ),
    .A2(_3167_),
    .B1(_0455_),
    .B2(_3109_),
    .X(_0456_));
 sky130_fd_sc_hd__mux4_1 _3956_ (.A0(\as2650.r123[1][5] ),
    .A1(\as2650.r123[0][5] ),
    .A2(\as2650.r123_2[1][5] ),
    .A3(\as2650.r123_2[0][5] ),
    .S0(_3070_),
    .S1(_3162_),
    .X(_0457_));
 sky130_fd_sc_hd__and3_1 _3957_ (.A(_3073_),
    .B(_3185_),
    .C(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__or2_1 _3958_ (.A(_0456_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_4 _3959_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _3960_ (.A(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _3961_ (.A1(_0404_),
    .A2(_0353_),
    .B1(_0400_),
    .B2(_3399_),
    .X(_0462_));
 sky130_fd_sc_hd__xnor2_2 _3962_ (.A(_0414_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__or2_1 _3963_ (.A(_3282_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__clkinv_4 _3964_ (.A(net5),
    .Y(_0465_));
 sky130_fd_sc_hd__a21oi_1 _3965_ (.A1(_0465_),
    .A2(_3282_),
    .B1(_3283_),
    .Y(_0466_));
 sky130_fd_sc_hd__a22o_1 _3966_ (.A1(_3283_),
    .A2(_0461_),
    .B1(_0464_),
    .B2(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(_0354_),
    .A1(_0467_),
    .S(_3195_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_2 _3968_ (.A(\as2650.r0[4] ),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _3969_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(_0468_),
    .A1(_0470_),
    .S(_3296_),
    .X(_0471_));
 sky130_fd_sc_hd__xnor2_1 _3971_ (.A(_0413_),
    .B(_0400_),
    .Y(_0472_));
 sky130_fd_sc_hd__and4_1 _3972_ (.A(_3395_),
    .B(_0335_),
    .C(_0352_),
    .D(_0439_),
    .X(_0473_));
 sky130_fd_sc_hd__a31o_1 _3973_ (.A1(_3395_),
    .A2(_0335_),
    .A3(_0352_),
    .B1(_0439_),
    .X(_0474_));
 sky130_fd_sc_hd__or2b_1 _3974_ (.A(_0473_),
    .B_N(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__or2b_1 _3975_ (.A(_3257_),
    .B_N(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__o221a_2 _3976_ (.A1(_3259_),
    .A2(_0439_),
    .B1(_0472_),
    .B2(_3258_),
    .C1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(_0471_),
    .A1(_0477_),
    .S(_3256_),
    .X(_0478_));
 sky130_fd_sc_hd__nand2_1 _3978_ (.A(_0305_),
    .B(_0475_),
    .Y(_0479_));
 sky130_fd_sc_hd__o221a_2 _3979_ (.A1(_3249_),
    .A2(_0439_),
    .B1(_0472_),
    .B2(_3248_),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__a21o_1 _3980_ (.A1(_3302_),
    .A2(_0480_),
    .B1(_3328_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_1 _3981_ (.A1(_3238_),
    .A2(_0478_),
    .B1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_2 _3982_ (.A1(_0309_),
    .A2(_0454_),
    .B1(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__mux4_1 _3983_ (.A0(\as2650.stack[7][12] ),
    .A1(\as2650.stack[4][12] ),
    .A2(\as2650.stack[5][12] ),
    .A3(\as2650.stack[6][12] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _3984_ (.A(_0317_),
    .B(\as2650.stack[3][12] ),
    .C(_3335_),
    .X(_0485_));
 sky130_fd_sc_hd__o22a_1 _3985_ (.A1(\as2650.stack[0][12] ),
    .A2(_3352_),
    .B1(_0329_),
    .B2(\as2650.stack[1][12] ),
    .X(_0486_));
 sky130_fd_sc_hd__o221a_1 _3986_ (.A1(\as2650.stack[2][12] ),
    .A2(_0316_),
    .B1(_0485_),
    .B2(_3334_),
    .C1(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a21o_2 _3987_ (.A1(_3338_),
    .A2(_0484_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__o221a_1 _3988_ (.A1(_0470_),
    .A2(_0314_),
    .B1(_3332_),
    .B2(_0488_),
    .C1(_3365_),
    .X(_0489_));
 sky130_fd_sc_hd__a211o_1 _3989_ (.A1(_3237_),
    .A2(_0483_),
    .B1(_0489_),
    .C1(_3367_),
    .X(_0490_));
 sky130_fd_sc_hd__o21a_1 _3990_ (.A1(\as2650.r123[0][4] ),
    .A2(_3236_),
    .B1(_0490_),
    .X(_0012_));
 sky130_fd_sc_hd__nor2_4 _3991_ (.A(_0456_),
    .B(_0458_),
    .Y(_0491_));
 sky130_fd_sc_hd__and3_2 _3992_ (.A(_0413_),
    .B(_0400_),
    .C(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_1 _3993_ (.A1(_0414_),
    .A2(_0400_),
    .B1(_0491_),
    .Y(_0493_));
 sky130_fd_sc_hd__or2_1 _3994_ (.A(_0492_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _3995_ (.A(_0460_),
    .B(_0473_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_1 _3996_ (.A(_0460_),
    .B(_0473_),
    .Y(_0496_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_0495_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__or2_1 _3998_ (.A(_3246_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o221a_2 _3999_ (.A1(_3249_),
    .A2(_0460_),
    .B1(_0494_),
    .B2(_3248_),
    .C1(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_2 _4000_ (.A0(\as2650.r123[2][6] ),
    .A1(\as2650.r123_2[2][6] ),
    .S(_3162_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _4001_ (.A1(\as2650.r0[6] ),
    .A2(_3167_),
    .B1(_0500_),
    .B2(_3109_),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _4002_ (.A0(\as2650.r123[1][6] ),
    .A1(\as2650.r123[0][6] ),
    .A2(\as2650.r123_2[1][6] ),
    .A3(\as2650.r123_2[0][6] ),
    .S0(_3178_),
    .S1(_3163_),
    .X(_0502_));
 sky130_fd_sc_hd__and3_1 _4003_ (.A(_3073_),
    .B(_3185_),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__nor2_4 _4004_ (.A(_0501_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__and3_1 _4005_ (.A(_3399_),
    .B(_0414_),
    .C(_0400_),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _4006_ (.A1(_3398_),
    .A2(_0473_),
    .B1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__xnor2_4 _4007_ (.A(_0460_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(_3139_),
    .B(_3201_),
    .Y(_0508_));
 sky130_fd_sc_hd__a211o_1 _4009_ (.A1(_3201_),
    .A2(_0507_),
    .B1(_0508_),
    .C1(_3283_),
    .X(_0509_));
 sky130_fd_sc_hd__o211a_1 _4010_ (.A1(_3225_),
    .A2(_0504_),
    .B1(_0509_),
    .C1(_3195_),
    .X(_0510_));
 sky130_fd_sc_hd__a21oi_1 _4011_ (.A1(_3264_),
    .A2(_0414_),
    .B1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__buf_2 _4012_ (.A(\as2650.r0[5] ),
    .X(_0512_));
 sky130_fd_sc_hd__buf_4 _4013_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(_0511_),
    .A1(_0513_),
    .S(_3296_),
    .X(_0514_));
 sky130_fd_sc_hd__or2_1 _4015_ (.A(_3257_),
    .B(_0497_),
    .X(_0515_));
 sky130_fd_sc_hd__o221a_2 _4016_ (.A1(_3259_),
    .A2(_0460_),
    .B1(_0494_),
    .B2(_3258_),
    .C1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(_0514_),
    .A1(_0516_),
    .S(_3256_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(_0499_),
    .A1(_0517_),
    .S(_3238_),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(\as2650.holding_reg[5] ),
    .B(_0460_),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _4020_ (.A(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(\as2650.holding_reg[5] ),
    .B(_0460_),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_2 _4022_ (.A(_0520_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21oi_1 _4023_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0437_),
    .Y(_0523_));
 sky130_fd_sc_hd__xor2_1 _4024_ (.A(_0522_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(_0435_),
    .B(_0437_),
    .X(_0525_));
 sky130_fd_sc_hd__and3_1 _4026_ (.A(_0447_),
    .B(_0522_),
    .C(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__a21o_1 _4027_ (.A1(_0447_),
    .A2(_0525_),
    .B1(_0522_),
    .X(_0527_));
 sky130_fd_sc_hd__or3b_1 _4028_ (.A(_3375_),
    .B(_0526_),
    .C_N(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(\as2650.holding_reg[5] ),
    .B(_3176_),
    .X(_0529_));
 sky130_fd_sc_hd__o21a_1 _4030_ (.A1(_3202_),
    .A2(_0461_),
    .B1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(\as2650.holding_reg[5] ),
    .A1(_0461_),
    .S(_3202_),
    .X(_0531_));
 sky130_fd_sc_hd__a221oi_1 _4032_ (.A1(_3220_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_3069_),
    .C1(_3319_),
    .Y(_0532_));
 sky130_fd_sc_hd__o211a_1 _4033_ (.A1(_3378_),
    .A2(_0524_),
    .B1(_0528_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__a21o_1 _4034_ (.A1(_3319_),
    .A2(_0519_),
    .B1(_0366_),
    .X(_0534_));
 sky130_fd_sc_hd__a2bb2o_2 _4035_ (.A1_N(_0533_),
    .A2_N(_0534_),
    .B1(_0366_),
    .B2(_0522_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_2 _4036_ (.A0(_0518_),
    .A1(_0535_),
    .S(_3328_),
    .X(_0536_));
 sky130_fd_sc_hd__o22a_1 _4037_ (.A1(\as2650.stack[3][13] ),
    .A2(_3342_),
    .B1(_3346_),
    .B2(\as2650.stack[2][13] ),
    .X(_0537_));
 sky130_fd_sc_hd__o221a_1 _4038_ (.A1(\as2650.stack[0][13] ),
    .A2(_3352_),
    .B1(_0329_),
    .B2(\as2650.stack[1][13] ),
    .C1(_0425_),
    .X(_0538_));
 sky130_fd_sc_hd__o22a_1 _4039_ (.A1(\as2650.stack[7][13] ),
    .A2(_3342_),
    .B1(_3346_),
    .B2(\as2650.stack[6][13] ),
    .X(_0539_));
 sky130_fd_sc_hd__o221a_1 _4040_ (.A1(\as2650.stack[4][13] ),
    .A2(_3352_),
    .B1(_0329_),
    .B2(\as2650.stack[5][13] ),
    .C1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__a22o_2 _4041_ (.A1(_0537_),
    .A2(_0538_),
    .B1(_0540_),
    .B2(_3338_),
    .X(_0541_));
 sky130_fd_sc_hd__o221a_1 _4042_ (.A1(_0513_),
    .A2(_0313_),
    .B1(_3332_),
    .B2(_0541_),
    .C1(_3365_),
    .X(_0542_));
 sky130_fd_sc_hd__a211o_1 _4043_ (.A1(_3237_),
    .A2(_0536_),
    .B1(_0542_),
    .C1(_3367_),
    .X(_0543_));
 sky130_fd_sc_hd__o21a_1 _4044_ (.A1(\as2650.r123[0][5] ),
    .A2(_3236_),
    .B1(_0543_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _4045_ (.A(\as2650.r0[6] ),
    .X(_0544_));
 sky130_fd_sc_hd__buf_4 _4046_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__o22a_1 _4047_ (.A1(\as2650.stack[7][14] ),
    .A2(_3342_),
    .B1(_3345_),
    .B2(\as2650.stack[6][14] ),
    .X(_0546_));
 sky130_fd_sc_hd__o221a_1 _4048_ (.A1(\as2650.stack[4][14] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[5][14] ),
    .C1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o22a_1 _4049_ (.A1(\as2650.stack[3][14] ),
    .A2(_3342_),
    .B1(_3346_),
    .B2(\as2650.stack[2][14] ),
    .X(_0548_));
 sky130_fd_sc_hd__o221a_1 _4050_ (.A1(\as2650.stack[0][14] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[1][14] ),
    .C1(_0425_),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_2 _4051_ (.A1(_3338_),
    .A2(_0547_),
    .B1(_0548_),
    .B2(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__o221a_1 _4052_ (.A1(_0545_),
    .A2(_0313_),
    .B1(_3332_),
    .B2(_0550_),
    .C1(_3365_),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _4053_ (.A(_3367_),
    .B(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _4054_ (.A(_0501_),
    .B(_0503_),
    .X(_0553_));
 sky130_fd_sc_hd__buf_2 _4055_ (.A(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__nand2_1 _4056_ (.A(\as2650.holding_reg[6] ),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__or2_1 _4057_ (.A(\as2650.holding_reg[6] ),
    .B(_0554_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__and2_1 _4059_ (.A(_0555_),
    .B(_0556_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(_0519_),
    .B(_0530_),
    .Y(_0559_));
 sky130_fd_sc_hd__and3_1 _4061_ (.A(_0527_),
    .B(_0558_),
    .C(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _4062_ (.A1(_0527_),
    .A2(_0559_),
    .B1(_0558_),
    .Y(_0561_));
 sky130_fd_sc_hd__or3_1 _4063_ (.A(_3375_),
    .B(_0560_),
    .C(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__o21ai_1 _4064_ (.A1(_0521_),
    .A2(_0523_),
    .B1(_0519_),
    .Y(_0563_));
 sky130_fd_sc_hd__xnor2_1 _4065_ (.A(_0557_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(\as2650.holding_reg[6] ),
    .A1(_0554_),
    .S(_3176_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_4 _4067_ (.A(_0554_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _4068_ (.A0(\as2650.holding_reg[6] ),
    .A1(_0566_),
    .S(_3202_),
    .X(_0567_));
 sky130_fd_sc_hd__a221o_1 _4069_ (.A1(_3220_),
    .A2(_0565_),
    .B1(_0567_),
    .B2(_3069_),
    .C1(_3319_),
    .X(_0568_));
 sky130_fd_sc_hd__a21oi_1 _4070_ (.A1(_3312_),
    .A2(_0564_),
    .B1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__a221o_1 _4071_ (.A1(_3319_),
    .A2(_0555_),
    .B1(_0562_),
    .B2(_0569_),
    .C1(_0366_),
    .X(_0570_));
 sky130_fd_sc_hd__o21a_1 _4072_ (.A1(_3324_),
    .A2(_0557_),
    .B1(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__and3_1 _4073_ (.A(_0460_),
    .B(_0473_),
    .C(_0554_),
    .X(_0572_));
 sky130_fd_sc_hd__nor2_1 _4074_ (.A(_0495_),
    .B(_0554_),
    .Y(_0573_));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_0572_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__xnor2_1 _4076_ (.A(_0492_),
    .B(_0504_),
    .Y(_0575_));
 sky130_fd_sc_hd__or2_1 _4077_ (.A(_3248_),
    .B(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__o221a_2 _4078_ (.A1(_3249_),
    .A2(_0554_),
    .B1(_0574_),
    .B2(_3246_),
    .C1(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__or2_1 _4079_ (.A(_3258_),
    .B(_0575_),
    .X(_0578_));
 sky130_fd_sc_hd__o221a_2 _4080_ (.A1(_3259_),
    .A2(_0554_),
    .B1(_0574_),
    .B2(_3257_),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a21oi_1 _4081_ (.A1(_3398_),
    .A2(_0495_),
    .B1(_0554_),
    .Y(_0580_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(_3399_),
    .A2(_0492_),
    .B1(_0572_),
    .B2(_3398_),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _4083_ (.A(_0413_),
    .B(_0491_),
    .C(_0504_),
    .X(_0582_));
 sky130_fd_sc_hd__and3_1 _4084_ (.A(_3399_),
    .B(_0400_),
    .C(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__o21ba_1 _4085_ (.A1(_0580_),
    .A2(_0581_),
    .B1_N(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__nor2_1 _4086_ (.A(_3282_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__a211o_1 _4087_ (.A1(_3144_),
    .A2(_3282_),
    .B1(_3283_),
    .C1(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__o211a_1 _4088_ (.A1(_3225_),
    .A2(_3271_),
    .B1(_0586_),
    .C1(_3195_),
    .X(_0587_));
 sky130_fd_sc_hd__a211o_1 _4089_ (.A1(_0357_),
    .A2(_0461_),
    .B1(_0587_),
    .C1(_3296_),
    .X(_0588_));
 sky130_fd_sc_hd__o211a_1 _4090_ (.A1(_0545_),
    .A2(_3208_),
    .B1(_3213_),
    .C1(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__a211o_1 _4091_ (.A1(_3256_),
    .A2(_0579_),
    .B1(_0589_),
    .C1(_3302_),
    .X(_0590_));
 sky130_fd_sc_hd__o211ai_1 _4092_ (.A1(_3238_),
    .A2(_0577_),
    .B1(_0590_),
    .C1(_0309_),
    .Y(_0591_));
 sky130_fd_sc_hd__o21ai_2 _4093_ (.A1(_0309_),
    .A2(_0571_),
    .B1(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__and2_1 _4094_ (.A(_3237_),
    .B(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__o22a_1 _4095_ (.A1(\as2650.r123[0][6] ),
    .A2(_3236_),
    .B1(_0552_),
    .B2(_0593_),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_1 _4096_ (.A(\as2650.holding_reg[7] ),
    .B(_3271_),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _4097_ (.A(\as2650.holding_reg[7] ),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_4 _4098_ (.A(_3266_),
    .B(_3268_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _4099_ (.A(_0595_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__and2_1 _4100_ (.A(_0594_),
    .B(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__and2_1 _4101_ (.A(_0555_),
    .B(_0565_),
    .X(_0599_));
 sky130_fd_sc_hd__or3_1 _4102_ (.A(_0561_),
    .B(_0598_),
    .C(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__o21ai_1 _4103_ (.A1(_0561_),
    .A2(_0599_),
    .B1(_0598_),
    .Y(_0601_));
 sky130_fd_sc_hd__a21o_1 _4104_ (.A1(_0600_),
    .A2(_0601_),
    .B1(_3375_),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_1 _4105_ (.A(_0594_),
    .B(_0597_),
    .Y(_0603_));
 sky130_fd_sc_hd__a21boi_1 _4106_ (.A1(_0558_),
    .A2(_0563_),
    .B1_N(_0555_),
    .Y(_0604_));
 sky130_fd_sc_hd__xnor2_1 _4107_ (.A(_0603_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(_0595_),
    .A1(_0596_),
    .S(_3202_),
    .X(_0606_));
 sky130_fd_sc_hd__o221a_1 _4109_ (.A1(_3378_),
    .A2(_0605_),
    .B1(_0606_),
    .B2(_3107_),
    .C1(_3377_),
    .X(_0607_));
 sky130_fd_sc_hd__a21oi_1 _4110_ (.A1(_3323_),
    .A2(_0597_),
    .B1(_3318_),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_1 _4111_ (.A1(_0602_),
    .A2(_0607_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__a31o_1 _4112_ (.A1(\as2650.holding_reg[7] ),
    .A2(_3319_),
    .A3(_3271_),
    .B1(_0366_),
    .X(_0610_));
 sky130_fd_sc_hd__o22a_2 _4113_ (.A1(_3324_),
    .A2(_0598_),
    .B1(_0609_),
    .B2(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__xnor2_1 _4114_ (.A(_0596_),
    .B(_0572_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _4115_ (.A(_0400_),
    .B(_0582_),
    .Y(_0613_));
 sky130_fd_sc_hd__xnor2_1 _4116_ (.A(_3270_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__or2_1 _4117_ (.A(_3270_),
    .B(_3249_),
    .X(_0615_));
 sky130_fd_sc_hd__o221a_2 _4118_ (.A1(_3246_),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_3248_),
    .C1(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _4119_ (.A(\as2650.r0[7] ),
    .X(_0617_));
 sky130_fd_sc_hd__buf_4 _4120_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__o21a_2 _4121_ (.A1(\as2650.psl[3] ),
    .A2(_3287_),
    .B1(_3272_),
    .X(_0619_));
 sky130_fd_sc_hd__a31o_1 _4122_ (.A1(_3398_),
    .A2(_0495_),
    .A3(_0554_),
    .B1(_0583_),
    .X(_0620_));
 sky130_fd_sc_hd__xnor2_2 _4123_ (.A(_3270_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _4124_ (.A(_3282_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__a211o_1 _4125_ (.A1(_3146_),
    .A2(_3282_),
    .B1(_3283_),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__o211a_1 _4126_ (.A1(_3225_),
    .A2(_0619_),
    .B1(_0623_),
    .C1(_3195_),
    .X(_0624_));
 sky130_fd_sc_hd__a211o_1 _4127_ (.A1(_3264_),
    .A2(_0566_),
    .B1(_0624_),
    .C1(_3296_),
    .X(_0625_));
 sky130_fd_sc_hd__o21a_1 _4128_ (.A1(_0618_),
    .A2(_3208_),
    .B1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or2_1 _4129_ (.A(_3270_),
    .B(_3259_),
    .X(_0627_));
 sky130_fd_sc_hd__o221a_4 _4130_ (.A1(_3257_),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_3258_),
    .C1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__o221a_1 _4131_ (.A1(_3256_),
    .A2(_0626_),
    .B1(_0628_),
    .B2(_3213_),
    .C1(_3218_),
    .X(_0629_));
 sky130_fd_sc_hd__a211o_1 _4132_ (.A1(_3302_),
    .A2(_0616_),
    .B1(_0629_),
    .C1(_3328_),
    .X(_0630_));
 sky130_fd_sc_hd__o21a_1 _4133_ (.A1(_0309_),
    .A2(_0611_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__a31o_1 _4134_ (.A1(_0618_),
    .A2(_3331_),
    .A3(_3365_),
    .B1(_3367_),
    .X(_0632_));
 sky130_fd_sc_hd__a21o_1 _4135_ (.A1(_3237_),
    .A2(_0631_),
    .B1(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__o21a_1 _4136_ (.A1(\as2650.r123[0][7] ),
    .A2(_3236_),
    .B1(_0633_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_4 _4137_ (.A(_3262_),
    .X(_0634_));
 sky130_fd_sc_hd__buf_2 _4138_ (.A(\as2650.pc[0] ),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_4 _4139_ (.A(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__inv_2 _4140_ (.A(_0317_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_2 _4141_ (.A(_3155_),
    .B(_3042_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_2 _4142_ (.A(_3151_),
    .B(_3097_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__clkbuf_4 _4144_ (.A(_3111_),
    .X(_0641_));
 sky130_fd_sc_hd__o22a_1 _4145_ (.A1(_3147_),
    .A2(_3084_),
    .B1(_0640_),
    .B2(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_2 _4146_ (.A(_3227_),
    .B(_3076_),
    .Y(_0643_));
 sky130_fd_sc_hd__or2b_1 _4147_ (.A(_3196_),
    .B_N(_3203_),
    .X(_0644_));
 sky130_fd_sc_hd__or3_1 _4148_ (.A(_0642_),
    .B(_0643_),
    .C(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_2 _4149_ (.A(_3065_),
    .B(_3110_),
    .Y(_0646_));
 sky130_fd_sc_hd__buf_4 _4150_ (.A(_3097_),
    .X(_0647_));
 sky130_fd_sc_hd__or3_1 _4151_ (.A(_3189_),
    .B(_0646_),
    .C(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__a21o_1 _4152_ (.A1(_0645_),
    .A2(_0648_),
    .B1(_3056_),
    .X(_0649_));
 sky130_fd_sc_hd__or3_1 _4153_ (.A(_0637_),
    .B(_3352_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__buf_4 _4154_ (.A(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _4155_ (.A0(_0636_),
    .A1(\as2650.stack[5][0] ),
    .S(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__nor3_4 _4156_ (.A(_3176_),
    .B(_3173_),
    .C(_3180_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_4 _4157_ (.A(_3120_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__or2_1 _4158_ (.A(_3056_),
    .B(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__or3_1 _4159_ (.A(_0637_),
    .B(_0329_),
    .C(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__buf_4 _4160_ (.A(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(_0634_),
    .A1(_0652_),
    .S(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _4162_ (.A(_0658_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _4163_ (.A(_3391_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_2 _4164_ (.A(\as2650.pc[1] ),
    .X(_0660_));
 sky130_fd_sc_hd__buf_4 _4165_ (.A(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(_0661_),
    .A1(\as2650.stack[5][1] ),
    .S(_0651_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(_0659_),
    .A1(_0662_),
    .S(_0657_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _4168_ (.A(_0663_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _4169_ (.A(_0326_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(\as2650.pc[2] ),
    .A1(\as2650.stack[5][2] ),
    .S(_0651_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(_0664_),
    .A1(_0665_),
    .S(_0657_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_1 _4172_ (.A(_0666_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _4173_ (.A(_0417_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_4 _4174_ (.A(\as2650.pc[3] ),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(_0668_),
    .A1(\as2650.stack[5][3] ),
    .S(_0651_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(_0667_),
    .A1(_0669_),
    .S(_0657_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _4177_ (.A(_0670_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _4178_ (.A(_0470_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_4 _4179_ (.A(\as2650.pc[4] ),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(_0672_),
    .A1(\as2650.stack[5][4] ),
    .S(_0651_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(_0671_),
    .A1(_0673_),
    .S(_0657_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _4182_ (.A(_0674_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_4 _4183_ (.A(_0513_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_4 _4184_ (.A(\as2650.pc[5] ),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(_0676_),
    .A1(\as2650.stack[5][5] ),
    .S(_0651_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(_0675_),
    .A1(_0677_),
    .S(_0657_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _4187_ (.A(_0678_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_4 _4188_ (.A(_0545_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_4 _4189_ (.A(\as2650.pc[6] ),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_4 _4190_ (.A(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(_0681_),
    .A1(\as2650.stack[5][6] ),
    .S(_0651_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(_0679_),
    .A1(_0682_),
    .S(_0657_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _4193_ (.A(_0683_),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_4 _4194_ (.A(_0618_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_4 _4195_ (.A(\as2650.pc[7] ),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _4196_ (.A0(_0685_),
    .A1(\as2650.stack[5][7] ),
    .S(_0651_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(_0684_),
    .A1(_0686_),
    .S(_0657_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _4198_ (.A(_0687_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_2 _4199_ (.A(_3165_),
    .B(_0654_),
    .Y(_0688_));
 sky130_fd_sc_hd__buf_4 _4200_ (.A(\as2650.pc[8] ),
    .X(_0689_));
 sky130_fd_sc_hd__buf_4 _4201_ (.A(_3102_),
    .X(_0690_));
 sky130_fd_sc_hd__buf_4 _4202_ (.A(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_1 _4203_ (.A(_0691_),
    .B(_0653_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor3_2 _4204_ (.A(_3184_),
    .B(_3056_),
    .C(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(\as2650.r123[0][0] ),
    .A1(\as2650.r123_2[0][0] ),
    .S(_3162_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_2 _4206_ (.A(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_4 _4207_ (.A(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__buf_4 _4208_ (.A(_0655_),
    .X(_0697_));
 sky130_fd_sc_hd__o22a_1 _4209_ (.A1(_0689_),
    .A2(_0693_),
    .B1(_0696_),
    .B2(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__a21o_2 _4210_ (.A1(\as2650.r123[0][0] ),
    .A2(_0688_),
    .B1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__buf_4 _4211_ (.A(_0637_),
    .X(_0700_));
 sky130_fd_sc_hd__or3_4 _4212_ (.A(_0700_),
    .B(_0329_),
    .C(_0649_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_4 _4213_ (.A(_0657_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(\as2650.stack[6][8] ),
    .A1(_0699_),
    .S(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_1 _4215_ (.A(_0703_),
    .X(_0024_));
 sky130_fd_sc_hd__buf_4 _4216_ (.A(\as2650.pc[9] ),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(\as2650.r123[0][1] ),
    .A1(\as2650.r123_2[0][1] ),
    .S(_3162_),
    .X(_0705_));
 sky130_fd_sc_hd__clkbuf_2 _4218_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_4 _4219_ (.A(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__o22a_1 _4220_ (.A1(_0704_),
    .A2(_0693_),
    .B1(_0707_),
    .B2(_0697_),
    .X(_0708_));
 sky130_fd_sc_hd__a21o_2 _4221_ (.A1(\as2650.r123[0][1] ),
    .A2(_0688_),
    .B1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _4222_ (.A0(\as2650.stack[6][9] ),
    .A1(_0709_),
    .S(_0702_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _4223_ (.A(_0710_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_2 _4224_ (.A0(\as2650.r123[0][2] ),
    .A1(\as2650.r123_2[0][2] ),
    .S(_3161_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_4 _4225_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__buf_4 _4226_ (.A(\as2650.pc[10] ),
    .X(_0713_));
 sky130_fd_sc_hd__o22a_1 _4227_ (.A1(_0712_),
    .A2(_0697_),
    .B1(_0693_),
    .B2(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_2 _4228_ (.A1(\as2650.r123[0][2] ),
    .A2(_0688_),
    .B1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(\as2650.stack[6][10] ),
    .A1(_0715_),
    .S(_0702_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _4230_ (.A(_0716_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_2 _4231_ (.A0(\as2650.r123[0][3] ),
    .A1(\as2650.r123_2[0][3] ),
    .S(_3161_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_4 _4232_ (.A(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_4 _4233_ (.A(\as2650.pc[11] ),
    .X(_0719_));
 sky130_fd_sc_hd__o22a_1 _4234_ (.A1(_0718_),
    .A2(_0697_),
    .B1(_0693_),
    .B2(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__a21o_2 _4235_ (.A1(\as2650.r123[0][3] ),
    .A2(_0688_),
    .B1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(\as2650.stack[6][11] ),
    .A1(_0721_),
    .S(_0702_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_1 _4237_ (.A(_0722_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(\as2650.r123[0][4] ),
    .A1(\as2650.r123_2[0][4] ),
    .S(_3161_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_4 _4239_ (.A(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__clkbuf_4 _4240_ (.A(_0655_),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _4241_ (.A(\as2650.pc[12] ),
    .X(_0726_));
 sky130_fd_sc_hd__o22a_1 _4242_ (.A1(_0724_),
    .A2(_0725_),
    .B1(_0693_),
    .B2(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_2 _4243_ (.A1(\as2650.r123[0][4] ),
    .A2(_0688_),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(\as2650.stack[6][12] ),
    .A1(_0728_),
    .S(_0702_),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_1 _4245_ (.A(_0729_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_2 _4246_ (.A0(\as2650.r123[0][5] ),
    .A1(\as2650.r123_2[0][5] ),
    .S(_3162_),
    .X(_0730_));
 sky130_fd_sc_hd__buf_2 _4247_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__o22a_1 _4248_ (.A1(_0731_),
    .A2(_0725_),
    .B1(_0693_),
    .B2(\as2650.pc[13] ),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_2 _4249_ (.A1(\as2650.r123[0][5] ),
    .A2(_0688_),
    .B1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(\as2650.stack[6][13] ),
    .A1(_0733_),
    .S(_0702_),
    .X(_0734_));
 sky130_fd_sc_hd__clkbuf_1 _4251_ (.A(_0734_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_2 _4252_ (.A0(\as2650.r123[0][6] ),
    .A1(\as2650.r123_2[0][6] ),
    .S(_3162_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_4 _4253_ (.A(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__o22a_1 _4254_ (.A1(_0736_),
    .A2(_0725_),
    .B1(_0693_),
    .B2(\as2650.pc[14] ),
    .X(_0737_));
 sky130_fd_sc_hd__a21o_2 _4255_ (.A1(\as2650.r123[0][6] ),
    .A2(_0688_),
    .B1(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\as2650.stack[6][14] ),
    .A1(_0738_),
    .S(_0702_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_1 _4257_ (.A(_0739_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _4258_ (.A(_3163_),
    .B(_3186_),
    .Y(_0740_));
 sky130_fd_sc_hd__or2_2 _4259_ (.A(_3056_),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__or4_1 _4260_ (.A(\as2650.ins_reg[3] ),
    .B(_3078_),
    .C(_3222_),
    .D(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__or3_1 _4261_ (.A(_3079_),
    .B(_3207_),
    .C(_0741_),
    .X(_0743_));
 sky130_fd_sc_hd__buf_2 _4262_ (.A(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__or2_1 _4263_ (.A(_3200_),
    .B(_0741_),
    .X(_0745_));
 sky130_fd_sc_hd__or4_4 _4264_ (.A(_3090_),
    .B(_3209_),
    .C(_3212_),
    .D(_0740_),
    .X(_0746_));
 sky130_fd_sc_hd__nor2_1 _4265_ (.A(_3055_),
    .B(_0740_),
    .Y(_0747_));
 sky130_fd_sc_hd__and3_2 _4266_ (.A(_3102_),
    .B(_0356_),
    .C(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__inv_2 _4267_ (.A(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__or2_2 _4268_ (.A(_3184_),
    .B(_3055_),
    .X(_0750_));
 sky130_fd_sc_hd__or2_1 _4269_ (.A(_3327_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__or3_1 _4270_ (.A(_3214_),
    .B(_3217_),
    .C(_0740_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _4271_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__and4_1 _4272_ (.A(_0746_),
    .B(_0749_),
    .C(_0751_),
    .D(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__o311a_1 _4273_ (.A1(_3226_),
    .A2(_3228_),
    .A3(_0741_),
    .B1(_0745_),
    .C1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__and3_1 _4274_ (.A(_0742_),
    .B(_0744_),
    .C(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__or2_1 _4275_ (.A(_3071_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_2 _4276_ (.A(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__clkinv_2 _4277_ (.A(\as2650.halted ),
    .Y(_0759_));
 sky130_fd_sc_hd__clkbuf_4 _4278_ (.A(_3181_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_2 _4279_ (.A(_3174_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(_3184_),
    .B(_3160_),
    .Y(_0762_));
 sky130_fd_sc_hd__a31o_1 _4281_ (.A1(_0759_),
    .A2(_0761_),
    .A3(_0762_),
    .B1(net9),
    .X(_0763_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__and2_1 _4283_ (.A(_0758_),
    .B(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_2 _4284_ (.A(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_4 _4285_ (.A(_3080_),
    .X(_0767_));
 sky130_fd_sc_hd__or3_4 _4286_ (.A(_0767_),
    .B(_3331_),
    .C(_0750_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_4 _4287_ (.A(_0759_),
    .X(_0769_));
 sky130_fd_sc_hd__and4_1 _4288_ (.A(_0769_),
    .B(_3153_),
    .C(_0761_),
    .D(_0762_),
    .X(_0770_));
 sky130_fd_sc_hd__o221a_1 _4289_ (.A1(_3262_),
    .A2(_0314_),
    .B1(_3360_),
    .B2(_0768_),
    .C1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__clkbuf_4 _4290_ (.A(_0751_),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_1 _4291_ (.A(_3184_),
    .B(_3167_),
    .Y(_0773_));
 sky130_fd_sc_hd__and4_2 _4292_ (.A(_3252_),
    .B(_3215_),
    .C(_3254_),
    .D(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__and3_2 _4293_ (.A(_3299_),
    .B(_3301_),
    .C(_0773_),
    .X(_0775_));
 sky130_fd_sc_hd__or2_2 _4294_ (.A(_3223_),
    .B(_0741_),
    .X(_0776_));
 sky130_fd_sc_hd__clkbuf_4 _4295_ (.A(_3192_),
    .X(_0777_));
 sky130_fd_sc_hd__or3_2 _4296_ (.A(_0777_),
    .B(_3193_),
    .C(_0741_),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_1 _4297_ (.A(_3200_),
    .B(_0741_),
    .Y(_0779_));
 sky130_fd_sc_hd__buf_2 _4298_ (.A(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__nor2_2 _4299_ (.A(_3223_),
    .B(_0741_),
    .Y(_0781_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(_3288_),
    .B(_0779_),
    .Y(_0782_));
 sky130_fd_sc_hd__a211o_1 _4301_ (.A1(_3028_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__o211a_1 _4302_ (.A1(_3280_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__and3_2 _4303_ (.A(_0690_),
    .B(_3294_),
    .C(_0747_),
    .X(_0785_));
 sky130_fd_sc_hd__a211o_1 _4304_ (.A1(_3273_),
    .A2(_0748_),
    .B1(_0784_),
    .C1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__o211a_1 _4305_ (.A1(_3262_),
    .A2(_0744_),
    .B1(_0786_),
    .C1(_0746_),
    .X(_0787_));
 sky130_fd_sc_hd__a211o_1 _4306_ (.A1(_3260_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__o21ai_1 _4307_ (.A1(_3250_),
    .A2(_0753_),
    .B1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nor2_1 _4308_ (.A(_3325_),
    .B(_0772_),
    .Y(_0790_));
 sky130_fd_sc_hd__a21o_1 _4309_ (.A1(_0772_),
    .A2(_0789_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _4310_ (.A(_0758_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__a211o_1 _4311_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_0766_),
    .B1(_0771_),
    .C1(_0792_),
    .X(_0031_));
 sky130_fd_sc_hd__inv_2 _4312_ (.A(_0751_),
    .Y(_0793_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_3128_),
    .A1(_3401_),
    .S(_0745_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(_3397_),
    .A1(_0794_),
    .S(_0742_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(_3287_),
    .A1(_0795_),
    .S(_0749_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(_3391_),
    .A1(_0796_),
    .S(_0744_),
    .X(_0797_));
 sky130_fd_sc_hd__a21o_1 _4317_ (.A1(_0303_),
    .A2(_0774_),
    .B1(_0775_),
    .X(_0798_));
 sky130_fd_sc_hd__a21o_1 _4318_ (.A1(_0746_),
    .A2(_0797_),
    .B1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__o21a_1 _4319_ (.A1(_0307_),
    .A2(_0753_),
    .B1(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__or2_1 _4320_ (.A(_3389_),
    .B(_0751_),
    .X(_0801_));
 sky130_fd_sc_hd__o21ai_2 _4321_ (.A1(_0793_),
    .A2(_0800_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(_0758_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _4323_ (.A(_3163_),
    .B(_0690_),
    .Y(_0804_));
 sky130_fd_sc_hd__and4b_2 _4324_ (.A_N(_0804_),
    .B(_0761_),
    .C(_3153_),
    .D(_0769_),
    .X(_0805_));
 sky130_fd_sc_hd__o221a_1 _4325_ (.A1(_0659_),
    .A2(_0314_),
    .B1(_0322_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__a211o_1 _4326_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_0766_),
    .B1(_0803_),
    .C1(_0806_),
    .X(_0032_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(_0345_),
    .B(_0780_),
    .Y(_0807_));
 sky130_fd_sc_hd__a211o_1 _4328_ (.A1(_3131_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__o211a_1 _4329_ (.A1(_0354_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a211o_1 _4330_ (.A1(_3280_),
    .A2(_0748_),
    .B1(_0809_),
    .C1(_0785_),
    .X(_0810_));
 sky130_fd_sc_hd__o211a_1 _4331_ (.A1(_0326_),
    .A2(_0744_),
    .B1(_0810_),
    .C1(_0746_),
    .X(_0811_));
 sky130_fd_sc_hd__a211o_1 _4332_ (.A1(_0342_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__o21ai_1 _4333_ (.A1(_0340_),
    .A2(_0753_),
    .B1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__nor2_1 _4334_ (.A(_0377_),
    .B(_0772_),
    .Y(_0814_));
 sky130_fd_sc_hd__a21o_2 _4335_ (.A1(_0772_),
    .A2(_0813_),
    .B1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _4336_ (.A(_0758_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__o221a_1 _4337_ (.A1(_0664_),
    .A2(_0314_),
    .B1(_0332_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0817_));
 sky130_fd_sc_hd__a211o_1 _4338_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_0766_),
    .B1(_0816_),
    .C1(_0817_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_4 _4339_ (.A(net4),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _4340_ (.A(_0406_),
    .B(_0780_),
    .Y(_0819_));
 sky130_fd_sc_hd__a211o_1 _4341_ (.A1(_0818_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__o211a_1 _4342_ (.A1(_0414_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__nor2_1 _4343_ (.A(_3397_),
    .B(_0778_),
    .Y(_0822_));
 sky130_fd_sc_hd__o21ai_1 _4344_ (.A1(_0821_),
    .A2(_0822_),
    .B1(_0744_),
    .Y(_0823_));
 sky130_fd_sc_hd__o211a_1 _4345_ (.A1(_0417_),
    .A2(_0744_),
    .B1(_0823_),
    .C1(_0746_),
    .X(_0824_));
 sky130_fd_sc_hd__a211o_1 _4346_ (.A1(_0420_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__o21ai_1 _4347_ (.A1(_0403_),
    .A2(_0753_),
    .B1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__mux2_2 _4348_ (.A0(_0397_),
    .A1(_0826_),
    .S(_0772_),
    .X(_0827_));
 sky130_fd_sc_hd__nor2_1 _4349_ (.A(_0758_),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__o221a_1 _4350_ (.A1(_0667_),
    .A2(_0314_),
    .B1(_0431_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0829_));
 sky130_fd_sc_hd__a211o_1 _4351_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_0766_),
    .B1(_0828_),
    .C1(_0829_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(_3137_),
    .A1(_0463_),
    .S(_0745_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(_0461_),
    .A1(_0830_),
    .S(_0742_),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(_0354_),
    .A1(_0831_),
    .S(_0749_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _4355_ (.A(_0785_),
    .B(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__o211a_1 _4356_ (.A1(_0470_),
    .A2(_0744_),
    .B1(_0833_),
    .C1(_0746_),
    .X(_0834_));
 sky130_fd_sc_hd__a211o_1 _4357_ (.A1(_0477_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _4358_ (.A(_0480_),
    .B(_0753_),
    .X(_0836_));
 sky130_fd_sc_hd__a21o_1 _4359_ (.A1(_0835_),
    .A2(_0836_),
    .B1(_0793_),
    .X(_0837_));
 sky130_fd_sc_hd__o21ai_4 _4360_ (.A1(_0454_),
    .A2(_0772_),
    .B1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _4361_ (.A(_0758_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__o221a_1 _4362_ (.A1(_0470_),
    .A2(_0314_),
    .B1(_0488_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0840_));
 sky130_fd_sc_hd__a211o_1 _4363_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_0766_),
    .B1(_0839_),
    .C1(_0840_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _4364_ (.A(_0507_),
    .B(_0780_),
    .Y(_0841_));
 sky130_fd_sc_hd__a211o_1 _4365_ (.A1(_3140_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__o211a_1 _4366_ (.A1(_0566_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__a211o_1 _4367_ (.A1(_0439_),
    .A2(_0748_),
    .B1(_0843_),
    .C1(_0785_),
    .X(_0844_));
 sky130_fd_sc_hd__o211a_1 _4368_ (.A1(_0513_),
    .A2(_0744_),
    .B1(_0844_),
    .C1(_0746_),
    .X(_0845_));
 sky130_fd_sc_hd__a211o_1 _4369_ (.A1(_0516_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__o21ai_1 _4370_ (.A1(_0499_),
    .A2(_0753_),
    .B1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _4371_ (.A(_0535_),
    .B(_0772_),
    .Y(_0848_));
 sky130_fd_sc_hd__a21o_2 _4372_ (.A1(_0772_),
    .A2(_0847_),
    .B1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__nor2_1 _4373_ (.A(_0758_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__o221a_1 _4374_ (.A1(_0513_),
    .A2(_0314_),
    .B1(_0541_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0851_));
 sky130_fd_sc_hd__a211o_1 _4375_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_0766_),
    .B1(_0850_),
    .C1(_0851_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(_0584_),
    .B(_0780_),
    .Y(_0852_));
 sky130_fd_sc_hd__a211o_1 _4377_ (.A1(_3143_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__o211a_1 _4378_ (.A1(_3271_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__a211o_1 _4379_ (.A1(_0461_),
    .A2(_0748_),
    .B1(_0854_),
    .C1(_0785_),
    .X(_0855_));
 sky130_fd_sc_hd__o211a_1 _4380_ (.A1(_0545_),
    .A2(_0744_),
    .B1(_0855_),
    .C1(_0746_),
    .X(_0856_));
 sky130_fd_sc_hd__a211o_1 _4381_ (.A1(_0579_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__o21ai_1 _4382_ (.A1(_0577_),
    .A2(_0753_),
    .B1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(_0571_),
    .A1(_0858_),
    .S(_0772_),
    .X(_0859_));
 sky130_fd_sc_hd__nor2_1 _4384_ (.A(_0758_),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__o221a_1 _4385_ (.A1(_0545_),
    .A2(_0314_),
    .B1(_0550_),
    .B2(_0768_),
    .C1(_0805_),
    .X(_0861_));
 sky130_fd_sc_hd__a211o_1 _4386_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_0766_),
    .B1(_0860_),
    .C1(_0861_),
    .X(_0037_));
 sky130_fd_sc_hd__nor2_1 _4387_ (.A(_0621_),
    .B(_0779_),
    .Y(_0862_));
 sky130_fd_sc_hd__a211o_1 _4388_ (.A1(_3147_),
    .A2(_0780_),
    .B1(_0781_),
    .C1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__o211a_1 _4389_ (.A1(_0619_),
    .A2(_0776_),
    .B1(_0778_),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__a211o_1 _4390_ (.A1(_0566_),
    .A2(_0748_),
    .B1(_0864_),
    .C1(_0785_),
    .X(_0865_));
 sky130_fd_sc_hd__inv_2 _4391_ (.A(_0618_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(_0866_),
    .B(_0785_),
    .Y(_0867_));
 sky130_fd_sc_hd__a21o_1 _4393_ (.A1(_0865_),
    .A2(_0867_),
    .B1(_0774_),
    .X(_0868_));
 sky130_fd_sc_hd__o211a_1 _4394_ (.A1(_0628_),
    .A2(_0746_),
    .B1(_0753_),
    .C1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a211o_1 _4395_ (.A1(_0616_),
    .A2(_0775_),
    .B1(_0869_),
    .C1(_0793_),
    .X(_0870_));
 sky130_fd_sc_hd__o21a_1 _4396_ (.A1(_0611_),
    .A2(_0772_),
    .B1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__a32o_1 _4397_ (.A1(_0618_),
    .A2(_0768_),
    .A3(_0805_),
    .B1(_0764_),
    .B2(\as2650.r123_2[0][7] ),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(_0871_),
    .A1(_0872_),
    .S(_0758_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_1 _4399_ (.A(_0873_),
    .X(_0038_));
 sky130_fd_sc_hd__nand3_4 _4400_ (.A(_3065_),
    .B(_3039_),
    .C(_3170_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_2 _4401_ (.A(_3197_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _4402_ (.A(_3222_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_0876_),
    .B(_3192_),
    .Y(_0877_));
 sky130_fd_sc_hd__buf_2 _4404_ (.A(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__nand2_2 _4405_ (.A(_3182_),
    .B(_3363_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_3071_),
    .B(_3202_),
    .Y(_0880_));
 sky130_fd_sc_hd__nor2_2 _4407_ (.A(_3173_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__or2_1 _4408_ (.A(_0653_),
    .B(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__or2_1 _4409_ (.A(_3178_),
    .B(_0880_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_1 _4410_ (.A(_3177_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_1 _4411_ (.A(_0882_),
    .B(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__or3b_1 _4412_ (.A(_3159_),
    .B(_0879_),
    .C_N(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__buf_4 _4413_ (.A(_3121_),
    .X(_0887_));
 sky130_fd_sc_hd__buf_4 _4414_ (.A(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__buf_4 _4415_ (.A(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_4 _4416_ (.A(\as2650.halted ),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_4 _4417_ (.A(_3119_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_4 _4418_ (.A(_3051_),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _4419_ (.A(_3065_),
    .B(_3104_),
    .X(_0893_));
 sky130_fd_sc_hd__or3b_1 _4420_ (.A(_3318_),
    .B(_3196_),
    .C_N(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__buf_2 _4421_ (.A(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nor2_2 _4422_ (.A(_3180_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__nor2_4 _4423_ (.A(_3040_),
    .B(_3045_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_4 _4424_ (.A(_3104_),
    .B(_3039_),
    .Y(_0898_));
 sky130_fd_sc_hd__or2_2 _4425_ (.A(_0897_),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__nor2_2 _4426_ (.A(_3065_),
    .B(_3196_),
    .Y(_0900_));
 sky130_fd_sc_hd__a2111o_1 _4427_ (.A1(_0892_),
    .A2(_0896_),
    .B1(_0899_),
    .C1(_0878_),
    .D1(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_4 _4428_ (.A(_3083_),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _4429_ (.A(_3109_),
    .B(_0895_),
    .Y(_0903_));
 sky130_fd_sc_hd__or4_1 _4430_ (.A(_0902_),
    .B(_0875_),
    .C(_0877_),
    .D(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__or4b_1 _4431_ (.A(_0890_),
    .B(_0891_),
    .C(_0901_),
    .D_N(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a2111oi_1 _4432_ (.A1(_0889_),
    .A2(_0881_),
    .B1(_0905_),
    .C1(_0879_),
    .D1(_0653_),
    .Y(_0906_));
 sky130_fd_sc_hd__buf_4 _4433_ (.A(_0690_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_4 _4434_ (.A(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _4435_ (.A(\as2650.psl[6] ),
    .B(_3178_),
    .Y(_0909_));
 sky130_fd_sc_hd__or2_1 _4436_ (.A(\as2650.psl[6] ),
    .B(_3178_),
    .X(_0910_));
 sky130_fd_sc_hd__xor2_1 _4437_ (.A(\as2650.psl[7] ),
    .B(_3071_),
    .X(_0911_));
 sky130_fd_sc_hd__a21oi_1 _4438_ (.A1(_0909_),
    .A2(_0910_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2_2 _4439_ (.A(_3109_),
    .B(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__a31o_1 _4440_ (.A1(_3323_),
    .A2(_0908_),
    .A3(_0913_),
    .B1(_0874_),
    .X(_0914_));
 sky130_fd_sc_hd__o311a_1 _4441_ (.A1(_0875_),
    .A2(_0878_),
    .A3(_0886_),
    .B1(_0906_),
    .C1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__or2_2 _4442_ (.A(_3186_),
    .B(_0895_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(\as2650.psu[5] ),
    .A1(_0916_),
    .S(_3140_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(_0513_),
    .A1(_0917_),
    .S(_0767_),
    .X(_0918_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(_0874_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__buf_2 _4446_ (.A(net9),
    .X(_0920_));
 sky130_fd_sc_hd__buf_6 _4447_ (.A(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a21oi_1 _4448_ (.A1(_0915_),
    .A2(_0919_),
    .B1(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__o21a_1 _4449_ (.A1(\as2650.psu[5] ),
    .A2(_0915_),
    .B1(_0922_),
    .X(_0039_));
 sky130_fd_sc_hd__or3_4 _4450_ (.A(_0700_),
    .B(_3352_),
    .C(_0725_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_4 _4451_ (.A(_0651_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(\as2650.stack[5][8] ),
    .A1(_0699_),
    .S(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _4453_ (.A(_0925_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(\as2650.stack[5][9] ),
    .A1(_0709_),
    .S(_0924_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _4455_ (.A(_0926_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4456_ (.A0(\as2650.stack[5][10] ),
    .A1(_0715_),
    .S(_0924_),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _4457_ (.A(_0927_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(\as2650.stack[5][11] ),
    .A1(_0721_),
    .S(_0924_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _4459_ (.A(_0928_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4460_ (.A0(\as2650.stack[5][12] ),
    .A1(_0728_),
    .S(_0924_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_1 _4461_ (.A(_0929_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(\as2650.stack[5][13] ),
    .A1(_0733_),
    .S(_0924_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _4463_ (.A(_0930_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(\as2650.stack[5][14] ),
    .A1(_0738_),
    .S(_0924_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _4465_ (.A(_0931_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_4 _4466_ (.A(_0649_),
    .X(_0932_));
 sky130_fd_sc_hd__or2_4 _4467_ (.A(_3336_),
    .B(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__or2_4 _4468_ (.A(_3336_),
    .B(_0725_),
    .X(_0934_));
 sky130_fd_sc_hd__nand2_4 _4469_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(\as2650.stack[4][8] ),
    .A1(_0699_),
    .S(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _4471_ (.A(_0936_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(\as2650.stack[4][9] ),
    .A1(_0709_),
    .S(_0935_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_1 _4473_ (.A(_0937_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(\as2650.stack[4][10] ),
    .A1(_0715_),
    .S(_0935_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_1 _4475_ (.A(_0938_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(\as2650.stack[4][11] ),
    .A1(_0721_),
    .S(_0935_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_1 _4477_ (.A(_0939_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(\as2650.stack[4][12] ),
    .A1(_0728_),
    .S(_0935_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _4479_ (.A(_0940_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(\as2650.stack[4][13] ),
    .A1(_0733_),
    .S(_0935_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_1 _4481_ (.A(_0941_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(\as2650.stack[4][14] ),
    .A1(_0738_),
    .S(_0935_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_1 _4483_ (.A(_0942_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _4484_ (.A(_0557_),
    .B(_0603_),
    .Y(_0943_));
 sky130_fd_sc_hd__or2_1 _4485_ (.A(_0364_),
    .B(_0383_),
    .X(_0944_));
 sky130_fd_sc_hd__or4_1 _4486_ (.A(_0887_),
    .B(_3371_),
    .C(_0441_),
    .D(_0522_),
    .X(_0945_));
 sky130_fd_sc_hd__inv_2 _4487_ (.A(\as2650.psl[1] ),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _4488_ (.A(_0946_),
    .B(_0598_),
    .Y(_0947_));
 sky130_fd_sc_hd__a21bo_1 _4489_ (.A1(_0603_),
    .A2(_0599_),
    .B1_N(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__and2_1 _4490_ (.A(_3306_),
    .B(_3308_),
    .X(_0949_));
 sky130_fd_sc_hd__o22a_1 _4491_ (.A1(_0949_),
    .A2(_3371_),
    .B1(_3387_),
    .B2(_3369_),
    .X(_0950_));
 sky130_fd_sc_hd__or3_1 _4492_ (.A(_0363_),
    .B(_0371_),
    .C(_0383_),
    .X(_0951_));
 sky130_fd_sc_hd__o211a_1 _4493_ (.A1(_0950_),
    .A2(_0944_),
    .B1(_0951_),
    .C1(_0445_),
    .X(_0952_));
 sky130_fd_sc_hd__o21a_1 _4494_ (.A1(_0441_),
    .A2(_0952_),
    .B1(_0525_),
    .X(_0953_));
 sky130_fd_sc_hd__o21a_1 _4495_ (.A1(_0522_),
    .A2(_0953_),
    .B1(_0559_),
    .X(_0954_));
 sky130_fd_sc_hd__o2bb2a_1 _4496_ (.A1_N(_0597_),
    .A2_N(_0606_),
    .B1(_0943_),
    .B2(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(_0947_),
    .A1(_0948_),
    .S(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a21o_1 _4498_ (.A1(_3229_),
    .A2(_0956_),
    .B1(_0888_),
    .X(_0957_));
 sky130_fd_sc_hd__o41a_1 _4499_ (.A1(_3310_),
    .A2(_0943_),
    .A3(_0944_),
    .A4(_0945_),
    .B1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__or4_1 _4500_ (.A(_3325_),
    .B(_3389_),
    .C(_0377_),
    .D(_0454_),
    .X(_0959_));
 sky130_fd_sc_hd__nor2_1 _4501_ (.A(_0535_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__a31o_1 _4502_ (.A1(_0397_),
    .A2(_0571_),
    .A3(_0960_),
    .B1(_0611_),
    .X(_0961_));
 sky130_fd_sc_hd__nor2_1 _4503_ (.A(_3229_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__and3_2 _4504_ (.A(_3049_),
    .B(_3189_),
    .C(_3170_),
    .X(_0963_));
 sky130_fd_sc_hd__or4_1 _4505_ (.A(_0544_),
    .B(_0513_),
    .C(_0470_),
    .D(_0417_),
    .X(_0964_));
 sky130_fd_sc_hd__or4_1 _4506_ (.A(_0326_),
    .B(_3391_),
    .C(_3262_),
    .D(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_0866_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__nor2_1 _4508_ (.A(_0963_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__a311o_1 _4509_ (.A1(_0596_),
    .A2(_0613_),
    .A3(_0963_),
    .B1(_0967_),
    .C1(_0767_),
    .X(_0968_));
 sky130_fd_sc_hd__buf_4 _4510_ (.A(_3049_),
    .X(_0969_));
 sky130_fd_sc_hd__buf_4 _4511_ (.A(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__o211a_1 _4512_ (.A1(_0958_),
    .A2(_0962_),
    .B1(_0968_),
    .C1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__buf_4 _4513_ (.A(_3104_),
    .X(_0972_));
 sky130_fd_sc_hd__clkbuf_4 _4514_ (.A(_0902_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _4515_ (.A(_3293_),
    .B(_3169_),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_2 _4516_ (.A(_3101_),
    .B(_3158_),
    .Y(_0975_));
 sky130_fd_sc_hd__a22o_1 _4517_ (.A1(_3121_),
    .A2(_0974_),
    .B1(_0975_),
    .B2(_3292_),
    .X(_0976_));
 sky130_fd_sc_hd__a31o_1 _4518_ (.A1(_0972_),
    .A2(_0973_),
    .A3(_3198_),
    .B1(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__nand2_1 _4519_ (.A(_0690_),
    .B(_0884_),
    .Y(_0978_));
 sky130_fd_sc_hd__or3b_1 _4520_ (.A(_0879_),
    .B(_0653_),
    .C_N(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__nor2_1 _4521_ (.A(_3227_),
    .B(_0969_),
    .Y(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _4522_ (.A(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__and3b_1 _4523_ (.A_N(_0904_),
    .B(_3189_),
    .C(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__clkbuf_4 _4524_ (.A(_3101_),
    .X(_0983_));
 sky130_fd_sc_hd__and3b_1 _4525_ (.A_N(\as2650.ins_reg[2] ),
    .B(_3038_),
    .C(_3319_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_2 _4526_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__nor2_2 _4527_ (.A(_3065_),
    .B(_3191_),
    .Y(_0986_));
 sky130_fd_sc_hd__nor2_1 _4528_ (.A(_0985_),
    .B(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__clkbuf_4 _4529_ (.A(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__and3_1 _4530_ (.A(_3065_),
    .B(_3038_),
    .C(_3170_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_4 _4531_ (.A(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_4 _4532_ (.A(_3227_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__and4_1 _4533_ (.A(_3119_),
    .B(_3197_),
    .C(_0988_),
    .D(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__or4_1 _4534_ (.A(_3158_),
    .B(_0900_),
    .C(_0990_),
    .D(_0877_),
    .X(_0993_));
 sky130_fd_sc_hd__or4bb_1 _4535_ (.A(_0898_),
    .B(_3170_),
    .C_N(_3181_),
    .D_N(_3363_),
    .X(_0994_));
 sky130_fd_sc_hd__nor2_1 _4536_ (.A(_0993_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__or3_1 _4537_ (.A(_0879_),
    .B(_0882_),
    .C(_0884_),
    .X(_0996_));
 sky130_fd_sc_hd__nor3_1 _4538_ (.A(_3073_),
    .B(_3292_),
    .C(_3177_),
    .Y(_0997_));
 sky130_fd_sc_hd__nor2_1 _4539_ (.A(_0996_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__a22oi_1 _4540_ (.A1(_0983_),
    .A2(_0992_),
    .B1(_0995_),
    .B2(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_2 _4541_ (.A(_3068_),
    .B(_0900_),
    .Y(_1000_));
 sky130_fd_sc_hd__or2_1 _4542_ (.A(\as2650.ins_reg[3] ),
    .B(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__o31a_1 _4543_ (.A1(_3227_),
    .A2(_3102_),
    .A3(_0988_),
    .B1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__nand2_4 _4544_ (.A(_3104_),
    .B(_0989_),
    .Y(_1003_));
 sky130_fd_sc_hd__nor2_1 _4545_ (.A(\as2650.halted ),
    .B(_3037_),
    .Y(_1004_));
 sky130_fd_sc_hd__or3_1 _4546_ (.A(_3038_),
    .B(_3221_),
    .C(_3169_),
    .X(_1005_));
 sky130_fd_sc_hd__or2_1 _4547_ (.A(_3079_),
    .B(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__and3_1 _4548_ (.A(_1003_),
    .B(_1004_),
    .C(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_2 _4549_ (.A(_3032_),
    .B(_3057_),
    .Y(_1008_));
 sky130_fd_sc_hd__or3_1 _4550_ (.A(_3101_),
    .B(_1008_),
    .C(_3156_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_4 _4551_ (.A(_3178_),
    .X(_1010_));
 sky130_fd_sc_hd__or3_2 _4552_ (.A(_1010_),
    .B(_0902_),
    .C(_0895_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_3102_),
    .B(_1005_),
    .Y(_1012_));
 sky130_fd_sc_hd__or4_1 _4554_ (.A(_3101_),
    .B(_3294_),
    .C(_0963_),
    .D(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__and4b_1 _4555_ (.A_N(_3053_),
    .B(_1009_),
    .C(_1011_),
    .D(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__and3_1 _4556_ (.A(_3066_),
    .B(_1007_),
    .C(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and3_1 _4557_ (.A(_0999_),
    .B(_1002_),
    .C(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__or4b_2 _4558_ (.A(_0977_),
    .B(_0979_),
    .C(_0982_),
    .D_N(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_4 _4559_ (.A(_0983_),
    .X(_1018_));
 sky130_fd_sc_hd__buf_2 _4560_ (.A(_3198_),
    .X(_1019_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_3149_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _4562_ (.A(_1018_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__clkinv_4 _4563_ (.A(_3142_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_1022_),
    .B(_1019_),
    .Y(_1023_));
 sky130_fd_sc_hd__or4_1 _4565_ (.A(_3132_),
    .B(_3135_),
    .C(_3137_),
    .D(_3140_),
    .X(_1024_));
 sky130_fd_sc_hd__or4_1 _4566_ (.A(_3029_),
    .B(_3129_),
    .C(_1023_),
    .D(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__inv_2 _4567_ (.A(_3273_),
    .Y(_1026_));
 sky130_fd_sc_hd__a211o_1 _4568_ (.A1(_1026_),
    .A2(_0492_),
    .B1(_0566_),
    .C1(_0777_),
    .X(_1027_));
 sky130_fd_sc_hd__inv_2 _4569_ (.A(_3178_),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_2 _4570_ (.A(\as2650.psl[6] ),
    .Y(_1029_));
 sky130_fd_sc_hd__mux2_1 _4571_ (.A0(_1029_),
    .A1(_3179_),
    .S(_3144_),
    .X(_1030_));
 sky130_fd_sc_hd__a21oi_1 _4572_ (.A1(_0881_),
    .A2(_0966_),
    .B1(_3160_),
    .Y(_1031_));
 sky130_fd_sc_hd__o21ai_1 _4573_ (.A1(_0545_),
    .A2(_0881_),
    .B1(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__o41a_1 _4574_ (.A1(_1028_),
    .A2(_0887_),
    .A3(_0895_),
    .A4(_1030_),
    .B1(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__or2_1 _4575_ (.A(_3397_),
    .B(_0354_),
    .X(_1034_));
 sky130_fd_sc_hd__or4b_1 _4576_ (.A(_3280_),
    .B(_3271_),
    .C(_1034_),
    .D_N(_0582_),
    .X(_1035_));
 sky130_fd_sc_hd__or3b_1 _4577_ (.A(_0876_),
    .B(_0619_),
    .C_N(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or2_2 _4578_ (.A(_3068_),
    .B(_3197_),
    .X(_1037_));
 sky130_fd_sc_hd__o211a_1 _4579_ (.A1(_0878_),
    .A2(_1033_),
    .B1(_1036_),
    .C1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_1027_),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__and3b_1 _4581_ (.A_N(_1021_),
    .B(_1025_),
    .C(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__a21oi_1 _4582_ (.A1(_1029_),
    .A2(_1017_),
    .B1(_0921_),
    .Y(_1041_));
 sky130_fd_sc_hd__o31a_1 _4583_ (.A1(_0971_),
    .A2(_1017_),
    .A3(_1040_),
    .B1(_1041_),
    .X(_0054_));
 sky130_fd_sc_hd__inv_2 _4584_ (.A(\as2650.psl[7] ),
    .Y(_1042_));
 sky130_fd_sc_hd__o221a_1 _4585_ (.A1(_0777_),
    .A2(_0566_),
    .B1(_0619_),
    .B2(_0876_),
    .C1(_1037_),
    .X(_1043_));
 sky130_fd_sc_hd__or2_2 _4586_ (.A(_3180_),
    .B(_0894_),
    .X(_1044_));
 sky130_fd_sc_hd__and4_1 _4587_ (.A(_3039_),
    .B(_3323_),
    .C(_3107_),
    .D(_0893_),
    .X(_1045_));
 sky130_fd_sc_hd__inv_2 _4588_ (.A(_3139_),
    .Y(_1046_));
 sky130_fd_sc_hd__clkinv_2 _4589_ (.A(_3128_),
    .Y(_1047_));
 sky130_fd_sc_hd__o22a_1 _4590_ (.A1(\as2650.psl[1] ),
    .A2(_1047_),
    .B1(_1022_),
    .B2(\as2650.psl[6] ),
    .X(_1048_));
 sky130_fd_sc_hd__o221a_1 _4591_ (.A1(_3163_),
    .A2(_0465_),
    .B1(_1046_),
    .B2(\as2650.psl[5] ),
    .C1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _4592_ (.A(net8),
    .Y(_1050_));
 sky130_fd_sc_hd__clkinv_2 _4593_ (.A(_3131_),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _4594_ (.A(_3028_),
    .Y(_1052_));
 sky130_fd_sc_hd__o22a_1 _4595_ (.A1(\as2650.carry ),
    .A2(_1052_),
    .B1(_0818_),
    .B2(\as2650.psl[3] ),
    .X(_1053_));
 sky130_fd_sc_hd__o221a_1 _4596_ (.A1(\as2650.psl[7] ),
    .A2(_1050_),
    .B1(_1051_),
    .B2(\as2650.overflow ),
    .C1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__and4_1 _4597_ (.A(_1010_),
    .B(_1045_),
    .C(_1049_),
    .D(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _4598_ (.A(_3178_),
    .B(_1045_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_3028_),
    .B(_3244_),
    .Y(_1057_));
 sky130_fd_sc_hd__o221a_1 _4600_ (.A1(_0818_),
    .A2(_0354_),
    .B1(_0461_),
    .B2(_1046_),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__o22a_1 _4601_ (.A1(_1051_),
    .A2(_3396_),
    .B1(_0439_),
    .B2(_0465_),
    .X(_1059_));
 sky130_fd_sc_hd__o221a_1 _4602_ (.A1(_1047_),
    .A2(_3280_),
    .B1(_0566_),
    .B2(_1022_),
    .C1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__o2111a_1 _4603_ (.A1(_1050_),
    .A2(_3271_),
    .B1(_1056_),
    .C1(_1058_),
    .D1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__a211o_1 _4604_ (.A1(_1028_),
    .A2(_1045_),
    .B1(_1055_),
    .C1(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__o22a_1 _4605_ (.A1(\as2650.psu[0] ),
    .A2(_1052_),
    .B1(_1022_),
    .B2(io_out[26]),
    .X(_1063_));
 sky130_fd_sc_hd__o221a_1 _4606_ (.A1(\as2650.psu[3] ),
    .A2(_0818_),
    .B1(_0465_),
    .B2(\as2650.psu[4] ),
    .C1(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__o221a_1 _4607_ (.A1(\as2650.psu[7] ),
    .A2(_1050_),
    .B1(_1046_),
    .B2(\as2650.psu[5] ),
    .C1(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__o221a_1 _4608_ (.A1(_3343_),
    .A2(_1047_),
    .B1(_1051_),
    .B2(\as2650.psu[2] ),
    .C1(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__or3b_1 _4609_ (.A(_1010_),
    .B(_1066_),
    .C_N(_1045_),
    .X(_1067_));
 sky130_fd_sc_hd__o211a_1 _4610_ (.A1(_3073_),
    .A2(_0895_),
    .B1(_1062_),
    .C1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__or4_1 _4611_ (.A(\as2650.psl[7] ),
    .B(_3147_),
    .C(_3073_),
    .D(_0895_),
    .X(_1069_));
 sky130_fd_sc_hd__or3b_1 _4612_ (.A(_0896_),
    .B(_1068_),
    .C_N(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__o31a_1 _4613_ (.A1(_1042_),
    .A2(_3149_),
    .A3(_1044_),
    .B1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__nor2_1 _4614_ (.A(_0888_),
    .B(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a211o_1 _4615_ (.A1(_0618_),
    .A2(_0889_),
    .B1(_0878_),
    .C1(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a21o_1 _4616_ (.A1(_1043_),
    .A2(_1073_),
    .B1(_1021_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(_0618_),
    .A1(_3271_),
    .S(_0963_),
    .X(_1075_));
 sky130_fd_sc_hd__o21ba_1 _4618_ (.A1(_3229_),
    .A2(_0611_),
    .B1_N(_0957_),
    .X(_1076_));
 sky130_fd_sc_hd__a211o_1 _4619_ (.A1(_0908_),
    .A2(_1075_),
    .B1(_1076_),
    .C1(_1018_),
    .X(_1077_));
 sky130_fd_sc_hd__a21oi_1 _4620_ (.A1(_1074_),
    .A2(_1077_),
    .B1(_1017_),
    .Y(_1078_));
 sky130_fd_sc_hd__a211oi_1 _4621_ (.A1(_1042_),
    .A2(_1017_),
    .B1(_1078_),
    .C1(_0921_),
    .Y(_0055_));
 sky130_fd_sc_hd__or2_2 _4622_ (.A(\as2650.psu[2] ),
    .B(_3345_),
    .X(_1079_));
 sky130_fd_sc_hd__or2_4 _4623_ (.A(_0725_),
    .B(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__or2_4 _4624_ (.A(_0932_),
    .B(_1079_),
    .X(_1081_));
 sky130_fd_sc_hd__nand2_4 _4625_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__mux2_1 _4626_ (.A0(\as2650.stack[3][8] ),
    .A1(_0699_),
    .S(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_1 _4627_ (.A(_1083_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(\as2650.stack[3][9] ),
    .A1(_0709_),
    .S(_1082_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _4629_ (.A(_1084_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(\as2650.stack[3][10] ),
    .A1(_0715_),
    .S(_1082_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _4631_ (.A(_1085_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4632_ (.A0(\as2650.stack[3][11] ),
    .A1(_0721_),
    .S(_1082_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _4633_ (.A(_1086_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(\as2650.stack[3][12] ),
    .A1(_0728_),
    .S(_1082_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_1 _4635_ (.A(_1087_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4636_ (.A0(\as2650.stack[3][13] ),
    .A1(_0733_),
    .S(_1082_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _4637_ (.A(_1088_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(\as2650.stack[3][14] ),
    .A1(_0738_),
    .S(_1082_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_1 _4639_ (.A(_1089_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_4 _4640_ (.A(_1050_),
    .X(_1090_));
 sky130_fd_sc_hd__buf_4 _4641_ (.A(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__or2_1 _4642_ (.A(_3032_),
    .B(_3036_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_4 _4643_ (.A(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _4644_ (.A1(_1091_),
    .A2(_0892_),
    .B1(_3076_),
    .B2(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__or4_1 _4645_ (.A(_3155_),
    .B(_3045_),
    .C(_3056_),
    .D(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__buf_2 _4646_ (.A(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nor2_2 _4647_ (.A(_1093_),
    .B(_3056_),
    .Y(_1097_));
 sky130_fd_sc_hd__buf_4 _4648_ (.A(_3066_),
    .X(_1098_));
 sky130_fd_sc_hd__nor3_1 _4649_ (.A(_1098_),
    .B(_3037_),
    .C(_1096_),
    .Y(_1099_));
 sky130_fd_sc_hd__a221o_1 _4650_ (.A1(_1010_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_3029_),
    .C1(_1099_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4651_ (.A0(_3129_),
    .A1(_3123_),
    .S(_1093_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _4652_ (.A0(_1100_),
    .A1(_3071_),
    .S(_1096_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _4653_ (.A(_1101_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _4654_ (.A1(_3081_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_3132_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(_3323_),
    .A1(_3140_),
    .S(_1097_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _4656_ (.A(_1102_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _4657_ (.A1(_3067_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_3144_),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _4658_ (.A1(_3068_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_3150_),
    .X(_0068_));
 sky130_fd_sc_hd__or3_1 _4659_ (.A(_0317_),
    .B(_0329_),
    .C(_0649_),
    .X(_1103_));
 sky130_fd_sc_hd__buf_4 _4660_ (.A(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__or3_4 _4661_ (.A(_0317_),
    .B(_0329_),
    .C(_0725_),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_4 _4662_ (.A(_1104_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(\as2650.stack[2][8] ),
    .A1(_0699_),
    .S(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _4664_ (.A(_1107_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(\as2650.stack[2][9] ),
    .A1(_0709_),
    .S(_1106_),
    .X(_1108_));
 sky130_fd_sc_hd__clkbuf_1 _4666_ (.A(_1108_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(\as2650.stack[2][10] ),
    .A1(_0715_),
    .S(_1106_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _4668_ (.A(_1109_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(\as2650.stack[2][11] ),
    .A1(_0721_),
    .S(_1106_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _4670_ (.A(_1110_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4671_ (.A0(\as2650.stack[2][12] ),
    .A1(_0728_),
    .S(_1106_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _4672_ (.A(_1111_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(\as2650.stack[2][13] ),
    .A1(_0733_),
    .S(_1106_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _4674_ (.A(_1112_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(\as2650.stack[2][14] ),
    .A1(_0738_),
    .S(_1106_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _4676_ (.A(_1113_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_2 _4677_ (.A(_1010_),
    .B(_0756_),
    .X(_1114_));
 sky130_fd_sc_hd__inv_2 _4678_ (.A(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__o31ai_4 _4679_ (.A1(\as2650.halted ),
    .A2(_3363_),
    .A3(_0804_),
    .B1(_3153_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2_4 _4680_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor4b_4 _4681_ (.A(_3330_),
    .B(_0750_),
    .C(_1117_),
    .D_N(_0879_),
    .Y(_1118_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(_0791_),
    .B(_1114_),
    .Y(_1119_));
 sky130_fd_sc_hd__a31o_1 _4683_ (.A1(_0634_),
    .A2(_0696_),
    .A3(_1118_),
    .B1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a21o_1 _4684_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_1117_),
    .B1(_1120_),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_4 _4685_ (.A(_1118_),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(_3390_),
    .B(_0695_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_3262_),
    .B(_0707_),
    .Y(_1123_));
 sky130_fd_sc_hd__and4_1 _4688_ (.A(_3391_),
    .B(_3261_),
    .C(_0696_),
    .D(_0707_),
    .X(_1124_));
 sky130_fd_sc_hd__a21oi_1 _4689_ (.A1(_1122_),
    .A2(_1123_),
    .B1(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__a2bb2o_1 _4690_ (.A1_N(_0802_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][1] ),
    .X(_1126_));
 sky130_fd_sc_hd__a21o_1 _4691_ (.A1(_1121_),
    .A2(_1125_),
    .B1(_1126_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _4692_ (.A1(_0325_),
    .A2(_0695_),
    .B1(_0707_),
    .B2(_3391_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2_1 _4693_ (.A(_0325_),
    .B(_0706_),
    .Y(_1128_));
 sky130_fd_sc_hd__or2_1 _4694_ (.A(_1122_),
    .B(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__and4_1 _4695_ (.A(_3261_),
    .B(_0712_),
    .C(_1127_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__a22oi_1 _4696_ (.A1(_3261_),
    .A2(_0712_),
    .B1(_1127_),
    .B2(_1129_),
    .Y(_1131_));
 sky130_fd_sc_hd__nor2_1 _4697_ (.A(_1130_),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_1124_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__or2_1 _4699_ (.A(_1124_),
    .B(_1132_),
    .X(_1134_));
 sky130_fd_sc_hd__and2_1 _4700_ (.A(_1133_),
    .B(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__a2bb2o_1 _4701_ (.A1_N(_0815_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][2] ),
    .X(_1136_));
 sky130_fd_sc_hd__a21o_1 _4702_ (.A1(_1121_),
    .A2(_1135_),
    .B1(_1136_),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_1 _4703_ (.A(_1122_),
    .B(_1128_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_0417_),
    .B(_0695_),
    .Y(_1138_));
 sky130_fd_sc_hd__and4_1 _4705_ (.A(_0348_),
    .B(_0325_),
    .C(_0695_),
    .D(_0706_),
    .X(_1139_));
 sky130_fd_sc_hd__a21o_1 _4706_ (.A1(_1128_),
    .A2(_1138_),
    .B1(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__and4_1 _4707_ (.A(_3390_),
    .B(\as2650.r0[0] ),
    .C(_0711_),
    .D(_0717_),
    .X(_1141_));
 sky130_fd_sc_hd__a22oi_1 _4708_ (.A1(_3390_),
    .A2(_0712_),
    .B1(_0718_),
    .B2(_3261_),
    .Y(_1142_));
 sky130_fd_sc_hd__or2_1 _4709_ (.A(_1141_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__xor2_1 _4710_ (.A(_1140_),
    .B(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__o21ai_2 _4711_ (.A1(_1137_),
    .A2(_1130_),
    .B1(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__o31ai_1 _4712_ (.A1(_1137_),
    .A2(_1130_),
    .A3(_1144_),
    .B1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__xor2_1 _4713_ (.A(_1133_),
    .B(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__a2bb2o_1 _4714_ (.A1_N(_0827_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][3] ),
    .X(_1148_));
 sky130_fd_sc_hd__a21o_1 _4715_ (.A1(_1121_),
    .A2(_1147_),
    .B1(_1148_),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _4716_ (.A(_1133_),
    .B(_1146_),
    .X(_1149_));
 sky130_fd_sc_hd__a21oi_1 _4717_ (.A1(_0348_),
    .A2(_0706_),
    .B1(_1141_),
    .Y(_1150_));
 sky130_fd_sc_hd__and3_1 _4718_ (.A(_0348_),
    .B(_0706_),
    .C(_1141_),
    .X(_1151_));
 sky130_fd_sc_hd__nor2_1 _4719_ (.A(_1150_),
    .B(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(_0469_),
    .B(_0695_),
    .Y(_1153_));
 sky130_fd_sc_hd__xor2_1 _4721_ (.A(_1152_),
    .B(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__nand2_1 _4722_ (.A(_0326_),
    .B(_0712_),
    .Y(_1155_));
 sky130_fd_sc_hd__and4_1 _4723_ (.A(\as2650.r0[1] ),
    .B(\as2650.r0[0] ),
    .C(_0717_),
    .D(_0723_),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _4724_ (.A1(\as2650.r0[1] ),
    .A2(_0717_),
    .B1(_0723_),
    .B2(\as2650.r0[0] ),
    .X(_1157_));
 sky130_fd_sc_hd__and2b_1 _4725_ (.A_N(_1156_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__xnor2_1 _4726_ (.A(_1155_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__xnor2_1 _4727_ (.A(_1154_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__o21bai_1 _4728_ (.A1(_1140_),
    .A2(_1143_),
    .B1_N(_1139_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__inv_2 _4730_ (.A(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_1 _4731_ (.A(_1160_),
    .B(_1161_),
    .Y(_1164_));
 sky130_fd_sc_hd__or2_1 _4732_ (.A(_1163_),
    .B(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_1 _4733_ (.A(_1149_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__and2_1 _4734_ (.A(_1149_),
    .B(_1165_),
    .X(_1167_));
 sky130_fd_sc_hd__or2_1 _4735_ (.A(_1166_),
    .B(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__nor2_1 _4736_ (.A(_1145_),
    .B(_1165_),
    .Y(_1169_));
 sky130_fd_sc_hd__a21oi_1 _4737_ (.A1(_1145_),
    .A2(_1168_),
    .B1(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__a2bb2o_1 _4738_ (.A1_N(_0838_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][4] ),
    .X(_1171_));
 sky130_fd_sc_hd__a21o_1 _4739_ (.A1(_1121_),
    .A2(_1170_),
    .B1(_1171_),
    .X(_0080_));
 sky130_fd_sc_hd__a31o_1 _4740_ (.A1(_0470_),
    .A2(_0696_),
    .A3(_1152_),
    .B1(_1151_),
    .X(_1172_));
 sky130_fd_sc_hd__or2b_1 _4741_ (.A(_1154_),
    .B_N(_1159_),
    .X(_1173_));
 sky130_fd_sc_hd__a22o_1 _4742_ (.A1(\as2650.r0[2] ),
    .A2(_0717_),
    .B1(_0723_),
    .B2(\as2650.r0[1] ),
    .X(_1174_));
 sky130_fd_sc_hd__nand4_1 _4743_ (.A(\as2650.r0[2] ),
    .B(_3390_),
    .C(_0717_),
    .D(_0723_),
    .Y(_1175_));
 sky130_fd_sc_hd__and2_1 _4744_ (.A(\as2650.r0[3] ),
    .B(_0711_),
    .X(_1176_));
 sky130_fd_sc_hd__a21o_1 _4745_ (.A1(_1174_),
    .A2(_1175_),
    .B1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__nand3_1 _4746_ (.A(_1176_),
    .B(_1174_),
    .C(_1175_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_3261_),
    .B(_0730_),
    .Y(_1179_));
 sky130_fd_sc_hd__inv_2 _4748_ (.A(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__and3_1 _4749_ (.A(_1177_),
    .B(_1178_),
    .C(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__a21oi_1 _4750_ (.A1(_1177_),
    .A2(_1178_),
    .B1(_1180_),
    .Y(_1182_));
 sky130_fd_sc_hd__or2_1 _4751_ (.A(_1181_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_0512_),
    .B(_0695_),
    .Y(_1184_));
 sky130_fd_sc_hd__a31o_1 _4753_ (.A1(_0325_),
    .A2(_0711_),
    .A3(_1157_),
    .B1(_1156_),
    .X(_1185_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_0469_),
    .B(_0706_),
    .Y(_1186_));
 sky130_fd_sc_hd__xnor2_1 _4755_ (.A(_1185_),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__xnor2_1 _4756_ (.A(_1184_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__xnor2_1 _4757_ (.A(_1183_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__xnor2_1 _4758_ (.A(_1173_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__xnor2_1 _4759_ (.A(_1172_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__a2111o_1 _4760_ (.A1(_1145_),
    .A2(_1149_),
    .B1(_1163_),
    .C1(_1164_),
    .D1(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__or2_1 _4761_ (.A(_1162_),
    .B(_1191_),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(_1162_),
    .B(_1191_),
    .Y(_1194_));
 sky130_fd_sc_hd__a211o_1 _4763_ (.A1(_1193_),
    .A2(_1194_),
    .B1(_1169_),
    .C1(_1166_),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _4764_ (.A(_1192_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__a2bb2o_1 _4765_ (.A1_N(_0849_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][5] ),
    .X(_1197_));
 sky130_fd_sc_hd__a21o_1 _4766_ (.A1(_1121_),
    .A2(_1196_),
    .B1(_1197_),
    .X(_0081_));
 sky130_fd_sc_hd__or2b_1 _4767_ (.A(_1173_),
    .B_N(_1189_),
    .X(_1198_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_1172_),
    .B(_1190_),
    .Y(_1199_));
 sky130_fd_sc_hd__and2b_1 _4769_ (.A_N(_1183_),
    .B(_1188_),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _4770_ (.A1(_0348_),
    .A2(_0718_),
    .B1(_0724_),
    .B2(_0325_),
    .X(_1201_));
 sky130_fd_sc_hd__nand4_1 _4771_ (.A(_0348_),
    .B(_0325_),
    .C(_0718_),
    .D(_0724_),
    .Y(_1202_));
 sky130_fd_sc_hd__and2_1 _4772_ (.A(_0469_),
    .B(_0711_),
    .X(_1203_));
 sky130_fd_sc_hd__a21o_1 _4773_ (.A1(_1201_),
    .A2(_1202_),
    .B1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__nand3_1 _4774_ (.A(_1201_),
    .B(_1202_),
    .C(_1203_),
    .Y(_1205_));
 sky130_fd_sc_hd__a22oi_1 _4775_ (.A1(_3390_),
    .A2(_0730_),
    .B1(_0736_),
    .B2(_3261_),
    .Y(_1206_));
 sky130_fd_sc_hd__and4_1 _4776_ (.A(_3390_),
    .B(_3261_),
    .C(_0730_),
    .D(_0735_),
    .X(_1207_));
 sky130_fd_sc_hd__nor2_1 _4777_ (.A(_1206_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__nand3_1 _4778_ (.A(_1204_),
    .B(_1205_),
    .C(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21o_1 _4779_ (.A1(_1204_),
    .A2(_1205_),
    .B1(_1208_),
    .X(_1210_));
 sky130_fd_sc_hd__nand3_2 _4780_ (.A(_1181_),
    .B(_1209_),
    .C(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__a21o_1 _4781_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1181_),
    .X(_1212_));
 sky130_fd_sc_hd__nand2_1 _4782_ (.A(_0544_),
    .B(_0695_),
    .Y(_1213_));
 sky130_fd_sc_hd__a21bo_1 _4783_ (.A1(_1176_),
    .A2(_1174_),
    .B1_N(_1175_),
    .X(_1214_));
 sky130_fd_sc_hd__nand2_1 _4784_ (.A(_0512_),
    .B(_0706_),
    .Y(_1215_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__xnor2_1 _4786_ (.A(_1213_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a21o_1 _4787_ (.A1(_1211_),
    .A2(_1212_),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__nand3_2 _4788_ (.A(_1211_),
    .B(_1212_),
    .C(_1217_),
    .Y(_1219_));
 sky130_fd_sc_hd__nand3_2 _4789_ (.A(_1200_),
    .B(_1218_),
    .C(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a21o_1 _4790_ (.A1(_1218_),
    .A2(_1219_),
    .B1(_1200_),
    .X(_1221_));
 sky130_fd_sc_hd__and3_1 _4791_ (.A(_0470_),
    .B(_0707_),
    .C(_1185_),
    .X(_1222_));
 sky130_fd_sc_hd__a31o_1 _4792_ (.A1(_0512_),
    .A2(_0696_),
    .A3(_1187_),
    .B1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a21oi_1 _4793_ (.A1(_1220_),
    .A2(_1221_),
    .B1(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__and3_1 _4794_ (.A(_1223_),
    .B(_1220_),
    .C(_1221_),
    .X(_1225_));
 sky130_fd_sc_hd__a211oi_2 _4795_ (.A1(_1198_),
    .A2(_1199_),
    .B1(_1224_),
    .C1(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__o211a_1 _4796_ (.A1(_1224_),
    .A2(_1225_),
    .B1(_1198_),
    .C1(_1199_),
    .X(_1227_));
 sky130_fd_sc_hd__a211oi_2 _4797_ (.A1(_1193_),
    .A2(_1192_),
    .B1(_1226_),
    .C1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__o211a_1 _4798_ (.A1(_1226_),
    .A2(_1227_),
    .B1(_1193_),
    .C1(_1192_),
    .X(_1229_));
 sky130_fd_sc_hd__nor2_1 _4799_ (.A(_1228_),
    .B(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__a2bb2o_1 _4800_ (.A1_N(_0859_),
    .A2_N(_1114_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][6] ),
    .X(_1231_));
 sky130_fd_sc_hd__a21o_1 _4801_ (.A1(_1121_),
    .A2(_1230_),
    .B1(_1231_),
    .X(_0082_));
 sky130_fd_sc_hd__nor2_1 _4802_ (.A(_1226_),
    .B(_1228_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand3_1 _4803_ (.A(_1223_),
    .B(_1220_),
    .C(_1221_),
    .Y(_1233_));
 sky130_fd_sc_hd__mux2_1 _4804_ (.A0(\as2650.r123[0][7] ),
    .A1(\as2650.r123_2[0][7] ),
    .S(_3161_),
    .X(_1234_));
 sky130_fd_sc_hd__a22o_1 _4805_ (.A1(_3261_),
    .A2(_1234_),
    .B1(_0735_),
    .B2(\as2650.r0[1] ),
    .X(_1235_));
 sky130_fd_sc_hd__nand4_1 _4806_ (.A(_3390_),
    .B(_3261_),
    .C(_1234_),
    .D(_0735_),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_0325_),
    .B(_0730_),
    .Y(_1237_));
 sky130_fd_sc_hd__a21bo_1 _4808_ (.A1(_1235_),
    .A2(_1236_),
    .B1_N(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__nand3b_1 _4809_ (.A_N(_1237_),
    .B(_1235_),
    .C(_1236_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand3_1 _4810_ (.A(_1207_),
    .B(_1238_),
    .C(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__a21o_1 _4811_ (.A1(_1238_),
    .A2(_1239_),
    .B1(_1207_),
    .X(_1241_));
 sky130_fd_sc_hd__nand2_1 _4812_ (.A(\as2650.r0[5] ),
    .B(_0711_),
    .Y(_1242_));
 sky130_fd_sc_hd__a22oi_1 _4813_ (.A1(_0469_),
    .A2(_0718_),
    .B1(_0724_),
    .B2(_0348_),
    .Y(_1243_));
 sky130_fd_sc_hd__and4_1 _4814_ (.A(\as2650.r0[4] ),
    .B(\as2650.r0[3] ),
    .C(_0717_),
    .D(_0723_),
    .X(_1244_));
 sky130_fd_sc_hd__nor2_1 _4815_ (.A(_1243_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__xnor2_1 _4816_ (.A(_1242_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a21oi_1 _4817_ (.A1(_1240_),
    .A2(_1241_),
    .B1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__and3_1 _4818_ (.A(_1240_),
    .B(_1241_),
    .C(_1246_),
    .X(_1248_));
 sky130_fd_sc_hd__or3_1 _4819_ (.A(_1209_),
    .B(_1247_),
    .C(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__o21ai_1 _4820_ (.A1(_1247_),
    .A2(_1248_),
    .B1(_1209_),
    .Y(_1250_));
 sky130_fd_sc_hd__a21bo_1 _4821_ (.A1(_1201_),
    .A2(_1203_),
    .B1_N(_1202_),
    .X(_1251_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(\as2650.r0[6] ),
    .B(_0706_),
    .Y(_1252_));
 sky130_fd_sc_hd__xnor2_1 _4823_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__and3_1 _4824_ (.A(\as2650.r0[7] ),
    .B(_0696_),
    .C(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a21oi_1 _4825_ (.A1(_0617_),
    .A2(_0696_),
    .B1(_1253_),
    .Y(_1255_));
 sky130_fd_sc_hd__nor2_1 _4826_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__a21oi_1 _4827_ (.A1(_1249_),
    .A2(_1250_),
    .B1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__and3_1 _4828_ (.A(_1249_),
    .B(_1250_),
    .C(_1256_),
    .X(_1258_));
 sky130_fd_sc_hd__o211ai_1 _4829_ (.A1(_1257_),
    .A2(_1258_),
    .B1(_1211_),
    .C1(_1219_),
    .Y(_1259_));
 sky130_fd_sc_hd__a211o_1 _4830_ (.A1(_1211_),
    .A2(_1219_),
    .B1(_1257_),
    .C1(_1258_),
    .X(_1260_));
 sky130_fd_sc_hd__and3_1 _4831_ (.A(_0513_),
    .B(_0707_),
    .C(_1214_),
    .X(_1261_));
 sky130_fd_sc_hd__a31o_1 _4832_ (.A1(_0544_),
    .A2(_0696_),
    .A3(_1216_),
    .B1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__a21oi_1 _4833_ (.A1(_1259_),
    .A2(_1260_),
    .B1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__and3_1 _4834_ (.A(_1262_),
    .B(_1259_),
    .C(_1260_),
    .X(_1264_));
 sky130_fd_sc_hd__a211o_1 _4835_ (.A1(_1220_),
    .A2(_1233_),
    .B1(_1263_),
    .C1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__o211ai_1 _4836_ (.A1(_1263_),
    .A2(_1264_),
    .B1(_1220_),
    .C1(_1233_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_1265_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__xor2_2 _4838_ (.A(_1232_),
    .B(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_1 _4839_ (.A1(_0871_),
    .A2(_1115_),
    .B1(_1117_),
    .B2(\as2650.r123_2[1][7] ),
    .X(_1269_));
 sky130_fd_sc_hd__a21o_1 _4840_ (.A1(_1121_),
    .A2(_1268_),
    .B1(_1269_),
    .X(_0083_));
 sky130_fd_sc_hd__or2_1 _4841_ (.A(_0317_),
    .B(_3352_),
    .X(_1270_));
 sky130_fd_sc_hd__or2_2 _4842_ (.A(_0932_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__or2_2 _4843_ (.A(_0725_),
    .B(_1270_),
    .X(_1272_));
 sky130_fd_sc_hd__nand2_4 _4844_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(\as2650.stack[1][8] ),
    .A1(_0699_),
    .S(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _4846_ (.A(_1274_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4847_ (.A0(\as2650.stack[1][9] ),
    .A1(_0709_),
    .S(_1273_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _4848_ (.A(_1275_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(\as2650.stack[1][10] ),
    .A1(_0715_),
    .S(_1273_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _4850_ (.A(_1276_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4851_ (.A0(\as2650.stack[1][11] ),
    .A1(_0721_),
    .S(_1273_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _4852_ (.A(_1277_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4853_ (.A0(\as2650.stack[1][12] ),
    .A1(_0728_),
    .S(_1273_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _4854_ (.A(_1278_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4855_ (.A0(\as2650.stack[1][13] ),
    .A1(_0733_),
    .S(_1273_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _4856_ (.A(_1279_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(\as2650.stack[1][14] ),
    .A1(_0738_),
    .S(_1273_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _4858_ (.A(_1280_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(_0700_),
    .B(_3335_),
    .Y(_1281_));
 sky130_fd_sc_hd__or2_2 _4860_ (.A(_0932_),
    .B(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__or2_2 _4861_ (.A(_0725_),
    .B(_1281_),
    .X(_1283_));
 sky130_fd_sc_hd__nand2_4 _4862_ (.A(_1282_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(\as2650.stack[0][8] ),
    .A1(_0699_),
    .S(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _4864_ (.A(_1285_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4865_ (.A0(\as2650.stack[0][9] ),
    .A1(_0709_),
    .S(_1284_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _4866_ (.A(_1286_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(\as2650.stack[0][10] ),
    .A1(_0715_),
    .S(_1284_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _4868_ (.A(_1287_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(\as2650.stack[0][11] ),
    .A1(_0721_),
    .S(_1284_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _4870_ (.A(_1288_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4871_ (.A0(\as2650.stack[0][12] ),
    .A1(_0728_),
    .S(_1284_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4872_ (.A(_1289_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(\as2650.stack[0][13] ),
    .A1(_0733_),
    .S(_1284_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _4874_ (.A(_1290_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4875_ (.A0(\as2650.stack[0][14] ),
    .A1(_0738_),
    .S(_1284_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _4876_ (.A(_1291_),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _4877_ (.A(\as2650.r123_2[3][0] ),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _4878_ (.A(_1292_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _4879_ (.A(\as2650.r123_2[3][1] ),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _4880_ (.A(_1293_),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_1 _4881_ (.A(\as2650.r123_2[3][2] ),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _4882_ (.A(_1294_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _4883_ (.A(\as2650.r123_2[3][3] ),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _4884_ (.A(_1295_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _4885_ (.A(\as2650.r123_2[3][4] ),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _4886_ (.A(_1296_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _4887_ (.A(\as2650.r123_2[3][5] ),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _4888_ (.A(_1297_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _4889_ (.A(\as2650.r123_2[3][6] ),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _4890_ (.A(_1298_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _4891_ (.A(\as2650.r123_2[3][7] ),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _4892_ (.A(_1299_),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _4893_ (.A(_3073_),
    .B(_0756_),
    .X(_1300_));
 sky130_fd_sc_hd__buf_2 _4894_ (.A(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__a211oi_1 _4895_ (.A1(_1220_),
    .A2(_1233_),
    .B1(_1263_),
    .C1(_1264_),
    .Y(_1302_));
 sky130_fd_sc_hd__o211a_1 _4896_ (.A1(_1226_),
    .A2(_1228_),
    .B1(_1265_),
    .C1(_1266_),
    .X(_1303_));
 sky130_fd_sc_hd__and3_1 _4897_ (.A(_0544_),
    .B(_0707_),
    .C(_1251_),
    .X(_1304_));
 sky130_fd_sc_hd__nand3_1 _4898_ (.A(_1249_),
    .B(_1250_),
    .C(_1256_),
    .Y(_1305_));
 sky130_fd_sc_hd__and3_1 _4899_ (.A(_0512_),
    .B(_0712_),
    .C(_1245_),
    .X(_1306_));
 sky130_fd_sc_hd__o211a_1 _4900_ (.A1(_1244_),
    .A2(_1306_),
    .B1(_0617_),
    .C1(_0707_),
    .X(_1307_));
 sky130_fd_sc_hd__a211oi_1 _4901_ (.A1(_0617_),
    .A2(_0707_),
    .B1(_1244_),
    .C1(_1306_),
    .Y(_1308_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(_1307_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__a22oi_1 _4903_ (.A1(_0512_),
    .A2(_0718_),
    .B1(_0724_),
    .B2(_0469_),
    .Y(_1310_));
 sky130_fd_sc_hd__and4_1 _4904_ (.A(\as2650.r0[5] ),
    .B(_0469_),
    .C(_0718_),
    .D(_0724_),
    .X(_1311_));
 sky130_fd_sc_hd__or2_1 _4905_ (.A(_1310_),
    .B(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(\as2650.r0[6] ),
    .B(_0712_),
    .Y(_1313_));
 sky130_fd_sc_hd__xnor2_1 _4907_ (.A(_1312_),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__clkbuf_4 _4908_ (.A(_1234_),
    .X(_1315_));
 sky130_fd_sc_hd__and4_1 _4909_ (.A(_0325_),
    .B(_3390_),
    .C(_1315_),
    .D(_0735_),
    .X(_1316_));
 sky130_fd_sc_hd__a22oi_1 _4910_ (.A1(_3390_),
    .A2(_1315_),
    .B1(_0736_),
    .B2(_0325_),
    .Y(_1317_));
 sky130_fd_sc_hd__nor2_1 _4911_ (.A(_1316_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(_0417_),
    .B(_0730_),
    .Y(_1319_));
 sky130_fd_sc_hd__xnor2_1 _4913_ (.A(_1318_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__and2_1 _4914_ (.A(_1236_),
    .B(_1239_),
    .X(_1321_));
 sky130_fd_sc_hd__xor2_1 _4915_ (.A(_1320_),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__xor2_1 _4916_ (.A(_1314_),
    .B(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a21boi_1 _4917_ (.A1(_1241_),
    .A2(_1246_),
    .B1_N(_1240_),
    .Y(_1324_));
 sky130_fd_sc_hd__xnor2_1 _4918_ (.A(_1323_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__and2_1 _4919_ (.A(_1309_),
    .B(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__nor2_1 _4920_ (.A(_1309_),
    .B(_1325_),
    .Y(_1327_));
 sky130_fd_sc_hd__a211o_1 _4921_ (.A1(_1249_),
    .A2(_1305_),
    .B1(_1326_),
    .C1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__o211ai_1 _4922_ (.A1(_1326_),
    .A2(_1327_),
    .B1(_1249_),
    .C1(_1305_),
    .Y(_1329_));
 sky130_fd_sc_hd__o211ai_2 _4923_ (.A1(_1304_),
    .A2(_1254_),
    .B1(_1328_),
    .C1(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a211o_1 _4924_ (.A1(_1328_),
    .A2(_1329_),
    .B1(_1304_),
    .C1(_1254_),
    .X(_1331_));
 sky130_fd_sc_hd__a21bo_1 _4925_ (.A1(_1262_),
    .A2(_1259_),
    .B1_N(_1260_),
    .X(_1332_));
 sky130_fd_sc_hd__nand3_1 _4926_ (.A(_1330_),
    .B(_1331_),
    .C(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__a21o_1 _4927_ (.A1(_1330_),
    .A2(_1331_),
    .B1(_1332_),
    .X(_1334_));
 sky130_fd_sc_hd__o211ai_1 _4928_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1333_),
    .C1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__a211o_1 _4929_ (.A1(_1333_),
    .A2(_1334_),
    .B1(_1302_),
    .C1(_1303_),
    .X(_1336_));
 sky130_fd_sc_hd__and2_1 _4930_ (.A(_1335_),
    .B(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__inv_2 _4931_ (.A(_1301_),
    .Y(_1338_));
 sky130_fd_sc_hd__nor2_2 _4932_ (.A(_1116_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__a22oi_1 _4933_ (.A1(_1118_),
    .A2(_1337_),
    .B1(_1339_),
    .B2(\as2650.r123_2[2][0] ),
    .Y(_1340_));
 sky130_fd_sc_hd__o21ai_1 _4934_ (.A1(_0791_),
    .A2(_1301_),
    .B1(_1340_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ba_1 _4935_ (.A1(_1310_),
    .A2(_1313_),
    .B1_N(_1311_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(\as2650.r0[2] ),
    .B(_1234_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_0348_),
    .B(_0735_),
    .Y(_1343_));
 sky130_fd_sc_hd__xor2_1 _4938_ (.A(_1342_),
    .B(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__and3_1 _4939_ (.A(_0469_),
    .B(_0730_),
    .C(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__a21oi_1 _4940_ (.A1(_0470_),
    .A2(_0731_),
    .B1(_1344_),
    .Y(_1346_));
 sky130_fd_sc_hd__nor2_1 _4941_ (.A(_1345_),
    .B(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__a31o_1 _4942_ (.A1(_0417_),
    .A2(_0731_),
    .A3(_1318_),
    .B1(_1316_),
    .X(_1348_));
 sky130_fd_sc_hd__xnor2_1 _4943_ (.A(_1347_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4944_ (.A(\as2650.r0[5] ),
    .B(_0724_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(\as2650.r0[6] ),
    .B(_0718_),
    .Y(_1351_));
 sky130_fd_sc_hd__xor2_1 _4946_ (.A(_1350_),
    .B(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__and3_1 _4947_ (.A(\as2650.r0[7] ),
    .B(_0712_),
    .C(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__a21oi_1 _4948_ (.A1(\as2650.r0[7] ),
    .A2(_0712_),
    .B1(_1352_),
    .Y(_1354_));
 sky130_fd_sc_hd__or2_1 _4949_ (.A(_1353_),
    .B(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__xor2_1 _4950_ (.A(_1349_),
    .B(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__or2b_1 _4951_ (.A(_1321_),
    .B_N(_1320_),
    .X(_1357_));
 sky130_fd_sc_hd__o21a_1 _4952_ (.A1(_1314_),
    .A2(_1322_),
    .B1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__xnor2_1 _4953_ (.A(_1356_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__xnor2_1 _4954_ (.A(_1341_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__and2b_1 _4955_ (.A_N(_1324_),
    .B(_1323_),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_1 _4956_ (.A(_1361_),
    .B(_1326_),
    .Y(_1362_));
 sky130_fd_sc_hd__xnor2_1 _4957_ (.A(_1360_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__xnor2_1 _4958_ (.A(_1307_),
    .B(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(_1328_),
    .B(_1330_),
    .Y(_1365_));
 sky130_fd_sc_hd__xor2_1 _4960_ (.A(_1364_),
    .B(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__a21o_1 _4961_ (.A1(_1333_),
    .A2(_1335_),
    .B1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nand3_1 _4962_ (.A(_1333_),
    .B(_1335_),
    .C(_1366_),
    .Y(_1368_));
 sky130_fd_sc_hd__and2_1 _4963_ (.A(_1367_),
    .B(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a22oi_1 _4964_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1339_),
    .B1(_1369_),
    .B2(_1121_),
    .Y(_1370_));
 sky130_fd_sc_hd__o21ai_1 _4965_ (.A1(_0802_),
    .A2(_1301_),
    .B1(_1370_),
    .Y(_0107_));
 sky130_fd_sc_hd__or2b_1 _4966_ (.A(_1364_),
    .B_N(_1365_),
    .X(_1371_));
 sky130_fd_sc_hd__and2b_1 _4967_ (.A_N(_1362_),
    .B(_1360_),
    .X(_1372_));
 sky130_fd_sc_hd__and2_1 _4968_ (.A(_1307_),
    .B(_1363_),
    .X(_1373_));
 sky130_fd_sc_hd__and2_1 _4969_ (.A(_1347_),
    .B(_1348_),
    .X(_1374_));
 sky130_fd_sc_hd__nor2_1 _4970_ (.A(_1349_),
    .B(_1355_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0348_),
    .B(_1315_),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_0469_),
    .B(_0736_),
    .Y(_1377_));
 sky130_fd_sc_hd__xor2_1 _4973_ (.A(_1376_),
    .B(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__and3_1 _4974_ (.A(_0512_),
    .B(_0731_),
    .C(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__a21oi_1 _4975_ (.A1(_0512_),
    .A2(_0731_),
    .B1(_1378_),
    .Y(_1380_));
 sky130_fd_sc_hd__nor2_1 _4976_ (.A(_1379_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__o21bai_1 _4977_ (.A1(_1342_),
    .A2(_1343_),
    .B1_N(_1345_),
    .Y(_1382_));
 sky130_fd_sc_hd__xnor2_1 _4978_ (.A(_1381_),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0617_),
    .B(_0724_),
    .Y(_1384_));
 sky130_fd_sc_hd__a22o_1 _4980_ (.A1(_0617_),
    .A2(_0718_),
    .B1(_0724_),
    .B2(_0544_),
    .X(_1385_));
 sky130_fd_sc_hd__o21ai_1 _4981_ (.A1(_1351_),
    .A2(_1384_),
    .B1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__xor2_1 _4982_ (.A(_1383_),
    .B(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__o21a_1 _4983_ (.A1(_1374_),
    .A2(_1375_),
    .B1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__nor3_1 _4984_ (.A(_1374_),
    .B(_1375_),
    .C(_1387_),
    .Y(_1389_));
 sky130_fd_sc_hd__nor2_1 _4985_ (.A(_1388_),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__o21ba_1 _4986_ (.A1(_1350_),
    .A2(_1351_),
    .B1_N(_1353_),
    .X(_1391_));
 sky130_fd_sc_hd__xnor2_1 _4987_ (.A(_1390_),
    .B(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and2b_1 _4988_ (.A_N(_1358_),
    .B(_1356_),
    .X(_1393_));
 sky130_fd_sc_hd__and2b_1 _4989_ (.A_N(_1341_),
    .B(_1359_),
    .X(_1394_));
 sky130_fd_sc_hd__nor2_1 _4990_ (.A(_1393_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__xnor2_1 _4991_ (.A(_1392_),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__o21a_1 _4992_ (.A1(_1372_),
    .A2(_1373_),
    .B1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__nor3_1 _4993_ (.A(_1372_),
    .B(_1373_),
    .C(_1396_),
    .Y(_1398_));
 sky130_fd_sc_hd__or2_1 _4994_ (.A(_1397_),
    .B(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__a21oi_2 _4995_ (.A1(_1371_),
    .A2(_1367_),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__and3_1 _4996_ (.A(_1371_),
    .B(_1367_),
    .C(_1399_),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_1400_),
    .B(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__a22oi_1 _4998_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_1339_),
    .B1(_1402_),
    .B2(_1118_),
    .Y(_1403_));
 sky130_fd_sc_hd__o21ai_1 _4999_ (.A1(_0815_),
    .A2(_1301_),
    .B1(_1403_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_1 _5000_ (.A(_1351_),
    .B(_1384_),
    .Y(_1404_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_0512_),
    .B(_1315_),
    .Y(_1405_));
 sky130_fd_sc_hd__a22o_1 _5002_ (.A1(_0469_),
    .A2(_1315_),
    .B1(_0736_),
    .B2(_0512_),
    .X(_1406_));
 sky130_fd_sc_hd__o21a_1 _5003_ (.A1(_1377_),
    .A2(_1405_),
    .B1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__and3_1 _5004_ (.A(_0544_),
    .B(_0731_),
    .C(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__a21oi_1 _5005_ (.A1(_0544_),
    .A2(_0731_),
    .B1(_1407_),
    .Y(_1409_));
 sky130_fd_sc_hd__or2_1 _5006_ (.A(_1408_),
    .B(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__o21ba_1 _5007_ (.A1(_1376_),
    .A2(_1377_),
    .B1_N(_1379_),
    .X(_1411_));
 sky130_fd_sc_hd__xnor2_1 _5008_ (.A(_1410_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__xnor2_1 _5009_ (.A(_1384_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__o2bb2a_1 _5010_ (.A1_N(_1381_),
    .A2_N(_1382_),
    .B1(_1383_),
    .B2(_1386_),
    .X(_1414_));
 sky130_fd_sc_hd__xor2_1 _5011_ (.A(_1413_),
    .B(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__nand2_1 _5012_ (.A(_1404_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__or2_1 _5013_ (.A(_1404_),
    .B(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__nand2_1 _5014_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__o21ba_1 _5015_ (.A1(_1389_),
    .A2(_1391_),
    .B1_N(_1388_),
    .X(_1419_));
 sky130_fd_sc_hd__or2_1 _5016_ (.A(_1418_),
    .B(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_1418_),
    .B(_1419_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_1420_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__inv_2 _5019_ (.A(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__and2b_1 _5020_ (.A_N(_1395_),
    .B(_1392_),
    .X(_1424_));
 sky130_fd_sc_hd__nor2_1 _5021_ (.A(_1424_),
    .B(_1397_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux2_1 _5022_ (.A0(_1425_),
    .A1(_1424_),
    .S(_1400_),
    .X(_1426_));
 sky130_fd_sc_hd__xnor2_2 _5023_ (.A(_1423_),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__a22oi_1 _5024_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_1339_),
    .B1(_1427_),
    .B2(_1118_),
    .Y(_1428_));
 sky130_fd_sc_hd__o21ai_1 _5025_ (.A1(_0827_),
    .A2(_1301_),
    .B1(_1428_),
    .Y(_0109_));
 sky130_fd_sc_hd__nor2_1 _5026_ (.A(_1377_),
    .B(_1405_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_0544_),
    .B(_0736_),
    .Y(_1430_));
 sky130_fd_sc_hd__xor2_1 _5028_ (.A(_1405_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__and3_1 _5029_ (.A(_0617_),
    .B(_0731_),
    .C(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a21oi_1 _5030_ (.A1(_0617_),
    .A2(_0731_),
    .B1(_1431_),
    .Y(_1433_));
 sky130_fd_sc_hd__nor2_1 _5031_ (.A(_1432_),
    .B(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__o21ai_2 _5032_ (.A1(_1429_),
    .A2(_1408_),
    .B1(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__or3_1 _5033_ (.A(_1429_),
    .B(_1408_),
    .C(_1434_),
    .X(_1436_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_1435_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__o32a_1 _5035_ (.A1(_1408_),
    .A2(_1409_),
    .A3(_1411_),
    .B1(_1412_),
    .B2(_1384_),
    .X(_1438_));
 sky130_fd_sc_hd__xor2_1 _5036_ (.A(_1437_),
    .B(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__o21a_1 _5037_ (.A1(_1413_),
    .A2(_1414_),
    .B1(_1416_),
    .X(_1440_));
 sky130_fd_sc_hd__xor2_1 _5038_ (.A(_1439_),
    .B(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__nor2_1 _5039_ (.A(_1420_),
    .B(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__and2_1 _5040_ (.A(_1420_),
    .B(_1441_),
    .X(_1443_));
 sky130_fd_sc_hd__nor2_1 _5041_ (.A(_1442_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__o31ai_2 _5042_ (.A1(_1424_),
    .A2(_1397_),
    .A3(_1400_),
    .B1(_1423_),
    .Y(_1445_));
 sky130_fd_sc_hd__xnor2_2 _5043_ (.A(_1444_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__a22oi_1 _5044_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1339_),
    .B1(_1446_),
    .B2(_1118_),
    .Y(_1447_));
 sky130_fd_sc_hd__o21ai_1 _5045_ (.A1(_0838_),
    .A2(_1301_),
    .B1(_1447_),
    .Y(_0110_));
 sky130_fd_sc_hd__o311a_1 _5046_ (.A1(_1424_),
    .A2(_1397_),
    .A3(_1400_),
    .B1(_1423_),
    .C1(_1444_),
    .X(_1448_));
 sky130_fd_sc_hd__or2b_1 _5047_ (.A(_1440_),
    .B_N(_1439_),
    .X(_1449_));
 sky130_fd_sc_hd__o21bai_2 _5048_ (.A1(_1405_),
    .A2(_1430_),
    .B1_N(_1432_),
    .Y(_1450_));
 sky130_fd_sc_hd__a22oi_1 _5049_ (.A1(_0545_),
    .A2(_1315_),
    .B1(_0736_),
    .B2(_0617_),
    .Y(_1451_));
 sky130_fd_sc_hd__and4_1 _5050_ (.A(_0617_),
    .B(_0544_),
    .C(_1315_),
    .D(_0736_),
    .X(_1452_));
 sky130_fd_sc_hd__nor2_1 _5051_ (.A(_1451_),
    .B(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__xnor2_2 _5052_ (.A(_1450_),
    .B(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__o21ai_1 _5053_ (.A1(_1437_),
    .A2(_1438_),
    .B1(_1435_),
    .Y(_1455_));
 sky130_fd_sc_hd__xnor2_1 _5054_ (.A(_1454_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__xnor2_1 _5055_ (.A(_1449_),
    .B(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__o21ai_1 _5056_ (.A1(_1442_),
    .A2(_1448_),
    .B1(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__or3_1 _5057_ (.A(_1442_),
    .B(_1448_),
    .C(_1457_),
    .X(_1459_));
 sky130_fd_sc_hd__and2_1 _5058_ (.A(_1458_),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a22oi_1 _5059_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_1339_),
    .B1(_1460_),
    .B2(_1118_),
    .Y(_1461_));
 sky130_fd_sc_hd__o21ai_1 _5060_ (.A1(_0849_),
    .A2(_1301_),
    .B1(_1461_),
    .Y(_0111_));
 sky130_fd_sc_hd__or2b_1 _5061_ (.A(_1449_),
    .B_N(_1456_),
    .X(_1462_));
 sky130_fd_sc_hd__or3_2 _5062_ (.A(_1437_),
    .B(_1438_),
    .C(_1454_),
    .X(_1463_));
 sky130_fd_sc_hd__and3_1 _5063_ (.A(_0618_),
    .B(_1315_),
    .C(_1430_),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_1450_),
    .B(_1453_),
    .Y(_1465_));
 sky130_fd_sc_hd__o21ai_2 _5065_ (.A1(_1435_),
    .A2(_1454_),
    .B1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__xnor2_2 _5066_ (.A(_1464_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__xnor2_1 _5067_ (.A(_1463_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__a21o_1 _5068_ (.A1(_1462_),
    .A2(_1458_),
    .B1(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__nand3_1 _5069_ (.A(_1462_),
    .B(_1458_),
    .C(_1468_),
    .Y(_1470_));
 sky130_fd_sc_hd__and2_1 _5070_ (.A(_1469_),
    .B(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__a2bb2o_1 _5071_ (.A1_N(_0859_),
    .A2_N(_1301_),
    .B1(_1339_),
    .B2(\as2650.r123_2[2][6] ),
    .X(_1472_));
 sky130_fd_sc_hd__a21o_1 _5072_ (.A1(_1121_),
    .A2(_1471_),
    .B1(_1472_),
    .X(_0112_));
 sky130_fd_sc_hd__a21oi_1 _5073_ (.A1(_0545_),
    .A2(_0736_),
    .B1(_1466_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_0684_),
    .B(_1315_),
    .Y(_1474_));
 sky130_fd_sc_hd__o221ai_4 _5075_ (.A1(_1463_),
    .A2(_1467_),
    .B1(_1473_),
    .B2(_1474_),
    .C1(_1469_),
    .Y(_1475_));
 sky130_fd_sc_hd__a22o_1 _5076_ (.A1(_0871_),
    .A2(_1338_),
    .B1(_1339_),
    .B2(\as2650.r123_2[2][7] ),
    .X(_1476_));
 sky130_fd_sc_hd__a21o_1 _5077_ (.A1(_1121_),
    .A2(_1475_),
    .B1(_1476_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5078_ (.A0(_0636_),
    .A1(\as2650.stack[4][0] ),
    .S(_0933_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _5079_ (.A0(_0634_),
    .A1(_1477_),
    .S(_0923_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _5080_ (.A(_1478_),
    .X(_0114_));
 sky130_fd_sc_hd__nor3_4 _5081_ (.A(_0700_),
    .B(_3352_),
    .C(_0697_),
    .Y(_1479_));
 sky130_fd_sc_hd__nor2_4 _5082_ (.A(_3336_),
    .B(_0932_),
    .Y(_1480_));
 sky130_fd_sc_hd__or2_1 _5083_ (.A(\as2650.stack[4][1] ),
    .B(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__o21a_1 _5084_ (.A1(_0661_),
    .A2(_0933_),
    .B1(_0923_),
    .X(_1482_));
 sky130_fd_sc_hd__a22o_1 _5085_ (.A1(_0659_),
    .A2(_1479_),
    .B1(_1481_),
    .B2(_1482_),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _5086_ (.A(\as2650.stack[4][2] ),
    .B(_1480_),
    .X(_1483_));
 sky130_fd_sc_hd__inv_2 _5087_ (.A(\as2650.pc[2] ),
    .Y(_1484_));
 sky130_fd_sc_hd__a21oi_1 _5088_ (.A1(_1484_),
    .A2(_1480_),
    .B1(_1479_),
    .Y(_1485_));
 sky130_fd_sc_hd__a22o_1 _5089_ (.A1(_0664_),
    .A2(_1479_),
    .B1(_1483_),
    .B2(_1485_),
    .X(_0116_));
 sky130_fd_sc_hd__or2_1 _5090_ (.A(\as2650.stack[4][3] ),
    .B(_1480_),
    .X(_1486_));
 sky130_fd_sc_hd__inv_2 _5091_ (.A(\as2650.pc[3] ),
    .Y(_1487_));
 sky130_fd_sc_hd__a21oi_1 _5092_ (.A1(_1487_),
    .A2(_1480_),
    .B1(_1479_),
    .Y(_1488_));
 sky130_fd_sc_hd__a22o_1 _5093_ (.A1(_0667_),
    .A2(_1479_),
    .B1(_1486_),
    .B2(_1488_),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _5094_ (.A(\as2650.stack[4][4] ),
    .B(_1480_),
    .X(_1489_));
 sky130_fd_sc_hd__inv_2 _5095_ (.A(\as2650.pc[4] ),
    .Y(_1490_));
 sky130_fd_sc_hd__a21oi_1 _5096_ (.A1(_1490_),
    .A2(_1480_),
    .B1(_1479_),
    .Y(_1491_));
 sky130_fd_sc_hd__a22o_1 _5097_ (.A1(_0671_),
    .A2(_1479_),
    .B1(_1489_),
    .B2(_1491_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_1 _5098_ (.A(\as2650.stack[4][5] ),
    .B(_1480_),
    .X(_1492_));
 sky130_fd_sc_hd__o21a_1 _5099_ (.A1(_0676_),
    .A2(_0933_),
    .B1(_0923_),
    .X(_1493_));
 sky130_fd_sc_hd__a22o_1 _5100_ (.A1(_0675_),
    .A2(_1479_),
    .B1(_1492_),
    .B2(_1493_),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _5101_ (.A(\as2650.stack[4][6] ),
    .B(_1480_),
    .X(_1494_));
 sky130_fd_sc_hd__o21a_1 _5102_ (.A1(_0681_),
    .A2(_0933_),
    .B1(_0923_),
    .X(_1495_));
 sky130_fd_sc_hd__a22o_1 _5103_ (.A1(_0679_),
    .A2(_1479_),
    .B1(_1494_),
    .B2(_1495_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _5104_ (.A(\as2650.stack[4][7] ),
    .B(_1480_),
    .X(_1496_));
 sky130_fd_sc_hd__o21a_1 _5105_ (.A1(_0685_),
    .A2(_0933_),
    .B1(_0923_),
    .X(_1497_));
 sky130_fd_sc_hd__a22o_1 _5106_ (.A1(_0684_),
    .A2(_1479_),
    .B1(_1496_),
    .B2(_1497_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(_0636_),
    .A1(\as2650.stack[2][0] ),
    .S(_1104_),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(_0634_),
    .A1(_1498_),
    .S(_1080_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _5109_ (.A(_1499_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(_0661_),
    .A1(\as2650.stack[2][1] ),
    .S(_1104_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(_0659_),
    .A1(_1500_),
    .S(_1080_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _5112_ (.A(_1501_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(\as2650.pc[2] ),
    .A1(\as2650.stack[2][2] ),
    .S(_1104_),
    .X(_1502_));
 sky130_fd_sc_hd__or3_2 _5114_ (.A(_3056_),
    .B(_0692_),
    .C(_1079_),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(_0664_),
    .A1(_1502_),
    .S(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _5116_ (.A(_1504_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(_0668_),
    .A1(\as2650.stack[2][3] ),
    .S(_1104_),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(_0667_),
    .A1(_1505_),
    .S(_1503_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _5119_ (.A(_1506_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(_0672_),
    .A1(\as2650.stack[2][4] ),
    .S(_1104_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(_0671_),
    .A1(_1507_),
    .S(_1080_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _5122_ (.A(_1508_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(_0676_),
    .A1(\as2650.stack[2][5] ),
    .S(_1104_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _5124_ (.A0(_0675_),
    .A1(_1509_),
    .S(_1080_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _5125_ (.A(_1510_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(_0681_),
    .A1(\as2650.stack[2][6] ),
    .S(_1104_),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(_0679_),
    .A1(_1511_),
    .S(_1080_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _5128_ (.A(_1512_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(_0685_),
    .A1(\as2650.stack[2][7] ),
    .S(_1104_),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _5130_ (.A0(_0684_),
    .A1(_1513_),
    .S(_1503_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _5131_ (.A(_1514_),
    .X(_0129_));
 sky130_fd_sc_hd__nor3_2 _5132_ (.A(_0317_),
    .B(_0329_),
    .C(_0697_),
    .Y(_1515_));
 sky130_fd_sc_hd__buf_2 _5133_ (.A(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__nor2_1 _5134_ (.A(_0932_),
    .B(_1270_),
    .Y(_1517_));
 sky130_fd_sc_hd__buf_2 _5135_ (.A(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__or2_1 _5136_ (.A(\as2650.stack[1][0] ),
    .B(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__inv_2 _5137_ (.A(_0635_),
    .Y(_1520_));
 sky130_fd_sc_hd__a21oi_1 _5138_ (.A1(_1520_),
    .A2(_1518_),
    .B1(_1516_),
    .Y(_1521_));
 sky130_fd_sc_hd__a22o_1 _5139_ (.A1(_0634_),
    .A2(_1516_),
    .B1(_1519_),
    .B2(_1521_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_1 _5140_ (.A(\as2650.stack[1][1] ),
    .B(_1518_),
    .X(_1522_));
 sky130_fd_sc_hd__o21a_1 _5141_ (.A1(_0661_),
    .A2(_1271_),
    .B1(_1105_),
    .X(_1523_));
 sky130_fd_sc_hd__a22o_1 _5142_ (.A1(_0659_),
    .A2(_1516_),
    .B1(_1522_),
    .B2(_1523_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _5143_ (.A(\as2650.stack[1][2] ),
    .B(_1518_),
    .X(_1524_));
 sky130_fd_sc_hd__a21oi_1 _5144_ (.A1(_1484_),
    .A2(_1518_),
    .B1(_1516_),
    .Y(_1525_));
 sky130_fd_sc_hd__a22o_1 _5145_ (.A1(_0664_),
    .A2(_1516_),
    .B1(_1524_),
    .B2(_1525_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _5146_ (.A(\as2650.stack[1][3] ),
    .B(_1518_),
    .X(_1526_));
 sky130_fd_sc_hd__a21oi_1 _5147_ (.A1(_1487_),
    .A2(_1518_),
    .B1(_1515_),
    .Y(_1527_));
 sky130_fd_sc_hd__a22o_1 _5148_ (.A1(_0667_),
    .A2(_1516_),
    .B1(_1526_),
    .B2(_1527_),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _5149_ (.A(\as2650.stack[1][4] ),
    .B(_1518_),
    .X(_1528_));
 sky130_fd_sc_hd__a21oi_1 _5150_ (.A1(_1490_),
    .A2(_1518_),
    .B1(_1515_),
    .Y(_1529_));
 sky130_fd_sc_hd__a22o_1 _5151_ (.A1(_0671_),
    .A2(_1516_),
    .B1(_1528_),
    .B2(_1529_),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _5152_ (.A(\as2650.stack[1][5] ),
    .B(_1518_),
    .X(_1530_));
 sky130_fd_sc_hd__o21a_1 _5153_ (.A1(_0676_),
    .A2(_1271_),
    .B1(_1105_),
    .X(_1531_));
 sky130_fd_sc_hd__a22o_1 _5154_ (.A1(_0675_),
    .A2(_1516_),
    .B1(_1530_),
    .B2(_1531_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _5155_ (.A(\as2650.stack[1][6] ),
    .B(_1517_),
    .X(_1532_));
 sky130_fd_sc_hd__o21a_1 _5156_ (.A1(_0681_),
    .A2(_1271_),
    .B1(_1105_),
    .X(_1533_));
 sky130_fd_sc_hd__a22o_1 _5157_ (.A1(_0679_),
    .A2(_1516_),
    .B1(_1532_),
    .B2(_1533_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _5158_ (.A(\as2650.stack[1][7] ),
    .B(_1517_),
    .X(_1534_));
 sky130_fd_sc_hd__o21a_1 _5159_ (.A1(_0685_),
    .A2(_1271_),
    .B1(_1105_),
    .X(_1535_));
 sky130_fd_sc_hd__a22o_1 _5160_ (.A1(_0684_),
    .A2(_1516_),
    .B1(_1534_),
    .B2(_1535_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _5161_ (.A(\as2650.r123[3][0] ),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _5162_ (.A(_1536_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _5163_ (.A(\as2650.r123[3][1] ),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _5164_ (.A(_1537_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _5165_ (.A(\as2650.r123[3][2] ),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_1538_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _5167_ (.A(\as2650.r123[3][3] ),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _5168_ (.A(_1539_),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(\as2650.r123[3][4] ),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _5170_ (.A(_1540_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _5171_ (.A(\as2650.r123[3][5] ),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _5172_ (.A(_1541_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _5173_ (.A(\as2650.r123[3][6] ),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _5174_ (.A(_1542_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _5175_ (.A(\as2650.r123[3][7] ),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _5176_ (.A(_1543_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _5177_ (.A0(_0636_),
    .A1(\as2650.stack[3][0] ),
    .S(_1081_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _5178_ (.A0(_0634_),
    .A1(_1544_),
    .S(_0934_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _5179_ (.A(_1545_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5180_ (.A0(_0661_),
    .A1(\as2650.stack[3][1] ),
    .S(_1081_),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(_0659_),
    .A1(_1546_),
    .S(_0934_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _5182_ (.A(_1547_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_2 _5183_ (.A(_3336_),
    .B(_0697_),
    .Y(_1548_));
 sky130_fd_sc_hd__nor2_2 _5184_ (.A(_0932_),
    .B(_1079_),
    .Y(_1549_));
 sky130_fd_sc_hd__or2_1 _5185_ (.A(\as2650.stack[3][2] ),
    .B(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__a21oi_1 _5186_ (.A1(_1484_),
    .A2(_1549_),
    .B1(_1548_),
    .Y(_1551_));
 sky130_fd_sc_hd__a22o_1 _5187_ (.A1(_0664_),
    .A2(_1548_),
    .B1(_1550_),
    .B2(_1551_),
    .X(_0148_));
 sky130_fd_sc_hd__or2_1 _5188_ (.A(\as2650.stack[3][3] ),
    .B(_1549_),
    .X(_1552_));
 sky130_fd_sc_hd__a21oi_1 _5189_ (.A1(_1487_),
    .A2(_1549_),
    .B1(_1548_),
    .Y(_1553_));
 sky130_fd_sc_hd__a22o_1 _5190_ (.A1(_0667_),
    .A2(_1548_),
    .B1(_1552_),
    .B2(_1553_),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _5191_ (.A(\as2650.stack[3][4] ),
    .B(_1549_),
    .X(_1554_));
 sky130_fd_sc_hd__a21oi_1 _5192_ (.A1(_1490_),
    .A2(_1549_),
    .B1(_1548_),
    .Y(_1555_));
 sky130_fd_sc_hd__a22o_1 _5193_ (.A1(_0671_),
    .A2(_1548_),
    .B1(_1554_),
    .B2(_1555_),
    .X(_0150_));
 sky130_fd_sc_hd__or2_1 _5194_ (.A(\as2650.stack[3][5] ),
    .B(_1549_),
    .X(_1556_));
 sky130_fd_sc_hd__o21a_1 _5195_ (.A1(_0676_),
    .A2(_1081_),
    .B1(_0934_),
    .X(_1557_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(_0675_),
    .A2(_1548_),
    .B1(_1556_),
    .B2(_1557_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(_0681_),
    .A1(\as2650.stack[3][6] ),
    .S(_1081_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _5198_ (.A0(_0679_),
    .A1(_1558_),
    .S(_0934_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _5199_ (.A(_1559_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5200_ (.A0(_0685_),
    .A1(\as2650.stack[3][7] ),
    .S(_1081_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(_0684_),
    .A1(_1560_),
    .S(_0934_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _5202_ (.A(_1561_),
    .X(_0153_));
 sky130_fd_sc_hd__buf_4 _5203_ (.A(_3153_),
    .X(_1562_));
 sky130_fd_sc_hd__and2_1 _5204_ (.A(_1562_),
    .B(\lfsr[1] ),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _5205_ (.A(_1563_),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _5206_ (.A(_0920_),
    .B(\lfsr[2] ),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _5207_ (.A(_1564_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _5208_ (.A(_1562_),
    .B(\lfsr[3] ),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _5209_ (.A(_1565_),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _5210_ (.A(_0920_),
    .B(\lfsr[4] ),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _5211_ (.A(_1566_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _5212_ (.A(_1562_),
    .B(\as2650.sense ),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _5213_ (.A(_1567_),
    .X(_0158_));
 sky130_fd_sc_hd__or2_1 _5214_ (.A(_0920_),
    .B(\lfsr[6] ),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _5215_ (.A(_1568_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _5216_ (.A(_1562_),
    .B(\lfsr[7] ),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _5217_ (.A(_1569_),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _5218_ (.A(_0920_),
    .B(\lfsr[8] ),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _5219_ (.A(_1570_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _5220_ (.A(_1562_),
    .B(\lfsr[9] ),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _5221_ (.A(_1571_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _5222_ (.A(_0920_),
    .B(\lfsr[10] ),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(_1572_),
    .X(_0163_));
 sky130_fd_sc_hd__a21oi_1 _5224_ (.A1(\lfsr[0] ),
    .A2(\lfsr[11] ),
    .B1(_0921_),
    .Y(_1573_));
 sky130_fd_sc_hd__o21a_1 _5225_ (.A1(\lfsr[0] ),
    .A2(\lfsr[11] ),
    .B1(_1573_),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _5226_ (.A(_0920_),
    .B(\lfsr[12] ),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _5227_ (.A(_1574_),
    .X(_0165_));
 sky130_fd_sc_hd__a21oi_1 _5228_ (.A1(\lfsr[0] ),
    .A2(\lfsr[13] ),
    .B1(_0921_),
    .Y(_1575_));
 sky130_fd_sc_hd__o21a_1 _5229_ (.A1(\lfsr[0] ),
    .A2(\lfsr[13] ),
    .B1(_1575_),
    .X(_0166_));
 sky130_fd_sc_hd__inv_2 _5230_ (.A(\lfsr[0] ),
    .Y(_1576_));
 sky130_fd_sc_hd__a21oi_1 _5231_ (.A1(_1576_),
    .A2(\lfsr[14] ),
    .B1(_0920_),
    .Y(_1577_));
 sky130_fd_sc_hd__o21ai_1 _5232_ (.A1(_1576_),
    .A2(\lfsr[14] ),
    .B1(_1577_),
    .Y(_0167_));
 sky130_fd_sc_hd__and2_1 _5233_ (.A(_1562_),
    .B(\lfsr[15] ),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _5234_ (.A(_1578_),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _5235_ (.A(_0920_),
    .B(\lfsr[0] ),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _5236_ (.A(_1579_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _5237_ (.A(_0697_),
    .B(_1270_),
    .Y(_1580_));
 sky130_fd_sc_hd__buf_2 _5238_ (.A(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__nor2_1 _5239_ (.A(_0932_),
    .B(_1281_),
    .Y(_1582_));
 sky130_fd_sc_hd__clkbuf_2 _5240_ (.A(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__or2_1 _5241_ (.A(\as2650.stack[0][0] ),
    .B(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__a21oi_1 _5242_ (.A1(_1520_),
    .A2(_1583_),
    .B1(_1581_),
    .Y(_1585_));
 sky130_fd_sc_hd__a22o_1 _5243_ (.A1(_0634_),
    .A2(_1581_),
    .B1(_1584_),
    .B2(_1585_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _5244_ (.A(\as2650.stack[0][1] ),
    .B(_1583_),
    .X(_1586_));
 sky130_fd_sc_hd__o21a_1 _5245_ (.A1(_0661_),
    .A2(_1282_),
    .B1(_1272_),
    .X(_1587_));
 sky130_fd_sc_hd__a22o_1 _5246_ (.A1(_0659_),
    .A2(_1581_),
    .B1(_1586_),
    .B2(_1587_),
    .X(_0171_));
 sky130_fd_sc_hd__or2_1 _5247_ (.A(\as2650.stack[0][2] ),
    .B(_1583_),
    .X(_1588_));
 sky130_fd_sc_hd__a21oi_1 _5248_ (.A1(_1484_),
    .A2(_1583_),
    .B1(_1581_),
    .Y(_1589_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(_0664_),
    .A2(_1581_),
    .B1(_1588_),
    .B2(_1589_),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(\as2650.stack[0][3] ),
    .B(_1583_),
    .X(_1590_));
 sky130_fd_sc_hd__a21oi_1 _5251_ (.A1(_1487_),
    .A2(_1583_),
    .B1(_1580_),
    .Y(_1591_));
 sky130_fd_sc_hd__a22o_1 _5252_ (.A1(_0667_),
    .A2(_1581_),
    .B1(_1590_),
    .B2(_1591_),
    .X(_0173_));
 sky130_fd_sc_hd__or2_1 _5253_ (.A(\as2650.stack[0][4] ),
    .B(_1583_),
    .X(_1592_));
 sky130_fd_sc_hd__a21oi_1 _5254_ (.A1(_1490_),
    .A2(_1583_),
    .B1(_1580_),
    .Y(_1593_));
 sky130_fd_sc_hd__a22o_1 _5255_ (.A1(_0671_),
    .A2(_1581_),
    .B1(_1592_),
    .B2(_1593_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _5256_ (.A(\as2650.stack[0][5] ),
    .B(_1583_),
    .X(_1594_));
 sky130_fd_sc_hd__o21a_1 _5257_ (.A1(_0676_),
    .A2(_1282_),
    .B1(_1272_),
    .X(_1595_));
 sky130_fd_sc_hd__a22o_1 _5258_ (.A1(_0675_),
    .A2(_1581_),
    .B1(_1594_),
    .B2(_1595_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _5259_ (.A(\as2650.stack[0][6] ),
    .B(_1582_),
    .X(_1596_));
 sky130_fd_sc_hd__o21a_1 _5260_ (.A1(_0681_),
    .A2(_1282_),
    .B1(_1272_),
    .X(_1597_));
 sky130_fd_sc_hd__a22o_1 _5261_ (.A1(_0679_),
    .A2(_1581_),
    .B1(_1596_),
    .B2(_1597_),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _5262_ (.A(\as2650.stack[0][7] ),
    .B(_1582_),
    .X(_1598_));
 sky130_fd_sc_hd__o21a_1 _5263_ (.A1(_0685_),
    .A2(_1282_),
    .B1(_1272_),
    .X(_1599_));
 sky130_fd_sc_hd__a22o_1 _5264_ (.A1(_0684_),
    .A2(_1581_),
    .B1(_1598_),
    .B2(_1599_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _5265_ (.A1(_0983_),
    .A2(_0892_),
    .B1(_3043_),
    .B2(_3155_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_4 _5266_ (.A(_1008_),
    .X(_1601_));
 sky130_fd_sc_hd__nand2_1 _5267_ (.A(_1601_),
    .B(_3103_),
    .Y(_1602_));
 sky130_fd_sc_hd__and3b_1 _5268_ (.A_N(_3053_),
    .B(_3199_),
    .C(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__and3_1 _5269_ (.A(_3112_),
    .B(_3206_),
    .C(_0893_),
    .X(_1604_));
 sky130_fd_sc_hd__nor2_1 _5270_ (.A(\as2650.halted ),
    .B(_3123_),
    .Y(_1605_));
 sky130_fd_sc_hd__or3b_1 _5271_ (.A(_0990_),
    .B(_1604_),
    .C_N(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nor2_4 _5272_ (.A(_3114_),
    .B(_3047_),
    .Y(_1607_));
 sky130_fd_sc_hd__clkbuf_4 _5273_ (.A(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_4 _5274_ (.A(_3156_),
    .X(_1609_));
 sky130_fd_sc_hd__o32a_1 _5275_ (.A1(_1608_),
    .A2(_1609_),
    .A3(_1001_),
    .B1(_1000_),
    .B2(_3160_),
    .X(_1610_));
 sky130_fd_sc_hd__nor2_1 _5276_ (.A(_0900_),
    .B(_0990_),
    .Y(_1611_));
 sky130_fd_sc_hd__a21oi_1 _5277_ (.A1(_0981_),
    .A2(_1611_),
    .B1(_0975_),
    .Y(_1612_));
 sky130_fd_sc_hd__and3b_1 _5278_ (.A_N(_1606_),
    .B(_1610_),
    .C(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__o211a_1 _5279_ (.A1(_3095_),
    .A2(_1009_),
    .B1(_1603_),
    .C1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(io_out[23]),
    .A1(_1600_),
    .S(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _5281_ (.A(_1562_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _5282_ (.A(_1616_),
    .X(_0178_));
 sky130_fd_sc_hd__buf_4 _5283_ (.A(_3227_),
    .X(_1617_));
 sky130_fd_sc_hd__buf_4 _5284_ (.A(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_0759_),
    .B(_1093_),
    .Y(_1619_));
 sky130_fd_sc_hd__or4_1 _5286_ (.A(_1618_),
    .B(_0767_),
    .C(_3197_),
    .D(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(_3067_),
    .A1(io_out[25]),
    .S(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__and2_1 _5288_ (.A(_1562_),
    .B(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _5289_ (.A(_1622_),
    .X(_0179_));
 sky130_fd_sc_hd__a21oi_1 _5290_ (.A1(_0891_),
    .A2(_1019_),
    .B1(_0898_),
    .Y(_1623_));
 sky130_fd_sc_hd__clkbuf_4 _5291_ (.A(_3062_),
    .X(_1624_));
 sky130_fd_sc_hd__or3_1 _5292_ (.A(_3118_),
    .B(_1008_),
    .C(_1001_),
    .X(_1625_));
 sky130_fd_sc_hd__o221a_1 _5293_ (.A1(_0897_),
    .A2(_1003_),
    .B1(_1001_),
    .B2(_0902_),
    .C1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__o221a_1 _5294_ (.A1(_0875_),
    .A2(_0899_),
    .B1(_1623_),
    .B2(_1624_),
    .C1(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__a21boi_1 _5295_ (.A1(_1004_),
    .A2(_1627_),
    .B1_N(io_out[24]),
    .Y(_1628_));
 sky130_fd_sc_hd__buf_4 _5296_ (.A(_0920_),
    .X(_1629_));
 sky130_fd_sc_hd__a311o_1 _5297_ (.A1(_3077_),
    .A2(_1004_),
    .A3(_1627_),
    .B1(_1628_),
    .C1(_1629_),
    .X(_0180_));
 sky130_fd_sc_hd__or4_2 _5298_ (.A(_3120_),
    .B(_0898_),
    .C(_0875_),
    .D(_0877_),
    .X(_1630_));
 sky130_fd_sc_hd__or2_1 _5299_ (.A(_0983_),
    .B(_0897_),
    .X(_1631_));
 sky130_fd_sc_hd__or4b_2 _5300_ (.A(_3158_),
    .B(_3292_),
    .C(_0974_),
    .D_N(_1005_),
    .X(_1632_));
 sky130_fd_sc_hd__o22ai_1 _5301_ (.A1(_0897_),
    .A2(_1630_),
    .B1(_1631_),
    .B2(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__nor3_1 _5302_ (.A(_3066_),
    .B(_3122_),
    .C(_0897_),
    .Y(_1634_));
 sky130_fd_sc_hd__buf_4 _5303_ (.A(_3048_),
    .X(_1635_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_0969_),
    .B(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__or2_1 _5305_ (.A(_3100_),
    .B(_3299_),
    .X(_1637_));
 sky130_fd_sc_hd__nor2_1 _5306_ (.A(_3171_),
    .B(_0913_),
    .Y(_1638_));
 sky130_fd_sc_hd__a31o_1 _5307_ (.A1(_3101_),
    .A2(_3107_),
    .A3(_0912_),
    .B1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__buf_2 _5308_ (.A(_3074_),
    .X(_1640_));
 sky130_fd_sc_hd__nor2_2 _5309_ (.A(_3104_),
    .B(_3158_),
    .Y(_1641_));
 sky130_fd_sc_hd__and4_1 _5310_ (.A(_1640_),
    .B(_1093_),
    .C(_3048_),
    .D(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__nand2_1 _5311_ (.A(_1639_),
    .B(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__o41a_1 _5312_ (.A1(_3121_),
    .A2(_3037_),
    .A3(_1636_),
    .A4(_1637_),
    .B1(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__and3_1 _5313_ (.A(_3178_),
    .B(_3120_),
    .C(_0881_),
    .X(_1645_));
 sky130_fd_sc_hd__a21oi_1 _5314_ (.A1(_3121_),
    .A2(_0884_),
    .B1(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__o21a_1 _5315_ (.A1(_0897_),
    .A2(_3263_),
    .B1(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__o21a_1 _5316_ (.A1(_0876_),
    .A2(_0899_),
    .B1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__or2_1 _5317_ (.A(_3173_),
    .B(_0880_),
    .X(_1649_));
 sky130_fd_sc_hd__nor2_2 _5318_ (.A(_1010_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__nor3_1 _5319_ (.A(_1650_),
    .B(_0997_),
    .C(_0974_),
    .Y(_1651_));
 sky130_fd_sc_hd__or2_2 _5320_ (.A(_3193_),
    .B(_3363_),
    .X(_1652_));
 sky130_fd_sc_hd__nor2_1 _5321_ (.A(_3037_),
    .B(_3043_),
    .Y(_1653_));
 sky130_fd_sc_hd__o221a_1 _5322_ (.A1(_3197_),
    .A2(_0899_),
    .B1(_1003_),
    .B2(_0897_),
    .C1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__o2111a_1 _5323_ (.A1(_3159_),
    .A2(_1651_),
    .B1(_1652_),
    .C1(_1654_),
    .D1(_0654_),
    .X(_1655_));
 sky130_fd_sc_hd__nand3_1 _5324_ (.A(_1644_),
    .B(_1648_),
    .C(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__a21o_1 _5325_ (.A1(_3174_),
    .A2(_3181_),
    .B1(_3159_),
    .X(_1657_));
 sky130_fd_sc_hd__a21oi_1 _5326_ (.A1(_3045_),
    .A2(_3117_),
    .B1(\as2650.halted ),
    .Y(_1658_));
 sky130_fd_sc_hd__and4_1 _5327_ (.A(_3052_),
    .B(_1602_),
    .C(_1657_),
    .D(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__or4b_2 _5328_ (.A(_1633_),
    .B(_1634_),
    .C(_1656_),
    .D_N(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_2 _5329_ (.A(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__or2_2 _5330_ (.A(_3158_),
    .B(_1005_),
    .X(_1662_));
 sky130_fd_sc_hd__nor2_1 _5331_ (.A(_3401_),
    .B(_0406_),
    .Y(_1663_));
 sky130_fd_sc_hd__and4_1 _5332_ (.A(_3288_),
    .B(_0345_),
    .C(_0584_),
    .D(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__and4b_1 _5333_ (.A_N(_0463_),
    .B(_0507_),
    .C(_0621_),
    .D(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__and3_1 _5334_ (.A(_3101_),
    .B(_3067_),
    .C(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__nand2_1 _5335_ (.A(_1642_),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_4 _5336_ (.A(_1662_),
    .B(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__nor2_1 _5337_ (.A(_1661_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__buf_2 _5338_ (.A(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__a21oi_1 _5339_ (.A1(_3254_),
    .A2(_3260_),
    .B1(_1052_),
    .Y(_1671_));
 sky130_fd_sc_hd__a31o_1 _5340_ (.A1(_1052_),
    .A2(_3254_),
    .A3(_3260_),
    .B1(_3091_),
    .X(_1672_));
 sky130_fd_sc_hd__buf_2 _5341_ (.A(_3216_),
    .X(_1673_));
 sky130_fd_sc_hd__and3_1 _5342_ (.A(_3029_),
    .B(_1673_),
    .C(_3250_),
    .X(_1674_));
 sky130_fd_sc_hd__a21oi_1 _5343_ (.A1(_1673_),
    .A2(_3250_),
    .B1(_3029_),
    .Y(_1675_));
 sky130_fd_sc_hd__or2_2 _5344_ (.A(_3088_),
    .B(_3059_),
    .X(_1676_));
 sky130_fd_sc_hd__nor2_2 _5345_ (.A(\as2650.cycle[7] ),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__nor2_4 _5346_ (.A(_3252_),
    .B(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__o21ai_1 _5347_ (.A1(_1674_),
    .A2(_1675_),
    .B1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o21ai_1 _5348_ (.A1(_1671_),
    .A2(_1672_),
    .B1(_1679_),
    .Y(_1680_));
 sky130_fd_sc_hd__clkbuf_4 _5349_ (.A(_3092_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_4 _5350_ (.A(_3061_),
    .X(_1682_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(\as2650.pc[0] ),
    .B(net1),
    .Y(_1683_));
 sky130_fd_sc_hd__or2_1 _5352_ (.A(_0635_),
    .B(_3028_),
    .X(_1684_));
 sky130_fd_sc_hd__and2_1 _5353_ (.A(_1683_),
    .B(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_3049_),
    .B(_3078_),
    .Y(_1686_));
 sky130_fd_sc_hd__clkbuf_4 _5355_ (.A(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__a221o_1 _5356_ (.A1(io_out[8]),
    .A2(_1681_),
    .B1(_1682_),
    .B2(_1685_),
    .C1(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__a21oi_1 _5357_ (.A1(_3060_),
    .A2(_1680_),
    .B1(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__nand2_4 _5358_ (.A(_1617_),
    .B(_3079_),
    .Y(_1690_));
 sky130_fd_sc_hd__and2_1 _5359_ (.A(_3081_),
    .B(_3051_),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_4 _5360_ (.A(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__nor2_2 _5361_ (.A(_1690_),
    .B(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(io_out[8]),
    .B(_0639_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_4 _5363_ (.A(_3151_),
    .B(_1008_),
    .Y(_1695_));
 sky130_fd_sc_hd__clkbuf_4 _5364_ (.A(_3117_),
    .X(_1696_));
 sky130_fd_sc_hd__nor2_2 _5365_ (.A(_0892_),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__o221a_1 _5366_ (.A1(io_out[8]),
    .A2(_1608_),
    .B1(_1695_),
    .B2(_1052_),
    .C1(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__nor2_4 _5367_ (.A(_3081_),
    .B(_3083_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_2 _5368_ (.A(_1696_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(io_out[8]),
    .A1(_1685_),
    .S(_3148_),
    .X(_1701_));
 sky130_fd_sc_hd__o2bb2a_1 _5370_ (.A1_N(_1694_),
    .A2_N(_1698_),
    .B1(_1700_),
    .B2(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__o221a_1 _5371_ (.A1(_0636_),
    .A2(_1693_),
    .B1(_1702_),
    .B2(_1690_),
    .C1(_1018_),
    .X(_1703_));
 sky130_fd_sc_hd__o21a_1 _5372_ (.A1(_1689_),
    .A2(_1703_),
    .B1(_1635_),
    .X(_1704_));
 sky130_fd_sc_hd__nor2_2 _5373_ (.A(_3062_),
    .B(_0975_),
    .Y(_1705_));
 sky130_fd_sc_hd__buf_2 _5374_ (.A(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_2 _5375_ (.A(_1669_),
    .X(_1707_));
 sky130_fd_sc_hd__o21ai_1 _5376_ (.A1(_1520_),
    .A2(_1706_),
    .B1(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__buf_4 _5377_ (.A(_3154_),
    .X(_1709_));
 sky130_fd_sc_hd__o221a_1 _5378_ (.A1(io_out[8]),
    .A2(_1670_),
    .B1(_1704_),
    .B2(_1708_),
    .C1(_1709_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_4 _5379_ (.A(_3252_),
    .X(_1710_));
 sky130_fd_sc_hd__xnor2_1 _5380_ (.A(_1047_),
    .B(_0303_),
    .Y(_1711_));
 sky130_fd_sc_hd__and2_1 _5381_ (.A(net1),
    .B(_3260_),
    .X(_1712_));
 sky130_fd_sc_hd__xor2_1 _5382_ (.A(_1711_),
    .B(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(_3129_),
    .A1(_1713_),
    .S(_3254_),
    .X(_1714_));
 sky130_fd_sc_hd__and2_1 _5384_ (.A(_3128_),
    .B(_0307_),
    .X(_1715_));
 sky130_fd_sc_hd__or2_1 _5385_ (.A(_3128_),
    .B(_0307_),
    .X(_1716_));
 sky130_fd_sc_hd__or2b_1 _5386_ (.A(_1715_),
    .B_N(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__and2_1 _5387_ (.A(net1),
    .B(_3250_),
    .X(_1718_));
 sky130_fd_sc_hd__xnor2_1 _5388_ (.A(_1717_),
    .B(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(_3129_),
    .A1(_1719_),
    .S(_1673_),
    .X(_1720_));
 sky130_fd_sc_hd__a22o_1 _5390_ (.A1(_1710_),
    .A2(_1714_),
    .B1(_1720_),
    .B2(_1678_),
    .X(_1721_));
 sky130_fd_sc_hd__xor2_1 _5391_ (.A(io_out[9]),
    .B(io_out[8]),
    .X(_1722_));
 sky130_fd_sc_hd__and2_1 _5392_ (.A(_0660_),
    .B(_3128_),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_1 _5393_ (.A(_0660_),
    .B(net2),
    .Y(_1724_));
 sky130_fd_sc_hd__nor2_1 _5394_ (.A(_1723_),
    .B(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _5395_ (.A(_1684_),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__or2_1 _5396_ (.A(_1684_),
    .B(_1725_),
    .X(_1727_));
 sky130_fd_sc_hd__and3_1 _5397_ (.A(_3061_),
    .B(_1726_),
    .C(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__a221o_1 _5398_ (.A1(_3060_),
    .A2(_1721_),
    .B1(_1722_),
    .B2(_1681_),
    .C1(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__nor2_1 _5399_ (.A(_0972_),
    .B(_3102_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _5400_ (.A(_3081_),
    .B(_3051_),
    .Y(_1731_));
 sky130_fd_sc_hd__clkbuf_4 _5401_ (.A(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_1730_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_3076_),
    .B(_3085_),
    .Y(_1734_));
 sky130_fd_sc_hd__xnor2_1 _5404_ (.A(_1683_),
    .B(_1725_),
    .Y(_1735_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(io_out[9]),
    .A1(_1735_),
    .S(_3147_),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(io_out[9]),
    .A1(_3129_),
    .S(_3151_),
    .X(_1737_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(_1722_),
    .A1(_1737_),
    .S(_1608_),
    .X(_1738_));
 sky130_fd_sc_hd__a22o_1 _5408_ (.A1(_1734_),
    .A2(_1736_),
    .B1(_1738_),
    .B2(_1697_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_4 _5409_ (.A(_1730_),
    .X(_1740_));
 sky130_fd_sc_hd__a221o_1 _5410_ (.A1(_0660_),
    .A2(_1733_),
    .B1(_1739_),
    .B2(_1740_),
    .C1(_0969_),
    .X(_1741_));
 sky130_fd_sc_hd__o21ai_1 _5411_ (.A1(_1687_),
    .A2(_1729_),
    .B1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a2bb2o_1 _5412_ (.A1_N(_0661_),
    .A2_N(_1706_),
    .B1(_1742_),
    .B2(_1635_),
    .X(_1743_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_1670_),
    .B(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__buf_4 _5414_ (.A(_3154_),
    .X(_1745_));
 sky130_fd_sc_hd__o211a_1 _5415_ (.A1(io_out[9]),
    .A2(_1670_),
    .B1(_1744_),
    .C1(_1745_),
    .X(_0182_));
 sky130_fd_sc_hd__and3_1 _5416_ (.A(io_out[10]),
    .B(io_out[9]),
    .C(io_out[8]),
    .X(_1746_));
 sky130_fd_sc_hd__a21oi_1 _5417_ (.A1(io_out[9]),
    .A2(io_out[8]),
    .B1(io_out[10]),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(_1746_),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__nor2_1 _5419_ (.A(_1676_),
    .B(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(_0660_),
    .B(_3128_),
    .Y(_1750_));
 sky130_fd_sc_hd__nand2_1 _5421_ (.A(\as2650.pc[2] ),
    .B(net3),
    .Y(_1751_));
 sky130_fd_sc_hd__or2_1 _5422_ (.A(\as2650.pc[2] ),
    .B(net3),
    .X(_1752_));
 sky130_fd_sc_hd__nand2_2 _5423_ (.A(_1751_),
    .B(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__a21o_1 _5424_ (.A1(_1750_),
    .A2(_1726_),
    .B1(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__nand3_1 _5425_ (.A(_1750_),
    .B(_1726_),
    .C(_1753_),
    .Y(_1755_));
 sky130_fd_sc_hd__a21o_1 _5426_ (.A1(_1716_),
    .A2(_1718_),
    .B1(_1715_),
    .X(_1756_));
 sky130_fd_sc_hd__or2_1 _5427_ (.A(net3),
    .B(_0340_),
    .X(_1757_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_3131_),
    .B(_0340_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1757_),
    .B(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2_1 _5430_ (.A(_1756_),
    .B(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__a21o_1 _5431_ (.A1(_1756_),
    .A2(_1759_),
    .B1(_3300_),
    .X(_1761_));
 sky130_fd_sc_hd__o22a_1 _5432_ (.A1(_3132_),
    .A2(_1673_),
    .B1(_1760_),
    .B2(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__and2_1 _5433_ (.A(_3128_),
    .B(_0303_),
    .X(_1763_));
 sky130_fd_sc_hd__a21o_1 _5434_ (.A1(_1711_),
    .A2(_1712_),
    .B1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__or2_1 _5435_ (.A(_3131_),
    .B(_0342_),
    .X(_1765_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_3131_),
    .B(_0342_),
    .Y(_1766_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_1765_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__xnor2_1 _5438_ (.A(_1764_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(_3131_),
    .A1(_1768_),
    .S(_3254_),
    .X(_1769_));
 sky130_fd_sc_hd__a22o_1 _5440_ (.A1(_1678_),
    .A2(_1762_),
    .B1(_1769_),
    .B2(_1710_),
    .X(_1770_));
 sky130_fd_sc_hd__a32o_1 _5441_ (.A1(_1682_),
    .A2(_1754_),
    .A3(_1755_),
    .B1(_1770_),
    .B2(_3060_),
    .X(_1771_));
 sky130_fd_sc_hd__buf_4 _5442_ (.A(_0647_),
    .X(_1772_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(_1772_),
    .B(_1748_),
    .Y(_1773_));
 sky130_fd_sc_hd__inv_2 _5444_ (.A(_3151_),
    .Y(_1774_));
 sky130_fd_sc_hd__nand2_2 _5445_ (.A(_1774_),
    .B(_1601_),
    .Y(_1775_));
 sky130_fd_sc_hd__o22a_1 _5446_ (.A1(io_out[10]),
    .A2(_1775_),
    .B1(_1695_),
    .B2(_3132_),
    .X(_1776_));
 sky130_fd_sc_hd__o21a_1 _5447_ (.A1(_1683_),
    .A2(_1724_),
    .B1(_1750_),
    .X(_1777_));
 sky130_fd_sc_hd__xnor2_2 _5448_ (.A(_1753_),
    .B(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(_3148_),
    .B(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__o211a_1 _5450_ (.A1(io_out[10]),
    .A2(_3148_),
    .B1(_1734_),
    .C1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__a31o_1 _5451_ (.A1(_1697_),
    .A2(_1773_),
    .A3(_1776_),
    .B1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__a221o_1 _5452_ (.A1(\as2650.pc[2] ),
    .A2(_1733_),
    .B1(_1781_),
    .B2(_1740_),
    .C1(_0970_),
    .X(_1782_));
 sky130_fd_sc_hd__o31a_1 _5453_ (.A1(_1687_),
    .A2(_1749_),
    .A3(_1771_),
    .B1(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__o22a_1 _5454_ (.A1(\as2650.pc[2] ),
    .A2(_1706_),
    .B1(_1783_),
    .B2(_1624_),
    .X(_1784_));
 sky130_fd_sc_hd__or2_1 _5455_ (.A(io_out[10]),
    .B(_1707_),
    .X(_1785_));
 sky130_fd_sc_hd__buf_4 _5456_ (.A(_3154_),
    .X(_1786_));
 sky130_fd_sc_hd__o311a_1 _5457_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_1784_),
    .B1(_1785_),
    .C1(_1786_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_0767_),
    .B(_1732_),
    .Y(_1787_));
 sky130_fd_sc_hd__or2_1 _5459_ (.A(_0668_),
    .B(_3134_),
    .X(_1788_));
 sky130_fd_sc_hd__nand2_2 _5460_ (.A(\as2650.pc[3] ),
    .B(_3134_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(_1788_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__o21a_1 _5462_ (.A1(_1753_),
    .A2(_1777_),
    .B1(_1751_),
    .X(_1791_));
 sky130_fd_sc_hd__xor2_1 _5463_ (.A(_1790_),
    .B(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(io_out[11]),
    .A1(_1792_),
    .S(_3147_),
    .X(_1793_));
 sky130_fd_sc_hd__and2_1 _5465_ (.A(io_out[11]),
    .B(_1746_),
    .X(_1794_));
 sky130_fd_sc_hd__nor2_1 _5466_ (.A(io_out[11]),
    .B(_1746_),
    .Y(_1795_));
 sky130_fd_sc_hd__or2_1 _5467_ (.A(_1794_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o21ai_1 _5468_ (.A1(_1608_),
    .A2(_1796_),
    .B1(_1697_),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_4 _5469_ (.A(_1774_),
    .B(_3097_),
    .Y(_1798_));
 sky130_fd_sc_hd__a22o_1 _5470_ (.A1(io_out[11]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(_3135_),
    .X(_1799_));
 sky130_fd_sc_hd__or2_1 _5471_ (.A(_1797_),
    .B(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__o21a_1 _5472_ (.A1(_1700_),
    .A2(_1793_),
    .B1(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o2bb2a_1 _5473_ (.A1_N(_1487_),
    .A2_N(_1787_),
    .B1(_1801_),
    .B2(_0907_),
    .X(_1802_));
 sky130_fd_sc_hd__buf_4 _5474_ (.A(_3103_),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_4 _5475_ (.A(\as2650.cycle[7] ),
    .B(_1681_),
    .Y(_1804_));
 sky130_fd_sc_hd__a221o_1 _5476_ (.A1(net3),
    .A2(_0342_),
    .B1(_1711_),
    .B2(_1712_),
    .C1(_1763_),
    .X(_1805_));
 sky130_fd_sc_hd__nor2_1 _5477_ (.A(_3134_),
    .B(_0420_),
    .Y(_1806_));
 sky130_fd_sc_hd__and2_1 _5478_ (.A(_3134_),
    .B(_0420_),
    .X(_1807_));
 sky130_fd_sc_hd__nor2_1 _5479_ (.A(_1806_),
    .B(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__a21oi_1 _5480_ (.A1(_1765_),
    .A2(_1805_),
    .B1(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__a31o_1 _5481_ (.A1(_1765_),
    .A2(_1808_),
    .A3(_1805_),
    .B1(_3212_),
    .X(_1810_));
 sky130_fd_sc_hd__a2bb2o_1 _5482_ (.A1_N(_1809_),
    .A2_N(_1810_),
    .B1(_3135_),
    .B2(_3212_),
    .X(_1811_));
 sky130_fd_sc_hd__a221o_1 _5483_ (.A1(net3),
    .A2(_0340_),
    .B1(_1716_),
    .B2(_1718_),
    .C1(_1715_),
    .X(_1812_));
 sky130_fd_sc_hd__nor2_1 _5484_ (.A(_3134_),
    .B(_0403_),
    .Y(_1813_));
 sky130_fd_sc_hd__and2_1 _5485_ (.A(_3134_),
    .B(_0403_),
    .X(_1814_));
 sky130_fd_sc_hd__nor2_1 _5486_ (.A(_1813_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__a21oi_1 _5487_ (.A1(_1757_),
    .A2(_1812_),
    .B1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__a31o_1 _5488_ (.A1(_1757_),
    .A2(_1815_),
    .A3(_1812_),
    .B1(_3300_),
    .X(_1817_));
 sky130_fd_sc_hd__o22a_1 _5489_ (.A1(_0818_),
    .A2(_1673_),
    .B1(_1816_),
    .B2(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__a2bb2o_1 _5490_ (.A1_N(_3090_),
    .A2_N(_1811_),
    .B1(_1818_),
    .B2(_1678_),
    .X(_1819_));
 sky130_fd_sc_hd__a221o_1 _5491_ (.A1(_1681_),
    .A2(_1796_),
    .B1(_1804_),
    .B2(_1819_),
    .C1(_1682_),
    .X(_1820_));
 sky130_fd_sc_hd__nand2_1 _5492_ (.A(_1751_),
    .B(_1754_),
    .Y(_1821_));
 sky130_fd_sc_hd__or2_1 _5493_ (.A(\as2650.cycle[6] ),
    .B(_3060_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_4 _5494_ (.A(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__a31o_1 _5495_ (.A1(_1788_),
    .A2(_1789_),
    .A3(_1821_),
    .B1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__a31o_1 _5496_ (.A1(_1751_),
    .A2(_1754_),
    .A3(_1790_),
    .B1(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__nand3_1 _5497_ (.A(_1803_),
    .B(_1820_),
    .C(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__o221a_1 _5498_ (.A1(_0668_),
    .A2(_0898_),
    .B1(_1802_),
    .B2(_1098_),
    .C1(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__o22a_1 _5499_ (.A1(_0668_),
    .A2(_1706_),
    .B1(_1827_),
    .B2(_1624_),
    .X(_1828_));
 sky130_fd_sc_hd__or2_1 _5500_ (.A(io_out[11]),
    .B(_1707_),
    .X(_1829_));
 sky130_fd_sc_hd__o311a_1 _5501_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_1828_),
    .B1(_1829_),
    .C1(_1786_),
    .X(_0184_));
 sky130_fd_sc_hd__xnor2_1 _5502_ (.A(_0465_),
    .B(_0480_),
    .Y(_1830_));
 sky130_fd_sc_hd__or2_1 _5503_ (.A(_3134_),
    .B(_0403_),
    .X(_1831_));
 sky130_fd_sc_hd__a31o_1 _5504_ (.A1(_1757_),
    .A2(_1831_),
    .A3(_1812_),
    .B1(_1814_),
    .X(_1832_));
 sky130_fd_sc_hd__xnor2_1 _5505_ (.A(_1830_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(_0465_),
    .A1(_1833_),
    .S(_1673_),
    .X(_1834_));
 sky130_fd_sc_hd__xnor2_1 _5507_ (.A(net5),
    .B(_0477_),
    .Y(_1835_));
 sky130_fd_sc_hd__or2_1 _5508_ (.A(_3134_),
    .B(_0420_),
    .X(_1836_));
 sky130_fd_sc_hd__a31oi_2 _5509_ (.A1(_1765_),
    .A2(_1836_),
    .A3(_1805_),
    .B1(_1807_),
    .Y(_1837_));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(_1835_),
    .B(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(_3137_),
    .A1(_1838_),
    .S(_3254_),
    .X(_1839_));
 sky130_fd_sc_hd__a2bb2o_1 _5512_ (.A1_N(_3094_),
    .A2_N(_1834_),
    .B1(_1839_),
    .B2(_1710_),
    .X(_1840_));
 sky130_fd_sc_hd__nand2_1 _5513_ (.A(_1788_),
    .B(_1821_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(\as2650.pc[4] ),
    .B(net5),
    .Y(_1842_));
 sky130_fd_sc_hd__or2_1 _5515_ (.A(\as2650.pc[4] ),
    .B(net5),
    .X(_1843_));
 sky130_fd_sc_hd__nand2_1 _5516_ (.A(_1842_),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__a21oi_2 _5517_ (.A1(_1789_),
    .A2(_1841_),
    .B1(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__a31o_1 _5518_ (.A1(_1789_),
    .A2(_1844_),
    .A3(_1841_),
    .B1(_1823_),
    .X(_1846_));
 sky130_fd_sc_hd__xnor2_1 _5519_ (.A(io_out[12]),
    .B(_1794_),
    .Y(_1847_));
 sky130_fd_sc_hd__o21a_1 _5520_ (.A1(_1676_),
    .A2(_1847_),
    .B1(_3103_),
    .X(_1848_));
 sky130_fd_sc_hd__o21ai_1 _5521_ (.A1(_1845_),
    .A2(_1846_),
    .B1(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__a21o_1 _5522_ (.A1(_3060_),
    .A2(_1840_),
    .B1(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__a21o_1 _5523_ (.A1(_1487_),
    .A2(_0818_),
    .B1(_1791_),
    .X(_1851_));
 sky130_fd_sc_hd__a21o_1 _5524_ (.A1(_1789_),
    .A2(_1851_),
    .B1(_1844_),
    .X(_1852_));
 sky130_fd_sc_hd__nand3_1 _5525_ (.A(_1789_),
    .B(_1844_),
    .C(_1851_),
    .Y(_1853_));
 sky130_fd_sc_hd__nand2_1 _5526_ (.A(_1852_),
    .B(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _5527_ (.A(_3148_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__or2_1 _5528_ (.A(io_out[12]),
    .B(_3148_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_4 _5529_ (.A(_3326_),
    .X(_1857_));
 sky130_fd_sc_hd__o2bb2a_1 _5530_ (.A1_N(_1857_),
    .A2_N(_1847_),
    .B1(_1775_),
    .B2(io_out[12]),
    .X(_1858_));
 sky130_fd_sc_hd__o211a_1 _5531_ (.A1(_3137_),
    .A2(_1695_),
    .B1(_1858_),
    .C1(_1697_),
    .X(_1859_));
 sky130_fd_sc_hd__a31o_1 _5532_ (.A1(_1734_),
    .A2(_1855_),
    .A3(_1856_),
    .B1(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__a221o_1 _5533_ (.A1(_0672_),
    .A2(_1787_),
    .B1(_1860_),
    .B2(_0767_),
    .C1(_1098_),
    .X(_1861_));
 sky130_fd_sc_hd__o211a_1 _5534_ (.A1(_0672_),
    .A2(_0898_),
    .B1(_1850_),
    .C1(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__o22a_1 _5535_ (.A1(_0672_),
    .A2(_1706_),
    .B1(_1862_),
    .B2(_1624_),
    .X(_1863_));
 sky130_fd_sc_hd__or2_1 _5536_ (.A(io_out[12]),
    .B(_1707_),
    .X(_1864_));
 sky130_fd_sc_hd__o311a_1 _5537_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_1863_),
    .B1(_1864_),
    .C1(_1786_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_4 _5538_ (.A(_1601_),
    .X(_1865_));
 sky130_fd_sc_hd__and3_1 _5539_ (.A(io_out[13]),
    .B(io_out[12]),
    .C(_1794_),
    .X(_1866_));
 sky130_fd_sc_hd__a21oi_1 _5540_ (.A1(io_out[12]),
    .A2(_1794_),
    .B1(io_out[13]),
    .Y(_1867_));
 sky130_fd_sc_hd__or2_1 _5541_ (.A(_1866_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nor2_1 _5542_ (.A(_1865_),
    .B(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__a221o_1 _5543_ (.A1(io_out[13]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(_3140_),
    .C1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__nor2_2 _5544_ (.A(_0972_),
    .B(_3117_),
    .Y(_1871_));
 sky130_fd_sc_hd__nand2_2 _5545_ (.A(_3119_),
    .B(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__o22a_1 _5546_ (.A1(\as2650.pc[5] ),
    .A2(_1693_),
    .B1(_1870_),
    .B2(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(\as2650.pc[5] ),
    .B(net6),
    .Y(_1874_));
 sky130_fd_sc_hd__or2_1 _5548_ (.A(\as2650.pc[5] ),
    .B(net6),
    .X(_1875_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(_1874_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(_1842_),
    .B(_1852_),
    .Y(_1877_));
 sky130_fd_sc_hd__xnor2_1 _5551_ (.A(_1876_),
    .B(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__and2_1 _5552_ (.A(io_out[13]),
    .B(_1091_),
    .X(_1879_));
 sky130_fd_sc_hd__a2111o_1 _5553_ (.A1(_3150_),
    .A2(_1878_),
    .B1(_1879_),
    .C1(_1700_),
    .D1(_1690_),
    .X(_1880_));
 sky130_fd_sc_hd__nand2_2 _5554_ (.A(_3101_),
    .B(_1635_),
    .Y(_1881_));
 sky130_fd_sc_hd__clkbuf_4 _5555_ (.A(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__a21oi_1 _5556_ (.A1(_1873_),
    .A2(_1880_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__a21o_1 _5557_ (.A1(_0672_),
    .A2(_3137_),
    .B1(_1845_),
    .X(_1884_));
 sky130_fd_sc_hd__xor2_1 _5558_ (.A(_1876_),
    .B(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__and2_1 _5559_ (.A(net5),
    .B(_0480_),
    .X(_1886_));
 sky130_fd_sc_hd__a21oi_1 _5560_ (.A1(_1830_),
    .A2(_1832_),
    .B1(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__or2_1 _5561_ (.A(_3139_),
    .B(_0499_),
    .X(_1888_));
 sky130_fd_sc_hd__nand2_1 _5562_ (.A(_3139_),
    .B(_0499_),
    .Y(_1889_));
 sky130_fd_sc_hd__nand2_1 _5563_ (.A(_1888_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__xnor2_1 _5564_ (.A(_1887_),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(_1046_),
    .A1(_1891_),
    .S(_1673_),
    .X(_1892_));
 sky130_fd_sc_hd__and2_1 _5566_ (.A(_3139_),
    .B(_0516_),
    .X(_1893_));
 sky130_fd_sc_hd__or2_1 _5567_ (.A(_3139_),
    .B(_0516_),
    .X(_1894_));
 sky130_fd_sc_hd__and2b_1 _5568_ (.A_N(_1893_),
    .B(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(net5),
    .B(_0477_),
    .Y(_1896_));
 sky130_fd_sc_hd__o21ai_1 _5570_ (.A1(_1835_),
    .A2(_1837_),
    .B1(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__xnor2_1 _5571_ (.A(_1895_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(_1046_),
    .A1(_1898_),
    .S(_3254_),
    .X(_1899_));
 sky130_fd_sc_hd__a22o_1 _5573_ (.A1(_1678_),
    .A2(_1892_),
    .B1(_1899_),
    .B2(_1710_),
    .X(_1900_));
 sky130_fd_sc_hd__a221o_1 _5574_ (.A1(_1804_),
    .A2(_1900_),
    .B1(_1868_),
    .B2(_1681_),
    .C1(_3061_),
    .X(_1901_));
 sky130_fd_sc_hd__o211a_1 _5575_ (.A1(_1823_),
    .A2(_1885_),
    .B1(_1901_),
    .C1(_1803_),
    .X(_1902_));
 sky130_fd_sc_hd__a2bb2o_1 _5576_ (.A1_N(_0676_),
    .A2_N(_1705_),
    .B1(_1902_),
    .B2(_1635_),
    .X(_1903_));
 sky130_fd_sc_hd__o21ai_1 _5577_ (.A1(_1883_),
    .A2(_1903_),
    .B1(_1670_),
    .Y(_1904_));
 sky130_fd_sc_hd__o211a_1 _5578_ (.A1(io_out[13]),
    .A2(_1670_),
    .B1(_1904_),
    .C1(_1745_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _5579_ (.A(\as2650.pc[6] ),
    .B(net7),
    .X(_1905_));
 sky130_fd_sc_hd__nor2_1 _5580_ (.A(_0680_),
    .B(net7),
    .Y(_1906_));
 sky130_fd_sc_hd__nor2_2 _5581_ (.A(_1905_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_1 _5582_ (.A(_1842_),
    .B(_1874_),
    .Y(_1908_));
 sky130_fd_sc_hd__o21a_1 _5583_ (.A1(_1845_),
    .A2(_1908_),
    .B1(_1875_),
    .X(_1909_));
 sky130_fd_sc_hd__xor2_1 _5584_ (.A(_1907_),
    .B(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__and2_1 _5585_ (.A(io_out[14]),
    .B(_1866_),
    .X(_1911_));
 sky130_fd_sc_hd__nor2_1 _5586_ (.A(io_out[14]),
    .B(_1866_),
    .Y(_1912_));
 sky130_fd_sc_hd__or2_1 _5587_ (.A(_1911_),
    .B(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__o21ai_1 _5588_ (.A1(_1676_),
    .A2(_1913_),
    .B1(_3103_),
    .Y(_1914_));
 sky130_fd_sc_hd__and2_1 _5589_ (.A(_3143_),
    .B(_0577_),
    .X(_1915_));
 sky130_fd_sc_hd__or2_1 _5590_ (.A(_3143_),
    .B(_0577_),
    .X(_1916_));
 sky130_fd_sc_hd__or2b_1 _5591_ (.A(_1915_),
    .B_N(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__a221o_1 _5592_ (.A1(_3139_),
    .A2(_0499_),
    .B1(_1830_),
    .B2(_1832_),
    .C1(_1886_),
    .X(_1918_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_1888_),
    .B(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__xor2_1 _5594_ (.A(_1917_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__nand2_1 _5595_ (.A(_1022_),
    .B(_3300_),
    .Y(_1921_));
 sky130_fd_sc_hd__o211a_1 _5596_ (.A1(_3300_),
    .A2(_1920_),
    .B1(_1921_),
    .C1(_1678_),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(_3143_),
    .B(_0579_),
    .Y(_1923_));
 sky130_fd_sc_hd__or2_1 _5598_ (.A(_3143_),
    .B(_0579_),
    .X(_1924_));
 sky130_fd_sc_hd__nand2_1 _5599_ (.A(_1923_),
    .B(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__a21o_2 _5600_ (.A1(_1894_),
    .A2(_1897_),
    .B1(_1893_),
    .X(_1926_));
 sky130_fd_sc_hd__xnor2_1 _5601_ (.A(_1925_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_1022_),
    .B(_3212_),
    .Y(_1928_));
 sky130_fd_sc_hd__o211a_1 _5603_ (.A1(_3212_),
    .A2(_1927_),
    .B1(_1928_),
    .C1(_1710_),
    .X(_1929_));
 sky130_fd_sc_hd__o21a_1 _5604_ (.A1(_1922_),
    .A2(_1929_),
    .B1(_3060_),
    .X(_1930_));
 sky130_fd_sc_hd__a211o_1 _5605_ (.A1(_1682_),
    .A2(_1910_),
    .B1(_1914_),
    .C1(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_1772_),
    .B(_1913_),
    .Y(_1932_));
 sky130_fd_sc_hd__o221a_1 _5607_ (.A1(io_out[14]),
    .A2(_1775_),
    .B1(_1695_),
    .B2(_3144_),
    .C1(_1697_),
    .X(_1933_));
 sky130_fd_sc_hd__a21bo_1 _5608_ (.A1(_1875_),
    .A2(_1877_),
    .B1_N(_1874_),
    .X(_1934_));
 sky130_fd_sc_hd__xor2_2 _5609_ (.A(_1907_),
    .B(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(io_out[14]),
    .A1(_1935_),
    .S(_3148_),
    .X(_1936_));
 sky130_fd_sc_hd__a22o_1 _5611_ (.A1(_1932_),
    .A2(_1933_),
    .B1(_1936_),
    .B2(_1734_),
    .X(_1937_));
 sky130_fd_sc_hd__a221o_1 _5612_ (.A1(_0680_),
    .A2(_1733_),
    .B1(_1937_),
    .B2(_1740_),
    .C1(_0970_),
    .X(_1938_));
 sky130_fd_sc_hd__a21oi_1 _5613_ (.A1(_1931_),
    .A2(_1938_),
    .B1(_1624_),
    .Y(_1939_));
 sky130_fd_sc_hd__nor2_1 _5614_ (.A(_0681_),
    .B(_1706_),
    .Y(_1940_));
 sky130_fd_sc_hd__o21ai_1 _5615_ (.A1(_1939_),
    .A2(_1940_),
    .B1(_1707_),
    .Y(_1941_));
 sky130_fd_sc_hd__o211a_1 _5616_ (.A1(io_out[14]),
    .A2(_1670_),
    .B1(_1941_),
    .C1(_1745_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _5617_ (.A(io_out[15]),
    .B(_1911_),
    .Y(_1942_));
 sky130_fd_sc_hd__nor2_1 _5618_ (.A(_1865_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__a221o_1 _5619_ (.A1(io_out[15]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(_3148_),
    .C1(_1872_),
    .X(_1944_));
 sky130_fd_sc_hd__o22a_1 _5620_ (.A1(\as2650.pc[7] ),
    .A2(_1693_),
    .B1(_1943_),
    .B2(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__and2_1 _5621_ (.A(\as2650.pc[7] ),
    .B(net7),
    .X(_1946_));
 sky130_fd_sc_hd__nor2_1 _5622_ (.A(\as2650.pc[7] ),
    .B(_3142_),
    .Y(_1947_));
 sky130_fd_sc_hd__nor2_2 _5623_ (.A(_1946_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__a21oi_1 _5624_ (.A1(_1907_),
    .A2(_1934_),
    .B1(_1905_),
    .Y(_1949_));
 sky130_fd_sc_hd__xnor2_2 _5625_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__a211o_1 _5626_ (.A1(_3149_),
    .A2(_1950_),
    .B1(_1700_),
    .C1(_0691_),
    .X(_1951_));
 sky130_fd_sc_hd__a211o_1 _5627_ (.A1(io_out[15]),
    .A2(_1091_),
    .B1(_1098_),
    .C1(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__a21o_1 _5628_ (.A1(_1907_),
    .A2(_1909_),
    .B1(_1905_),
    .X(_1953_));
 sky130_fd_sc_hd__xnor2_1 _5629_ (.A(_1948_),
    .B(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__inv_2 _5630_ (.A(_1923_),
    .Y(_1955_));
 sky130_fd_sc_hd__a21oi_1 _5631_ (.A1(_1924_),
    .A2(_1926_),
    .B1(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__xnor2_1 _5632_ (.A(_3147_),
    .B(_0628_),
    .Y(_1957_));
 sky130_fd_sc_hd__a21oi_1 _5633_ (.A1(_1956_),
    .A2(_1957_),
    .B1(_3212_),
    .Y(_1958_));
 sky130_fd_sc_hd__o21ai_1 _5634_ (.A1(_1956_),
    .A2(_1957_),
    .B1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(_3148_),
    .B(_3212_),
    .Y(_1960_));
 sky130_fd_sc_hd__a31o_1 _5636_ (.A1(_1888_),
    .A2(_1916_),
    .A3(_1918_),
    .B1(_1915_),
    .X(_1961_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(_3146_),
    .B(_0616_),
    .X(_1962_));
 sky130_fd_sc_hd__or2_1 _5638_ (.A(_3146_),
    .B(_0616_),
    .X(_1963_));
 sky130_fd_sc_hd__and2b_1 _5639_ (.A_N(_1962_),
    .B(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__nand2_1 _5640_ (.A(_1961_),
    .B(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__o21a_1 _5641_ (.A1(_1961_),
    .A2(_1964_),
    .B1(_1673_),
    .X(_1966_));
 sky130_fd_sc_hd__o2bb2a_1 _5642_ (.A1_N(_1965_),
    .A2_N(_1966_),
    .B1(_1091_),
    .B2(_1673_),
    .X(_1967_));
 sky130_fd_sc_hd__a32o_1 _5643_ (.A1(_1710_),
    .A2(_1959_),
    .A3(_1960_),
    .B1(_1678_),
    .B2(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__a221o_1 _5644_ (.A1(_1804_),
    .A2(_1968_),
    .B1(_1942_),
    .B2(_1681_),
    .C1(_3061_),
    .X(_1969_));
 sky130_fd_sc_hd__o211ai_1 _5645_ (.A1(_1823_),
    .A2(_1954_),
    .B1(_1969_),
    .C1(_1803_),
    .Y(_1970_));
 sky130_fd_sc_hd__o211a_1 _5646_ (.A1(_0970_),
    .A2(_1945_),
    .B1(_1952_),
    .C1(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__o22a_1 _5647_ (.A1(_0685_),
    .A2(_1706_),
    .B1(_1971_),
    .B2(_1624_),
    .X(_1972_));
 sky130_fd_sc_hd__or2_1 _5648_ (.A(io_out[15]),
    .B(_1707_),
    .X(_1973_));
 sky130_fd_sc_hd__o311a_1 _5649_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_1972_),
    .B1(_1973_),
    .C1(_1786_),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _5650_ (.A(_1804_),
    .Y(_1974_));
 sky130_fd_sc_hd__a221oi_4 _5651_ (.A1(_3146_),
    .A2(_0628_),
    .B1(_1924_),
    .B2(_1926_),
    .C1(_1955_),
    .Y(_1975_));
 sky130_fd_sc_hd__o21ai_1 _5652_ (.A1(_3146_),
    .A2(_0628_),
    .B1(_3254_),
    .Y(_1976_));
 sky130_fd_sc_hd__or2_1 _5653_ (.A(_1975_),
    .B(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__xnor2_1 _5654_ (.A(_3030_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__a311o_1 _5655_ (.A1(_1888_),
    .A2(_1916_),
    .A3(_1918_),
    .B1(_1962_),
    .C1(_1915_),
    .X(_1979_));
 sky130_fd_sc_hd__and2_1 _5656_ (.A(_3216_),
    .B(_1963_),
    .X(_1980_));
 sky130_fd_sc_hd__nand2_1 _5657_ (.A(_1979_),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__xnor2_1 _5658_ (.A(_3030_),
    .B(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__o22a_1 _5659_ (.A1(_3090_),
    .A2(_1978_),
    .B1(_1982_),
    .B2(_3094_),
    .X(_1983_));
 sky130_fd_sc_hd__and3_1 _5660_ (.A(io_out[16]),
    .B(io_out[15]),
    .C(_1911_),
    .X(_1984_));
 sky130_fd_sc_hd__a21oi_1 _5661_ (.A1(io_out[15]),
    .A2(_1911_),
    .B1(io_out[16]),
    .Y(_1985_));
 sky130_fd_sc_hd__nor2_1 _5662_ (.A(_1984_),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__o221a_1 _5663_ (.A1(_1974_),
    .A2(_1983_),
    .B1(_1986_),
    .B2(_1676_),
    .C1(_1823_),
    .X(_1987_));
 sky130_fd_sc_hd__nand2_1 _5664_ (.A(\as2650.pc[8] ),
    .B(_3142_),
    .Y(_1988_));
 sky130_fd_sc_hd__or2_1 _5665_ (.A(\as2650.pc[8] ),
    .B(_3142_),
    .X(_1989_));
 sky130_fd_sc_hd__and2_1 _5666_ (.A(_1988_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__or4b_1 _5667_ (.A(_1876_),
    .B(_1905_),
    .C(_1906_),
    .D_N(_1948_),
    .X(_1991_));
 sky130_fd_sc_hd__inv_2 _5668_ (.A(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__a41o_1 _5669_ (.A1(_1875_),
    .A2(_1907_),
    .A3(_1908_),
    .A4(_1948_),
    .B1(_1905_),
    .X(_1993_));
 sky130_fd_sc_hd__or2_1 _5670_ (.A(_1946_),
    .B(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__a21o_1 _5671_ (.A1(_1845_),
    .A2(_1992_),
    .B1(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__nand2_1 _5672_ (.A(_1990_),
    .B(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__or2_1 _5673_ (.A(_1990_),
    .B(_1995_),
    .X(_1997_));
 sky130_fd_sc_hd__and3_1 _5674_ (.A(_1682_),
    .B(_1996_),
    .C(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__or4_1 _5675_ (.A(_1687_),
    .B(_3062_),
    .C(_1987_),
    .D(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__o21ba_1 _5676_ (.A1(_1852_),
    .A2(_1991_),
    .B1_N(_1994_),
    .X(_2000_));
 sky130_fd_sc_hd__xor2_1 _5677_ (.A(_1990_),
    .B(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__nor2_1 _5678_ (.A(_1700_),
    .B(_1690_),
    .Y(_2002_));
 sky130_fd_sc_hd__o21ai_1 _5679_ (.A1(io_out[16]),
    .A2(_3149_),
    .B1(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__a21o_1 _5680_ (.A1(_3150_),
    .A2(_2001_),
    .B1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__inv_2 _5681_ (.A(_0689_),
    .Y(_2005_));
 sky130_fd_sc_hd__o22a_1 _5682_ (.A1(io_out[16]),
    .A2(_1775_),
    .B1(_1695_),
    .B2(_3030_),
    .X(_2006_));
 sky130_fd_sc_hd__o21ai_1 _5683_ (.A1(_1608_),
    .A2(_1986_),
    .B1(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__nor2_4 _5684_ (.A(_0969_),
    .B(_3062_),
    .Y(_2008_));
 sky130_fd_sc_hd__o221a_1 _5685_ (.A1(_2005_),
    .A2(_1693_),
    .B1(_1872_),
    .B2(_2007_),
    .C1(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__o2bb2a_1 _5686_ (.A1_N(_2004_),
    .A2_N(_2009_),
    .B1(_0689_),
    .B2(_1705_),
    .X(_2010_));
 sky130_fd_sc_hd__a21bo_1 _5687_ (.A1(_1999_),
    .A2(_2010_),
    .B1_N(_1707_),
    .X(_2011_));
 sky130_fd_sc_hd__o211a_1 _5688_ (.A1(io_out[16]),
    .A2(_1670_),
    .B1(_2011_),
    .C1(_1745_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _5689_ (.A(io_out[17]),
    .B(_1984_),
    .X(_2012_));
 sky130_fd_sc_hd__nor2_1 _5690_ (.A(io_out[17]),
    .B(_1984_),
    .Y(_2013_));
 sky130_fd_sc_hd__or2_1 _5691_ (.A(_2012_),
    .B(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__inv_2 _5692_ (.A(\as2650.addr_buff[0] ),
    .Y(_2015_));
 sky130_fd_sc_hd__inv_2 _5693_ (.A(\as2650.addr_buff[1] ),
    .Y(_2016_));
 sky130_fd_sc_hd__o21a_1 _5694_ (.A1(_2015_),
    .A2(_1977_),
    .B1(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__nor2_1 _5695_ (.A(_2015_),
    .B(_2016_),
    .Y(_2018_));
 sky130_fd_sc_hd__or3b_1 _5696_ (.A(_1975_),
    .B(_1976_),
    .C_N(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__nand2_1 _5697_ (.A(_3252_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__o31a_1 _5698_ (.A1(_2015_),
    .A2(_2016_),
    .A3(_1981_),
    .B1(_1678_),
    .X(_2021_));
 sky130_fd_sc_hd__a31o_1 _5699_ (.A1(_3030_),
    .A2(_1979_),
    .A3(_1980_),
    .B1(\as2650.addr_buff[1] ),
    .X(_2022_));
 sky130_fd_sc_hd__a2bb2o_1 _5700_ (.A1_N(_2017_),
    .A2_N(_2020_),
    .B1(_2021_),
    .B2(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a2bb2o_1 _5701_ (.A1_N(_1676_),
    .A2_N(_2014_),
    .B1(_2023_),
    .B2(_1804_),
    .X(_2024_));
 sky130_fd_sc_hd__xnor2_2 _5702_ (.A(\as2650.pc[9] ),
    .B(_3142_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _5703_ (.A(_1988_),
    .B(_1996_),
    .Y(_2026_));
 sky130_fd_sc_hd__xnor2_1 _5704_ (.A(_2025_),
    .B(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(_2024_),
    .A1(_2027_),
    .S(_1682_),
    .X(_2028_));
 sky130_fd_sc_hd__nor2_1 _5706_ (.A(_1865_),
    .B(_2014_),
    .Y(_2029_));
 sky130_fd_sc_hd__a221o_1 _5707_ (.A1(io_out[17]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(\as2650.addr_buff[1] ),
    .C1(_1872_),
    .X(_2030_));
 sky130_fd_sc_hd__o22a_1 _5708_ (.A1(_0704_),
    .A2(_1693_),
    .B1(_2029_),
    .B2(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or2_1 _5709_ (.A(_0969_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__or2b_1 _5710_ (.A(_2000_),
    .B_N(_1990_),
    .X(_2033_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_1988_),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__xnor2_1 _5712_ (.A(_2025_),
    .B(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__a211o_1 _5713_ (.A1(_3149_),
    .A2(_2035_),
    .B1(_1700_),
    .C1(_0907_),
    .X(_2036_));
 sky130_fd_sc_hd__a211o_1 _5714_ (.A1(io_out[17]),
    .A2(_1091_),
    .B1(_1098_),
    .C1(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__o211a_1 _5715_ (.A1(_1687_),
    .A2(_2028_),
    .B1(_2032_),
    .C1(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__o22a_1 _5716_ (.A1(_0704_),
    .A2(_1706_),
    .B1(_2038_),
    .B2(_1624_),
    .X(_2039_));
 sky130_fd_sc_hd__or2_1 _5717_ (.A(io_out[17]),
    .B(_1707_),
    .X(_2040_));
 sky130_fd_sc_hd__o311a_1 _5718_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_2039_),
    .B1(_2040_),
    .C1(_1786_),
    .X(_0190_));
 sky130_fd_sc_hd__o21ai_1 _5719_ (.A1(_0704_),
    .A2(_0689_),
    .B1(_3143_),
    .Y(_2041_));
 sky130_fd_sc_hd__or2_1 _5720_ (.A(_1996_),
    .B(_2025_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(\as2650.pc[10] ),
    .B(_3143_),
    .Y(_2043_));
 sky130_fd_sc_hd__or2_1 _5722_ (.A(\as2650.pc[10] ),
    .B(_3142_),
    .X(_2044_));
 sky130_fd_sc_hd__nand2_2 _5723_ (.A(_2043_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__a21oi_1 _5724_ (.A1(_2041_),
    .A2(_2042_),
    .B1(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__a31o_1 _5725_ (.A1(_2045_),
    .A2(_2041_),
    .A3(_2042_),
    .B1(_1823_),
    .X(_2047_));
 sky130_fd_sc_hd__a21oi_1 _5726_ (.A1(_1710_),
    .A2(_2019_),
    .B1(_2021_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand3_1 _5727_ (.A(_1678_),
    .B(_1979_),
    .C(_1980_),
    .Y(_2049_));
 sky130_fd_sc_hd__o31ai_2 _5728_ (.A1(_3090_),
    .A2(_1975_),
    .A3(_1976_),
    .B1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__and3_1 _5729_ (.A(\as2650.addr_buff[0] ),
    .B(\as2650.addr_buff[1] ),
    .C(\as2650.addr_buff[2] ),
    .X(_2051_));
 sky130_fd_sc_hd__a2bb2o_1 _5730_ (.A1_N(\as2650.addr_buff[2] ),
    .A2_N(_2048_),
    .B1(_2050_),
    .B2(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__xnor2_1 _5731_ (.A(io_out[18]),
    .B(_2012_),
    .Y(_2053_));
 sky130_fd_sc_hd__a221o_1 _5732_ (.A1(_1804_),
    .A2(_2052_),
    .B1(_2053_),
    .B2(_1681_),
    .C1(_1682_),
    .X(_2054_));
 sky130_fd_sc_hd__o2111a_1 _5733_ (.A1(_2046_),
    .A2(_2047_),
    .B1(_1803_),
    .C1(_1635_),
    .D1(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__inv_2 _5734_ (.A(_2045_),
    .Y(_2056_));
 sky130_fd_sc_hd__or2_1 _5735_ (.A(_2033_),
    .B(_2025_),
    .X(_2057_));
 sky130_fd_sc_hd__nand2_1 _5736_ (.A(_2041_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__xnor2_1 _5737_ (.A(_2056_),
    .B(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_3150_),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__o211a_1 _5739_ (.A1(io_out[18]),
    .A2(_3150_),
    .B1(_2002_),
    .C1(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(_1772_),
    .B(_2053_),
    .Y(_2062_));
 sky130_fd_sc_hd__o221a_1 _5741_ (.A1(io_out[18]),
    .A2(_1775_),
    .B1(_1695_),
    .B2(\as2650.addr_buff[2] ),
    .C1(_0891_),
    .X(_2063_));
 sky130_fd_sc_hd__a22o_1 _5742_ (.A1(_0713_),
    .A2(_1692_),
    .B1(_2062_),
    .B2(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__a221o_1 _5743_ (.A1(_0713_),
    .A2(_1690_),
    .B1(_2064_),
    .B2(_1871_),
    .C1(_1881_),
    .X(_2065_));
 sky130_fd_sc_hd__o22ai_1 _5744_ (.A1(_0713_),
    .A2(_1706_),
    .B1(_2061_),
    .B2(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__o21ai_1 _5745_ (.A1(_2055_),
    .A2(_2066_),
    .B1(_1707_),
    .Y(_2067_));
 sky130_fd_sc_hd__o211a_1 _5746_ (.A1(io_out[18]),
    .A2(_1670_),
    .B1(_2067_),
    .C1(_1745_),
    .X(_0191_));
 sky130_fd_sc_hd__xor2_1 _5747_ (.A(\as2650.pc[11] ),
    .B(_3142_),
    .X(_2068_));
 sky130_fd_sc_hd__inv_2 _5748_ (.A(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__a21bo_1 _5749_ (.A1(_2056_),
    .A2(_2058_),
    .B1_N(_2043_),
    .X(_2070_));
 sky130_fd_sc_hd__xnor2_1 _5750_ (.A(_2069_),
    .B(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(io_out[19]),
    .A1(_2071_),
    .S(_3147_),
    .X(_2072_));
 sky130_fd_sc_hd__and3_1 _5752_ (.A(io_out[19]),
    .B(io_out[18]),
    .C(_2012_),
    .X(_2073_));
 sky130_fd_sc_hd__a21oi_1 _5753_ (.A1(io_out[18]),
    .A2(_2012_),
    .B1(io_out[19]),
    .Y(_2074_));
 sky130_fd_sc_hd__or2_1 _5754_ (.A(_2073_),
    .B(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__nor2_1 _5755_ (.A(_1601_),
    .B(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__a221o_1 _5756_ (.A1(io_out[19]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(\as2650.addr_buff[3] ),
    .C1(_1609_),
    .X(_2077_));
 sky130_fd_sc_hd__o22a_1 _5757_ (.A1(_0719_),
    .A2(_1732_),
    .B1(_2076_),
    .B2(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__o32a_1 _5758_ (.A1(_0691_),
    .A2(_1700_),
    .A3(_2072_),
    .B1(_2078_),
    .B2(_1696_),
    .X(_2079_));
 sky130_fd_sc_hd__o22a_1 _5759_ (.A1(_0719_),
    .A2(_1740_),
    .B1(_2079_),
    .B2(_0972_),
    .X(_2080_));
 sky130_fd_sc_hd__nor2_1 _5760_ (.A(\as2650.addr_buff[2] ),
    .B(_1677_),
    .Y(_2081_));
 sky130_fd_sc_hd__a2111o_1 _5761_ (.A1(_3252_),
    .A2(_2019_),
    .B1(_2081_),
    .C1(_2021_),
    .D1(\as2650.addr_buff[3] ),
    .X(_2082_));
 sky130_fd_sc_hd__a21bo_1 _5762_ (.A1(_2050_),
    .A2(_2051_),
    .B1_N(\as2650.addr_buff[3] ),
    .X(_2083_));
 sky130_fd_sc_hd__a32o_1 _5763_ (.A1(_1804_),
    .A2(_2082_),
    .A3(_2083_),
    .B1(_2075_),
    .B2(_1681_),
    .X(_2084_));
 sky130_fd_sc_hd__a21oi_1 _5764_ (.A1(_0713_),
    .A2(_3144_),
    .B1(_2046_),
    .Y(_2085_));
 sky130_fd_sc_hd__xnor2_1 _5765_ (.A(_2069_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(_2084_),
    .A1(_2086_),
    .S(_3061_),
    .X(_2087_));
 sky130_fd_sc_hd__a2bb2o_1 _5767_ (.A1_N(_0970_),
    .A2_N(_2080_),
    .B1(_2087_),
    .B2(_3103_),
    .X(_2088_));
 sky130_fd_sc_hd__a2bb2o_1 _5768_ (.A1_N(_0719_),
    .A2_N(_1705_),
    .B1(_2088_),
    .B2(_1635_),
    .X(_2089_));
 sky130_fd_sc_hd__nand2_1 _5769_ (.A(_1670_),
    .B(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__o211a_1 _5770_ (.A1(io_out[19]),
    .A2(_1670_),
    .B1(_2090_),
    .C1(_1745_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _5771_ (.A(\as2650.addr_buff[4] ),
    .Y(_2091_));
 sky130_fd_sc_hd__a31o_1 _5772_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2050_),
    .A3(_2051_),
    .B1(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__nand2_1 _5773_ (.A(\as2650.addr_buff[2] ),
    .B(\as2650.addr_buff[3] ),
    .Y(_2093_));
 sky130_fd_sc_hd__inv_2 _5774_ (.A(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__o211ai_1 _5775_ (.A1(_1677_),
    .A2(_2094_),
    .B1(_2048_),
    .C1(_2091_),
    .Y(_2095_));
 sky130_fd_sc_hd__xnor2_1 _5776_ (.A(io_out[20]),
    .B(_2073_),
    .Y(_2096_));
 sky130_fd_sc_hd__a32o_1 _5777_ (.A1(_1804_),
    .A2(_2092_),
    .A3(_2095_),
    .B1(_2096_),
    .B2(_1681_),
    .X(_2097_));
 sky130_fd_sc_hd__xor2_2 _5778_ (.A(\as2650.pc[12] ),
    .B(_3143_),
    .X(_2098_));
 sky130_fd_sc_hd__o41a_1 _5779_ (.A1(\as2650.pc[11] ),
    .A2(\as2650.pc[10] ),
    .A3(_0704_),
    .A4(\as2650.pc[8] ),
    .B1(_3143_),
    .X(_2099_));
 sky130_fd_sc_hd__inv_2 _5780_ (.A(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__o31a_1 _5781_ (.A1(_2045_),
    .A2(_2042_),
    .A3(_2069_),
    .B1(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__xnor2_1 _5782_ (.A(_2098_),
    .B(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(_1682_),
    .B(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__o21ai_1 _5784_ (.A1(_1682_),
    .A2(_2097_),
    .B1(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__o31a_1 _5785_ (.A1(_2045_),
    .A2(_2057_),
    .A3(_2069_),
    .B1(_2100_),
    .X(_2105_));
 sky130_fd_sc_hd__xnor2_1 _5786_ (.A(_2098_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(io_out[20]),
    .A1(_2106_),
    .S(_3147_),
    .X(_2107_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(_1601_),
    .B(_2096_),
    .Y(_2108_));
 sky130_fd_sc_hd__a221o_1 _5789_ (.A1(io_out[20]),
    .A2(_0639_),
    .B1(_1798_),
    .B2(\as2650.addr_buff[4] ),
    .C1(_1609_),
    .X(_2109_));
 sky130_fd_sc_hd__o22a_1 _5790_ (.A1(_0726_),
    .A2(_1732_),
    .B1(_2108_),
    .B2(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__o32a_1 _5791_ (.A1(_0887_),
    .A2(_1700_),
    .A3(_2107_),
    .B1(_2110_),
    .B2(_1696_),
    .X(_2111_));
 sky130_fd_sc_hd__o22a_1 _5792_ (.A1(_0726_),
    .A2(_1740_),
    .B1(_2111_),
    .B2(_0972_),
    .X(_2112_));
 sky130_fd_sc_hd__o22a_1 _5793_ (.A1(_1687_),
    .A2(_2104_),
    .B1(_2112_),
    .B2(_0970_),
    .X(_2113_));
 sky130_fd_sc_hd__o22a_1 _5794_ (.A1(_0726_),
    .A2(_1706_),
    .B1(_2113_),
    .B2(_1624_),
    .X(_2114_));
 sky130_fd_sc_hd__or2_1 _5795_ (.A(io_out[20]),
    .B(_1707_),
    .X(_2115_));
 sky130_fd_sc_hd__o311a_1 _5796_ (.A1(_1661_),
    .A2(_1668_),
    .A3(_2114_),
    .B1(_2115_),
    .C1(_1786_),
    .X(_0193_));
 sky130_fd_sc_hd__a211o_1 _5797_ (.A1(io_oeb),
    .A2(_3205_),
    .B1(_0638_),
    .C1(_0887_),
    .X(_2116_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_0969_),
    .B(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__o21ai_1 _5799_ (.A1(_3160_),
    .A2(_1000_),
    .B1(_0981_),
    .Y(_2118_));
 sky130_fd_sc_hd__a31o_1 _5800_ (.A1(io_out[21]),
    .A2(_3330_),
    .A3(_1019_),
    .B1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__buf_2 _5801_ (.A(_0641_),
    .X(_2120_));
 sky130_fd_sc_hd__a31o_1 _5802_ (.A1(io_out[21]),
    .A2(_2120_),
    .A3(_3080_),
    .B1(_1098_),
    .X(_2121_));
 sky130_fd_sc_hd__and4_1 _5803_ (.A(_1635_),
    .B(_2117_),
    .C(_2119_),
    .D(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__and3b_1 _5804_ (.A_N(_1633_),
    .B(_1647_),
    .C(_0654_),
    .X(_2123_));
 sky130_fd_sc_hd__nor2_1 _5805_ (.A(_3093_),
    .B(_1687_),
    .Y(_2124_));
 sky130_fd_sc_hd__and3_1 _5806_ (.A(_3146_),
    .B(_3061_),
    .C(_3063_),
    .X(_2125_));
 sky130_fd_sc_hd__or2_1 _5807_ (.A(_2124_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(_3039_),
    .B(_3090_),
    .Y(_2127_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_3151_),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__o31a_1 _5810_ (.A1(_3146_),
    .A2(_0902_),
    .A3(_3076_),
    .B1(_1093_),
    .X(_2129_));
 sky130_fd_sc_hd__o2111a_1 _5811_ (.A1(_0983_),
    .A2(_1804_),
    .B1(_2128_),
    .C1(_2129_),
    .D1(_1626_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _5812_ (.A(_3227_),
    .B(_1640_),
    .Y(_2131_));
 sky130_fd_sc_hd__or4_1 _5813_ (.A(_3121_),
    .B(_3037_),
    .C(_1881_),
    .D(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__and4b_1 _5814_ (.A_N(_2126_),
    .B(_2130_),
    .C(_2132_),
    .D(_1652_),
    .X(_2133_));
 sky130_fd_sc_hd__o2bb2a_1 _5815_ (.A1_N(_0969_),
    .A2_N(_3112_),
    .B1(_0876_),
    .B2(_0899_),
    .X(_2134_));
 sky130_fd_sc_hd__o211a_1 _5816_ (.A1(_3159_),
    .A2(_1651_),
    .B1(_2134_),
    .C1(_1662_),
    .X(_2135_));
 sky130_fd_sc_hd__and4_1 _5817_ (.A(_1644_),
    .B(_1659_),
    .C(_2133_),
    .D(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__and3_1 _5818_ (.A(_1667_),
    .B(_2123_),
    .C(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(io_out[21]),
    .A1(_2122_),
    .S(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__and2_1 _5820_ (.A(_3154_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_1 _5821_ (.A(_2139_),
    .X(_0194_));
 sky130_fd_sc_hd__and3_1 _5822_ (.A(_3146_),
    .B(_1699_),
    .C(_1871_),
    .X(_2140_));
 sky130_fd_sc_hd__a31o_1 _5823_ (.A1(_1640_),
    .A2(_1730_),
    .A3(_1692_),
    .B1(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__o21a_1 _5824_ (.A1(_0997_),
    .A2(_0974_),
    .B1(_0887_),
    .X(_2142_));
 sky130_fd_sc_hd__nor2_2 _5825_ (.A(_3051_),
    .B(_0646_),
    .Y(_2143_));
 sky130_fd_sc_hd__nor2_1 _5826_ (.A(_3158_),
    .B(_3174_),
    .Y(_2144_));
 sky130_fd_sc_hd__inv_2 _5827_ (.A(_1658_),
    .Y(_2145_));
 sky130_fd_sc_hd__a311o_1 _5828_ (.A1(_3046_),
    .A2(_2143_),
    .A3(_3115_),
    .B1(_2144_),
    .C1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__and3_1 _5829_ (.A(_3123_),
    .B(_3045_),
    .C(_3076_),
    .X(_2147_));
 sky130_fd_sc_hd__o21a_1 _5830_ (.A1(_3114_),
    .A2(_3077_),
    .B1(_0641_),
    .X(_2148_));
 sky130_fd_sc_hd__and3b_1 _5831_ (.A_N(_3115_),
    .B(_2147_),
    .C(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__or3b_1 _5832_ (.A(_2146_),
    .B(_2149_),
    .C_N(_1652_),
    .X(_2150_));
 sky130_fd_sc_hd__o31a_1 _5833_ (.A1(_1010_),
    .A2(_3160_),
    .A3(_1649_),
    .B1(_0654_),
    .X(_2151_));
 sky130_fd_sc_hd__or3b_1 _5834_ (.A(_2142_),
    .B(_2150_),
    .C_N(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__o221a_1 _5835_ (.A1(_3160_),
    .A2(_0760_),
    .B1(_1732_),
    .B2(_1640_),
    .C1(_1626_),
    .X(_2153_));
 sky130_fd_sc_hd__o211a_1 _5836_ (.A1(_1631_),
    .A2(_1632_),
    .B1(_1643_),
    .C1(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_1648_),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__a211o_1 _5838_ (.A1(_1018_),
    .A2(_2141_),
    .B1(_2152_),
    .C1(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__nor2_1 _5839_ (.A(_1668_),
    .B(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__clkbuf_4 _5840_ (.A(_0646_),
    .X(_2158_));
 sky130_fd_sc_hd__nor2_1 _5841_ (.A(_1608_),
    .B(_0638_),
    .Y(_2159_));
 sky130_fd_sc_hd__a21o_1 _5842_ (.A1(_2158_),
    .A2(_2159_),
    .B1(_1798_),
    .X(_2160_));
 sky130_fd_sc_hd__a32o_1 _5843_ (.A1(io_out[22]),
    .A2(_1697_),
    .A3(_2160_),
    .B1(_3149_),
    .B2(_1696_),
    .X(_2161_));
 sky130_fd_sc_hd__a311o_1 _5844_ (.A1(io_out[22]),
    .A2(_0973_),
    .A3(_1000_),
    .B1(_0691_),
    .C1(_1617_),
    .X(_2162_));
 sky130_fd_sc_hd__o21ai_1 _5845_ (.A1(_1690_),
    .A2(_2161_),
    .B1(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_1018_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__a31o_1 _5847_ (.A1(io_out[22]),
    .A2(_0973_),
    .A3(_2159_),
    .B1(_1687_),
    .X(_2165_));
 sky130_fd_sc_hd__a31o_1 _5848_ (.A1(_1093_),
    .A2(_2164_),
    .A3(_2165_),
    .B1(_1624_),
    .X(_2166_));
 sky130_fd_sc_hd__or3_1 _5849_ (.A(_1668_),
    .B(_2156_),
    .C(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__o211a_1 _5850_ (.A1(io_out[22]),
    .A2(_2157_),
    .B1(_2167_),
    .C1(_1745_),
    .X(_0195_));
 sky130_fd_sc_hd__or3_1 _5851_ (.A(_3121_),
    .B(_3099_),
    .C(_3037_),
    .X(_2168_));
 sky130_fd_sc_hd__or3_1 _5852_ (.A(_0897_),
    .B(_0975_),
    .C(_2127_),
    .X(_2169_));
 sky130_fd_sc_hd__or3b_2 _5853_ (.A(_0890_),
    .B(_2168_),
    .C_N(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__a21oi_1 _5854_ (.A1(\as2650.addr_buff[5] ),
    .A2(_1635_),
    .B1(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__a211oi_1 _5855_ (.A1(_3247_),
    .A2(_2170_),
    .B1(_2171_),
    .C1(_0921_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21oi_1 _5856_ (.A1(\as2650.addr_buff[6] ),
    .A2(_1635_),
    .B1(_2170_),
    .Y(_2172_));
 sky130_fd_sc_hd__a211oi_1 _5857_ (.A1(_3245_),
    .A2(_2170_),
    .B1(_2172_),
    .C1(_0921_),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(_3262_),
    .A1(_3029_),
    .S(_3080_),
    .X(_2173_));
 sky130_fd_sc_hd__a31o_1 _5859_ (.A1(_0690_),
    .A2(_3202_),
    .A3(_0963_),
    .B1(_3209_),
    .X(_2174_));
 sky130_fd_sc_hd__a21o_1 _5860_ (.A1(_0973_),
    .A2(_1012_),
    .B1(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__nor2_1 _5861_ (.A(_3293_),
    .B(_1632_),
    .Y(_2176_));
 sky130_fd_sc_hd__or3_1 _5862_ (.A(_0976_),
    .B(_2175_),
    .C(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__clkbuf_4 _5863_ (.A(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(_2173_),
    .A1(\as2650.holding_reg[0] ),
    .S(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__clkbuf_1 _5865_ (.A(_2179_),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_1047_),
    .B(_3079_),
    .Y(_2180_));
 sky130_fd_sc_hd__or2_1 _5867_ (.A(_3391_),
    .B(_0767_),
    .X(_2181_));
 sky130_fd_sc_hd__and2_1 _5868_ (.A(_2180_),
    .B(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(_2182_),
    .A1(\as2650.holding_reg[1] ),
    .S(_2178_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _5870_ (.A(_2183_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(_0326_),
    .A1(_3132_),
    .S(_3080_),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(_2184_),
    .A1(\as2650.holding_reg[2] ),
    .S(_2178_),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _5873_ (.A(_2185_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _5874_ (.A(_0417_),
    .B(_0907_),
    .Y(_2186_));
 sky130_fd_sc_hd__o21a_1 _5875_ (.A1(_0818_),
    .A2(_0889_),
    .B1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__inv_2 _5876_ (.A(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(_2188_),
    .A1(\as2650.holding_reg[3] ),
    .S(_2178_),
    .X(_2189_));
 sky130_fd_sc_hd__clkbuf_1 _5878_ (.A(_2189_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_0470_),
    .B(_0907_),
    .Y(_2190_));
 sky130_fd_sc_hd__o21a_1 _5880_ (.A1(_0465_),
    .A2(_0889_),
    .B1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__inv_2 _5881_ (.A(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(_2192_),
    .A1(\as2650.holding_reg[4] ),
    .S(_2178_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_1 _5883_ (.A(_2193_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(_0513_),
    .A1(_3140_),
    .S(_3080_),
    .X(_2194_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(_2194_),
    .A1(\as2650.holding_reg[5] ),
    .S(_2178_),
    .X(_2195_));
 sky130_fd_sc_hd__clkbuf_1 _5886_ (.A(_2195_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5887_ (.A0(_0545_),
    .A1(_3144_),
    .S(_0767_),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(_2196_),
    .A1(\as2650.holding_reg[6] ),
    .S(_2178_),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _5889_ (.A(_2197_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5890_ (.A0(_0618_),
    .A1(_3150_),
    .S(_0767_),
    .X(_2198_));
 sky130_fd_sc_hd__mux2_1 _5891_ (.A0(_2198_),
    .A1(\as2650.holding_reg[7] ),
    .S(_2178_),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _5892_ (.A(_2199_),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _5893_ (.A1(_0769_),
    .A2(_1006_),
    .B1(_1629_),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _5894_ (.A(_1631_),
    .Y(_2200_));
 sky130_fd_sc_hd__nor2_1 _5895_ (.A(_3251_),
    .B(_3205_),
    .Y(_2201_));
 sky130_fd_sc_hd__a21o_1 _5896_ (.A1(_3151_),
    .A2(_3252_),
    .B1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__a21oi_1 _5897_ (.A1(_1091_),
    .A2(_3205_),
    .B1(_1823_),
    .Y(_2203_));
 sky130_fd_sc_hd__a211o_1 _5898_ (.A1(_3046_),
    .A2(_3251_),
    .B1(_2202_),
    .C1(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__or4_1 _5899_ (.A(_1608_),
    .B(_0907_),
    .C(_1604_),
    .D(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_0889_),
    .B(_0893_),
    .Y(_2206_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_3155_),
    .B(_3119_),
    .Y(_2207_));
 sky130_fd_sc_hd__or2_4 _5902_ (.A(_1639_),
    .B(_1666_),
    .X(_2208_));
 sky130_fd_sc_hd__or2_1 _5903_ (.A(_3159_),
    .B(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__o211a_1 _5904_ (.A1(_3115_),
    .A2(_2207_),
    .B1(_2209_),
    .C1(_1640_),
    .X(_2210_));
 sky130_fd_sc_hd__a211o_1 _5905_ (.A1(_3155_),
    .A2(_3114_),
    .B1(_1798_),
    .C1(_2158_),
    .X(_2211_));
 sky130_fd_sc_hd__and3b_1 _5906_ (.A_N(_2210_),
    .B(_2211_),
    .C(_1618_),
    .X(_2212_));
 sky130_fd_sc_hd__or4_1 _5907_ (.A(_3046_),
    .B(_0990_),
    .C(_0878_),
    .D(_0882_),
    .X(_2213_));
 sky130_fd_sc_hd__or2_1 _5908_ (.A(_0879_),
    .B(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__a2bb2o_1 _5909_ (.A1_N(_1857_),
    .A2_N(_1000_),
    .B1(_2207_),
    .B2(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__o211ai_1 _5910_ (.A1(_0891_),
    .A2(_0913_),
    .B1(_0990_),
    .C1(_3155_),
    .Y(_2216_));
 sky130_fd_sc_hd__a21oi_1 _5911_ (.A1(_2215_),
    .A2(_2216_),
    .B1(_1618_),
    .Y(_2217_));
 sky130_fd_sc_hd__clkbuf_4 _5912_ (.A(_3076_),
    .X(_2218_));
 sky130_fd_sc_hd__o32ai_1 _5913_ (.A1(_0897_),
    .A2(_2212_),
    .A3(_2217_),
    .B1(_2218_),
    .B2(_3155_),
    .Y(_2219_));
 sky130_fd_sc_hd__a32o_1 _5914_ (.A1(_2200_),
    .A2(_2205_),
    .A3(_2206_),
    .B1(_2219_),
    .B2(_1018_),
    .X(_2220_));
 sky130_fd_sc_hd__o22a_1 _5915_ (.A1(_0769_),
    .A2(_3155_),
    .B1(_1619_),
    .B2(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__nor2_1 _5916_ (.A(_1629_),
    .B(_2221_),
    .Y(_0207_));
 sky130_fd_sc_hd__o21ai_1 _5917_ (.A1(_0641_),
    .A2(_0638_),
    .B1(_1617_),
    .Y(_2222_));
 sky130_fd_sc_hd__a211oi_1 _5918_ (.A1(_0891_),
    .A2(_2222_),
    .B1(_2148_),
    .C1(_1696_),
    .Y(_2223_));
 sky130_fd_sc_hd__xnor2_1 _5919_ (.A(_3040_),
    .B(_3046_),
    .Y(_2224_));
 sky130_fd_sc_hd__and3_1 _5920_ (.A(_3155_),
    .B(_1609_),
    .C(_0913_),
    .X(_2225_));
 sky130_fd_sc_hd__nor2_2 _5921_ (.A(_1617_),
    .B(_0874_),
    .Y(_2226_));
 sky130_fd_sc_hd__a211oi_1 _5922_ (.A1(_2225_),
    .A2(_2226_),
    .B1(_0969_),
    .C1(_0897_),
    .Y(_2227_));
 sky130_fd_sc_hd__o221a_1 _5923_ (.A1(_3193_),
    .A2(_2214_),
    .B1(_2223_),
    .B2(_2224_),
    .C1(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__o21a_1 _5924_ (.A1(_2131_),
    .A2(_2209_),
    .B1(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__o21a_1 _5925_ (.A1(_2224_),
    .A2(_2202_),
    .B1(_1823_),
    .X(_2230_));
 sky130_fd_sc_hd__or4_1 _5926_ (.A(_0907_),
    .B(_0638_),
    .C(_2203_),
    .D(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__a311o_1 _5927_ (.A1(_2200_),
    .A2(_2206_),
    .A3(_2231_),
    .B1(_1624_),
    .C1(_0890_),
    .X(_2232_));
 sky130_fd_sc_hd__o2bb2a_1 _5928_ (.A1_N(_0890_),
    .A2_N(_3040_),
    .B1(_2229_),
    .B2(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__nor2_1 _5929_ (.A(_1629_),
    .B(_2233_),
    .Y(_0208_));
 sky130_fd_sc_hd__and3_1 _5930_ (.A(_3034_),
    .B(_3040_),
    .C(_3046_),
    .X(_2234_));
 sky130_fd_sc_hd__a21oi_1 _5931_ (.A1(_3040_),
    .A2(_3046_),
    .B1(_3034_),
    .Y(_2235_));
 sky130_fd_sc_hd__nor3_1 _5932_ (.A(_1865_),
    .B(_2234_),
    .C(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__or4_1 _5933_ (.A(_3292_),
    .B(_3206_),
    .C(_0963_),
    .D(_1012_),
    .X(_2237_));
 sky130_fd_sc_hd__or2b_1 _5934_ (.A(_2236_),
    .B_N(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__a211o_1 _5935_ (.A1(_0892_),
    .A2(_0988_),
    .B1(_2234_),
    .C1(_2235_),
    .X(_2239_));
 sky130_fd_sc_hd__a31o_1 _5936_ (.A1(_3068_),
    .A2(_3098_),
    .A3(_0900_),
    .B1(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__nand3b_1 _5937_ (.A_N(_1000_),
    .B(_2239_),
    .C(_3098_),
    .Y(_2241_));
 sky130_fd_sc_hd__o2111ai_1 _5938_ (.A1(_3050_),
    .A2(_0874_),
    .B1(_2240_),
    .C1(_2241_),
    .D1(_0972_),
    .Y(_2242_));
 sky130_fd_sc_hd__o311a_1 _5939_ (.A1(_2158_),
    .A2(_3114_),
    .A3(_3077_),
    .B1(_3085_),
    .C1(_2236_),
    .X(_2243_));
 sky130_fd_sc_hd__nor2_1 _5940_ (.A(_2158_),
    .B(_1695_),
    .Y(_2244_));
 sky130_fd_sc_hd__o21ai_1 _5941_ (.A1(_3057_),
    .A2(_2218_),
    .B1(_1618_),
    .Y(_2245_));
 sky130_fd_sc_hd__o31a_1 _5942_ (.A1(_2243_),
    .A2(_2244_),
    .A3(_2245_),
    .B1(_2008_),
    .X(_2246_));
 sky130_fd_sc_hd__a221o_1 _5943_ (.A1(_3063_),
    .A2(_2238_),
    .B1(_2242_),
    .B2(_2246_),
    .C1(_0890_),
    .X(_2247_));
 sky130_fd_sc_hd__o211a_1 _5944_ (.A1(_0769_),
    .A2(_3034_),
    .B1(_1786_),
    .C1(_2247_),
    .X(_0209_));
 sky130_fd_sc_hd__o21ai_1 _5945_ (.A1(_3110_),
    .A2(_2159_),
    .B1(_3085_),
    .Y(_2248_));
 sky130_fd_sc_hd__nor2_1 _5946_ (.A(_3033_),
    .B(_2234_),
    .Y(_2249_));
 sky130_fd_sc_hd__and2_1 _5947_ (.A(_3033_),
    .B(_2234_),
    .X(_2250_));
 sky130_fd_sc_hd__or2_1 _5948_ (.A(_2249_),
    .B(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__a211oi_1 _5949_ (.A1(_1618_),
    .A2(_2248_),
    .B1(_2251_),
    .C1(_0970_),
    .Y(_2252_));
 sky130_fd_sc_hd__a32o_1 _5950_ (.A1(_3050_),
    .A2(_1640_),
    .A3(_1798_),
    .B1(_1699_),
    .B2(_3150_),
    .X(_2253_));
 sky130_fd_sc_hd__o211a_1 _5951_ (.A1(_3205_),
    .A2(_3214_),
    .B1(_2251_),
    .C1(_3091_),
    .X(_2254_));
 sky130_fd_sc_hd__o21a_1 _5952_ (.A1(_3151_),
    .A2(_3205_),
    .B1(_1710_),
    .X(_2255_));
 sky130_fd_sc_hd__o22a_1 _5953_ (.A1(_1823_),
    .A2(_3205_),
    .B1(_2254_),
    .B2(_2255_),
    .X(_2256_));
 sky130_fd_sc_hd__a2111o_1 _5954_ (.A1(_3150_),
    .A2(_1682_),
    .B1(_0638_),
    .C1(_1604_),
    .D1(_1018_),
    .X(_2257_));
 sky130_fd_sc_hd__nor2_1 _5955_ (.A(_2256_),
    .B(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__a211o_1 _5956_ (.A1(_3123_),
    .A2(_2253_),
    .B1(_2258_),
    .C1(_0890_),
    .X(_2259_));
 sky130_fd_sc_hd__o221a_1 _5957_ (.A1(_0769_),
    .A2(_3033_),
    .B1(_2252_),
    .B2(_2259_),
    .C1(_1709_),
    .X(_0210_));
 sky130_fd_sc_hd__a21oi_1 _5958_ (.A1(_0769_),
    .A2(_2250_),
    .B1(\as2650.cycle[4] ),
    .Y(_2260_));
 sky130_fd_sc_hd__and3_1 _5959_ (.A(_0769_),
    .B(\as2650.cycle[4] ),
    .C(_2250_),
    .X(_2261_));
 sky130_fd_sc_hd__nor3_1 _5960_ (.A(_1629_),
    .B(_2260_),
    .C(_2261_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _5961_ (.A1(\as2650.cycle[5] ),
    .A2(_2261_),
    .B1(_0921_),
    .Y(_2262_));
 sky130_fd_sc_hd__o21a_1 _5962_ (.A1(\as2650.cycle[5] ),
    .A2(_2261_),
    .B1(_2262_),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _5963_ (.A(\as2650.cycle[5] ),
    .B(\as2650.cycle[4] ),
    .C(_2250_),
    .X(_2263_));
 sky130_fd_sc_hd__and2_1 _5964_ (.A(\as2650.cycle[6] ),
    .B(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__or2_1 _5965_ (.A(\as2650.cycle[6] ),
    .B(_2263_),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_1774_),
    .B(_1710_),
    .Y(_2266_));
 sky130_fd_sc_hd__a31o_1 _5967_ (.A1(_1823_),
    .A2(_2266_),
    .A3(_3214_),
    .B1(_1636_),
    .X(_2267_));
 sky130_fd_sc_hd__and3b_1 _5968_ (.A_N(_2264_),
    .B(_2265_),
    .C(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__a311o_1 _5969_ (.A1(_3081_),
    .A2(_3063_),
    .A3(_1641_),
    .B1(_2125_),
    .C1(_0890_),
    .X(_2269_));
 sky130_fd_sc_hd__o221a_1 _5970_ (.A1(_0769_),
    .A2(\as2650.cycle[6] ),
    .B1(_2268_),
    .B2(_2269_),
    .C1(_1709_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_4 _5971_ (.A(_0975_),
    .X(_2270_));
 sky130_fd_sc_hd__xnor2_1 _5972_ (.A(\as2650.cycle[7] ),
    .B(_2264_),
    .Y(_2271_));
 sky130_fd_sc_hd__or4b_1 _5973_ (.A(_2270_),
    .B(_2271_),
    .C(_2127_),
    .D_N(_3064_),
    .X(_2272_));
 sky130_fd_sc_hd__a21oi_1 _5974_ (.A1(_1618_),
    .A2(_2270_),
    .B1(_0890_),
    .Y(_2273_));
 sky130_fd_sc_hd__a221oi_1 _5975_ (.A1(_0890_),
    .A2(_3058_),
    .B1(_2272_),
    .B2(_2273_),
    .C1(_0921_),
    .Y(_0214_));
 sky130_fd_sc_hd__mux2_1 _5976_ (.A0(\as2650.psu[7] ),
    .A1(_0916_),
    .S(_3150_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(_0978_),
    .B(_1011_),
    .Y(_2275_));
 sky130_fd_sc_hd__o22a_1 _5978_ (.A1(_0618_),
    .A2(_0978_),
    .B1(_2275_),
    .B2(\as2650.sense ),
    .X(_2276_));
 sky130_fd_sc_hd__o21a_1 _5979_ (.A1(_1011_),
    .A2(_2274_),
    .B1(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__or2_1 _5980_ (.A(\as2650.psu[7] ),
    .B(_0769_),
    .X(_2278_));
 sky130_fd_sc_hd__o211a_1 _5981_ (.A1(_0890_),
    .A2(_2277_),
    .B1(_2278_),
    .C1(_1745_),
    .X(_0215_));
 sky130_fd_sc_hd__a21o_1 _5982_ (.A1(_2159_),
    .A2(_2168_),
    .B1(_1636_),
    .X(_2279_));
 sky130_fd_sc_hd__and3_1 _5983_ (.A(_1640_),
    .B(_3112_),
    .C(_1730_),
    .X(_2280_));
 sky130_fd_sc_hd__a31o_1 _5984_ (.A1(_1617_),
    .A2(_1640_),
    .A3(_1798_),
    .B1(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__a21oi_1 _5985_ (.A1(_3123_),
    .A2(_2281_),
    .B1(_2150_),
    .Y(_2282_));
 sky130_fd_sc_hd__o311a_1 _5986_ (.A1(_3058_),
    .A2(\as2650.cycle[6] ),
    .A3(_0983_),
    .B1(_1093_),
    .C1(_3052_),
    .X(_2283_));
 sky130_fd_sc_hd__or4_1 _5987_ (.A(_3158_),
    .B(_0900_),
    .C(_3181_),
    .D(_0990_),
    .X(_2284_));
 sky130_fd_sc_hd__or3_1 _5988_ (.A(_3111_),
    .B(_3095_),
    .C(_1008_),
    .X(_2285_));
 sky130_fd_sc_hd__or4_1 _5989_ (.A(_3066_),
    .B(_3118_),
    .C(_3117_),
    .D(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__and3_1 _5990_ (.A(_3120_),
    .B(_0893_),
    .C(_1638_),
    .X(_2287_));
 sky130_fd_sc_hd__clkinv_2 _5991_ (.A(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a211o_1 _5992_ (.A1(_3102_),
    .A2(_3197_),
    .B1(_1611_),
    .C1(_0899_),
    .X(_2289_));
 sky130_fd_sc_hd__and4_1 _5993_ (.A(_2284_),
    .B(_2286_),
    .C(_2288_),
    .D(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__and4b_1 _5994_ (.A_N(_2244_),
    .B(_2283_),
    .C(_2290_),
    .D(_2135_),
    .X(_2291_));
 sky130_fd_sc_hd__and4_1 _5995_ (.A(_2123_),
    .B(_2279_),
    .C(_2282_),
    .D(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_2 _5996_ (.A(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__clkbuf_4 _5997_ (.A(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_0972_),
    .B(_0874_),
    .Y(_2295_));
 sky130_fd_sc_hd__buf_2 _5999_ (.A(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__buf_2 _6000_ (.A(_1003_),
    .X(_2297_));
 sky130_fd_sc_hd__o22a_1 _6001_ (.A1(\as2650.stack[3][0] ),
    .A2(_3341_),
    .B1(_3344_),
    .B2(\as2650.stack[2][0] ),
    .X(_2298_));
 sky130_fd_sc_hd__o221a_1 _6002_ (.A1(\as2650.stack[0][0] ),
    .A2(_3350_),
    .B1(_3353_),
    .B2(\as2650.stack[1][0] ),
    .C1(_0425_),
    .X(_2299_));
 sky130_fd_sc_hd__mux4_2 _6003_ (.A0(\as2650.stack[7][0] ),
    .A1(\as2650.stack[4][0] ),
    .A2(\as2650.stack[5][0] ),
    .A3(\as2650.stack[6][0] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_2300_));
 sky130_fd_sc_hd__a22oi_4 _6004_ (.A1(_2298_),
    .A2(_2299_),
    .B1(_2300_),
    .B2(_3337_),
    .Y(_2301_));
 sky130_fd_sc_hd__o221a_1 _6005_ (.A1(_3028_),
    .A2(_0647_),
    .B1(_1608_),
    .B2(_3030_),
    .C1(_0973_),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(_0635_),
    .A1(_1685_),
    .S(_1090_),
    .X(_2303_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_0635_),
    .B(_3081_),
    .Y(_2304_));
 sky130_fd_sc_hd__o211a_1 _6008_ (.A1(_3081_),
    .A2(_2303_),
    .B1(_2304_),
    .C1(_0892_),
    .X(_2305_));
 sky130_fd_sc_hd__nor2_1 _6009_ (.A(_2302_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__or2_1 _6010_ (.A(_0635_),
    .B(\as2650.ins_reg[2] ),
    .X(_2307_));
 sky130_fd_sc_hd__and2_1 _6011_ (.A(_2304_),
    .B(_2307_),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(_0635_),
    .A1(_2308_),
    .S(_1665_),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_1 _6013_ (.A(_1520_),
    .B(_1639_),
    .Y(_2310_));
 sky130_fd_sc_hd__a221o_1 _6014_ (.A1(_0983_),
    .A2(_3067_),
    .B1(_1639_),
    .B2(_2308_),
    .C1(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__o211a_1 _6015_ (.A1(_3226_),
    .A2(_2309_),
    .B1(_2311_),
    .C1(_0690_),
    .X(_2312_));
 sky130_fd_sc_hd__a211o_1 _6016_ (.A1(_3080_),
    .A2(_2306_),
    .B1(_2312_),
    .C1(_2120_),
    .X(_2313_));
 sky130_fd_sc_hd__a21oi_1 _6017_ (.A1(_1601_),
    .A2(_3239_),
    .B1(_3028_),
    .Y(_2314_));
 sky130_fd_sc_hd__and3_1 _6018_ (.A(_3028_),
    .B(_1601_),
    .C(_3239_),
    .X(_2315_));
 sky130_fd_sc_hd__o21a_1 _6019_ (.A1(_2314_),
    .A2(_2315_),
    .B1(_3119_),
    .X(_2316_));
 sky130_fd_sc_hd__a211o_1 _6020_ (.A1(_0635_),
    .A2(_1609_),
    .B1(_2316_),
    .C1(_2158_),
    .X(_2317_));
 sky130_fd_sc_hd__inv_2 _6021_ (.A(_2303_),
    .Y(_2318_));
 sky130_fd_sc_hd__clkbuf_4 _6022_ (.A(_0643_),
    .X(_2319_));
 sky130_fd_sc_hd__o221a_1 _6023_ (.A1(_0635_),
    .A2(_3228_),
    .B1(_1690_),
    .B2(_2318_),
    .C1(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__a31o_1 _6024_ (.A1(_2218_),
    .A2(_2313_),
    .A3(_2317_),
    .B1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__o221a_1 _6025_ (.A1(_0636_),
    .A2(_2296_),
    .B1(_2297_),
    .B2(_2301_),
    .C1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__buf_2 _6026_ (.A(_2008_),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _6027_ (.A0(_0636_),
    .A1(_2322_),
    .S(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__o21ai_1 _6028_ (.A1(_0636_),
    .A2(_2293_),
    .B1(_1786_),
    .Y(_2325_));
 sky130_fd_sc_hd__a21oi_1 _6029_ (.A1(_2294_),
    .A2(_2324_),
    .B1(_2325_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor2_1 _6030_ (.A(_3046_),
    .B(_2120_),
    .Y(_2326_));
 sky130_fd_sc_hd__or2_1 _6031_ (.A(_0660_),
    .B(_0635_),
    .X(_2327_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(_0660_),
    .B(_2307_),
    .Y(_2328_));
 sky130_fd_sc_hd__o21ai_1 _6033_ (.A1(_3081_),
    .A2(_2327_),
    .B1(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__o21a_1 _6034_ (.A1(_3046_),
    .A2(_2208_),
    .B1(_2158_),
    .X(_2330_));
 sky130_fd_sc_hd__inv_2 _6035_ (.A(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _6036_ (.A(\as2650.pc[1] ),
    .B(\as2650.pc[0] ),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(_2332_),
    .B(_2327_),
    .Y(_2333_));
 sky130_fd_sc_hd__a32o_1 _6038_ (.A1(_2208_),
    .A2(_2326_),
    .A3(_2329_),
    .B1(_2331_),
    .B2(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__xnor2_1 _6039_ (.A(net2),
    .B(_3276_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _6040_ (.A(net1),
    .B(_3239_),
    .Y(_2336_));
 sky130_fd_sc_hd__nor2_1 _6041_ (.A(_2335_),
    .B(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__a21o_1 _6042_ (.A1(_2335_),
    .A2(_2336_),
    .B1(_1772_),
    .X(_2338_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_3129_),
    .B(_3097_),
    .Y(_2339_));
 sky130_fd_sc_hd__o211ai_1 _6044_ (.A1(_2337_),
    .A2(_2338_),
    .B1(_2143_),
    .C1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__mux2_1 _6045_ (.A0(_0660_),
    .A1(_1735_),
    .S(_1091_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(_3129_),
    .A1(\as2650.addr_buff[1] ),
    .S(_1857_),
    .X(_2342_));
 sky130_fd_sc_hd__a2bb2o_1 _6047_ (.A1_N(_1732_),
    .A2_N(_2333_),
    .B1(_2342_),
    .B2(_0973_),
    .X(_2343_));
 sky130_fd_sc_hd__a211o_1 _6048_ (.A1(_1699_),
    .A2(_2341_),
    .B1(_2343_),
    .C1(_2120_),
    .X(_2344_));
 sky130_fd_sc_hd__a21oi_1 _6049_ (.A1(_2340_),
    .A2(_2344_),
    .B1(_0889_),
    .Y(_2345_));
 sky130_fd_sc_hd__a211o_1 _6050_ (.A1(_1609_),
    .A2(_2334_),
    .B1(_2345_),
    .C1(_2319_),
    .X(_2346_));
 sky130_fd_sc_hd__o22a_1 _6051_ (.A1(\as2650.stack[7][1] ),
    .A2(_3342_),
    .B1(_3346_),
    .B2(\as2650.stack[6][1] ),
    .X(_2347_));
 sky130_fd_sc_hd__o22a_1 _6052_ (.A1(\as2650.stack[4][1] ),
    .A2(_3351_),
    .B1(_3355_),
    .B2(\as2650.stack[5][1] ),
    .X(_2348_));
 sky130_fd_sc_hd__and3_1 _6053_ (.A(\as2650.psu[2] ),
    .B(\as2650.stack[3][1] ),
    .C(_3335_),
    .X(_2349_));
 sky130_fd_sc_hd__o22a_1 _6054_ (.A1(\as2650.stack[0][1] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[1][1] ),
    .X(_2350_));
 sky130_fd_sc_hd__o221a_1 _6055_ (.A1(\as2650.stack[2][1] ),
    .A2(_3345_),
    .B1(_2349_),
    .B2(_3334_),
    .C1(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__a31o_2 _6056_ (.A1(_3338_),
    .A2(_2347_),
    .A3(_2348_),
    .B1(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__inv_2 _6057_ (.A(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__nor2_1 _6058_ (.A(_0888_),
    .B(_2341_),
    .Y(_2354_));
 sky130_fd_sc_hd__a211o_1 _6059_ (.A1(_0889_),
    .A2(_2333_),
    .B1(_2354_),
    .C1(_2218_),
    .X(_2355_));
 sky130_fd_sc_hd__o221a_1 _6060_ (.A1(_2296_),
    .A2(_2333_),
    .B1(_2353_),
    .B2(_2297_),
    .C1(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__a21oi_1 _6061_ (.A1(_2346_),
    .A2(_2356_),
    .B1(_1882_),
    .Y(_2357_));
 sky130_fd_sc_hd__buf_2 _6062_ (.A(_2293_),
    .X(_2358_));
 sky130_fd_sc_hd__o21ai_1 _6063_ (.A1(_2323_),
    .A2(_2333_),
    .B1(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__o221a_1 _6064_ (.A1(_0661_),
    .A2(_2294_),
    .B1(_2357_),
    .B2(_2359_),
    .C1(_1709_),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _6065_ (.A(_1484_),
    .B(_2332_),
    .Y(_2360_));
 sky130_fd_sc_hd__and2_1 _6066_ (.A(_1484_),
    .B(_2332_),
    .X(_2361_));
 sky130_fd_sc_hd__nor2_1 _6067_ (.A(_2360_),
    .B(_2361_),
    .Y(_2362_));
 sky130_fd_sc_hd__and3_1 _6068_ (.A(\as2650.pc[2] ),
    .B(_0660_),
    .C(_2307_),
    .X(_2363_));
 sky130_fd_sc_hd__a21oi_1 _6069_ (.A1(_0660_),
    .A2(_2307_),
    .B1(\as2650.pc[2] ),
    .Y(_2364_));
 sky130_fd_sc_hd__nand2_2 _6070_ (.A(_3121_),
    .B(_2208_),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_2 _6071_ (.A(_0641_),
    .B(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__o21ai_1 _6072_ (.A1(_2363_),
    .A2(_2364_),
    .B1(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__and2_1 _6073_ (.A(_3128_),
    .B(_3276_),
    .X(_2368_));
 sky130_fd_sc_hd__nand2_1 _6074_ (.A(net3),
    .B(_3392_),
    .Y(_2369_));
 sky130_fd_sc_hd__or2_1 _6075_ (.A(net3),
    .B(_3392_),
    .X(_2370_));
 sky130_fd_sc_hd__o211ai_2 _6076_ (.A1(_2368_),
    .A2(_2337_),
    .B1(_2369_),
    .C1(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__a211o_1 _6077_ (.A1(_2369_),
    .A2(_2370_),
    .B1(_2368_),
    .C1(_2337_),
    .X(_2372_));
 sky130_fd_sc_hd__a21oi_1 _6078_ (.A1(_2371_),
    .A2(_2372_),
    .B1(_0647_),
    .Y(_2373_));
 sky130_fd_sc_hd__a21oi_1 _6079_ (.A1(_1051_),
    .A2(_1857_),
    .B1(_2373_),
    .Y(_2374_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(_1484_),
    .A1(_1778_),
    .S(_1091_),
    .X(_2375_));
 sky130_fd_sc_hd__nor2_1 _6081_ (.A(_3085_),
    .B(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(_3131_),
    .A1(\as2650.addr_buff[2] ),
    .S(_1857_),
    .X(_2377_));
 sky130_fd_sc_hd__a221o_1 _6083_ (.A1(_0973_),
    .A2(_2377_),
    .B1(_2362_),
    .B2(_1692_),
    .C1(_0641_),
    .X(_2378_));
 sky130_fd_sc_hd__o22a_1 _6084_ (.A1(_3113_),
    .A2(_2374_),
    .B1(_2376_),
    .B2(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__o21a_1 _6085_ (.A1(_0888_),
    .A2(_2379_),
    .B1(_2218_),
    .X(_2380_));
 sky130_fd_sc_hd__or2_1 _6086_ (.A(_0891_),
    .B(_2330_),
    .X(_2381_));
 sky130_fd_sc_hd__or2_1 _6087_ (.A(_2362_),
    .B(_2381_),
    .X(_2382_));
 sky130_fd_sc_hd__o21ai_1 _6088_ (.A1(_3228_),
    .A2(_2362_),
    .B1(_2319_),
    .Y(_2383_));
 sky130_fd_sc_hd__a21oi_1 _6089_ (.A1(_1740_),
    .A2(_2375_),
    .B1(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__a31o_1 _6090_ (.A1(_2367_),
    .A2(_2380_),
    .A3(_2382_),
    .B1(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__o22a_1 _6091_ (.A1(\as2650.stack[5][2] ),
    .A2(_3355_),
    .B1(_3346_),
    .B2(\as2650.stack[6][2] ),
    .X(_2386_));
 sky130_fd_sc_hd__o22a_1 _6092_ (.A1(\as2650.stack[7][2] ),
    .A2(_3342_),
    .B1(_3351_),
    .B2(\as2650.stack[4][2] ),
    .X(_2387_));
 sky130_fd_sc_hd__and3_1 _6093_ (.A(\as2650.psu[2] ),
    .B(\as2650.stack[3][2] ),
    .C(_3335_),
    .X(_2388_));
 sky130_fd_sc_hd__o22a_1 _6094_ (.A1(\as2650.stack[0][2] ),
    .A2(_3351_),
    .B1(_3354_),
    .B2(\as2650.stack[1][2] ),
    .X(_2389_));
 sky130_fd_sc_hd__o221a_1 _6095_ (.A1(\as2650.stack[2][2] ),
    .A2(_3346_),
    .B1(_2388_),
    .B2(_3334_),
    .C1(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__a31o_1 _6096_ (.A1(_3338_),
    .A2(_2386_),
    .A3(_2387_),
    .B1(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__o221a_1 _6097_ (.A1(_2296_),
    .A2(_2362_),
    .B1(_2391_),
    .B2(_2297_),
    .C1(_2008_),
    .X(_2392_));
 sky130_fd_sc_hd__clkinv_2 _6098_ (.A(_2293_),
    .Y(_2393_));
 sky130_fd_sc_hd__a221o_1 _6099_ (.A1(_1882_),
    .A2(_2362_),
    .B1(_2385_),
    .B2(_2392_),
    .C1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__o211a_1 _6100_ (.A1(\as2650.pc[2] ),
    .A2(_2294_),
    .B1(_2394_),
    .C1(_1745_),
    .X(_0218_));
 sky130_fd_sc_hd__and2_1 _6101_ (.A(\as2650.pc[3] ),
    .B(_2360_),
    .X(_2395_));
 sky130_fd_sc_hd__nor2_1 _6102_ (.A(_0668_),
    .B(_2360_),
    .Y(_2396_));
 sky130_fd_sc_hd__or2_2 _6103_ (.A(_2395_),
    .B(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__nor2_1 _6104_ (.A(_2323_),
    .B(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hd__o22a_1 _6105_ (.A1(\as2650.stack[7][3] ),
    .A2(_3341_),
    .B1(_3345_),
    .B2(\as2650.stack[6][3] ),
    .X(_2399_));
 sky130_fd_sc_hd__o221a_1 _6106_ (.A1(\as2650.stack[4][3] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[5][3] ),
    .C1(_3337_),
    .X(_2400_));
 sky130_fd_sc_hd__o22a_1 _6107_ (.A1(\as2650.stack[3][3] ),
    .A2(_3341_),
    .B1(_3345_),
    .B2(\as2650.stack[2][3] ),
    .X(_2401_));
 sky130_fd_sc_hd__o221a_1 _6108_ (.A1(\as2650.stack[0][3] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[1][3] ),
    .C1(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__a22o_1 _6109_ (.A1(_2399_),
    .A2(_2400_),
    .B1(_2402_),
    .B2(_0425_),
    .X(_2403_));
 sky130_fd_sc_hd__inv_2 _6110_ (.A(_2403_),
    .Y(_2404_));
 sky130_fd_sc_hd__and2_1 _6111_ (.A(net4),
    .B(_0349_),
    .X(_2405_));
 sky130_fd_sc_hd__nor2_1 _6112_ (.A(_3134_),
    .B(_0349_),
    .Y(_2406_));
 sky130_fd_sc_hd__o211a_1 _6113_ (.A1(_2405_),
    .A2(_2406_),
    .B1(_2369_),
    .C1(_2371_),
    .X(_2407_));
 sky130_fd_sc_hd__a211oi_2 _6114_ (.A1(_2369_),
    .A2(_2371_),
    .B1(_2405_),
    .C1(_2406_),
    .Y(_2408_));
 sky130_fd_sc_hd__nand2_1 _6115_ (.A(_3135_),
    .B(_0647_),
    .Y(_2409_));
 sky130_fd_sc_hd__nor2_1 _6116_ (.A(_2158_),
    .B(_1609_),
    .Y(_2410_));
 sky130_fd_sc_hd__o311a_1 _6117_ (.A1(_0647_),
    .A2(_2407_),
    .A3(_2408_),
    .B1(_2409_),
    .C1(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__a31o_1 _6118_ (.A1(_2120_),
    .A2(_1609_),
    .A3(_2397_),
    .B1(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _6119_ (.A0(_0668_),
    .A1(_1792_),
    .S(_1090_),
    .X(_2413_));
 sky130_fd_sc_hd__inv_2 _6120_ (.A(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__o221a_1 _6121_ (.A1(_1690_),
    .A2(_2414_),
    .B1(_2397_),
    .B2(_3228_),
    .C1(_2319_),
    .X(_2415_));
 sky130_fd_sc_hd__and2_1 _6122_ (.A(_0668_),
    .B(_2363_),
    .X(_2416_));
 sky130_fd_sc_hd__nor2_1 _6123_ (.A(_0668_),
    .B(_2363_),
    .Y(_2417_));
 sky130_fd_sc_hd__or3_1 _6124_ (.A(_2365_),
    .B(_2416_),
    .C(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__nand2_1 _6125_ (.A(\as2650.addr_buff[3] ),
    .B(_3097_),
    .Y(_2419_));
 sky130_fd_sc_hd__o211a_1 _6126_ (.A1(_0818_),
    .A2(_3097_),
    .B1(_2419_),
    .C1(_0902_),
    .X(_2420_));
 sky130_fd_sc_hd__a211o_1 _6127_ (.A1(_1692_),
    .A2(_2397_),
    .B1(_2420_),
    .C1(_3121_),
    .X(_2421_));
 sky130_fd_sc_hd__a21o_1 _6128_ (.A1(_1699_),
    .A2(_2414_),
    .B1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__o211a_1 _6129_ (.A1(_2209_),
    .A2(_2397_),
    .B1(_2422_),
    .C1(_1640_),
    .X(_2423_));
 sky130_fd_sc_hd__nand2_1 _6130_ (.A(_2418_),
    .B(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__or3b_1 _6131_ (.A(_2412_),
    .B(_2415_),
    .C_N(_2424_),
    .X(_2425_));
 sky130_fd_sc_hd__o221a_1 _6132_ (.A1(_2296_),
    .A2(_2397_),
    .B1(_2404_),
    .B2(_2297_),
    .C1(_2425_),
    .X(_2426_));
 sky130_fd_sc_hd__o21ai_1 _6133_ (.A1(_1882_),
    .A2(_2426_),
    .B1(_2358_),
    .Y(_2427_));
 sky130_fd_sc_hd__o221a_1 _6134_ (.A1(_0668_),
    .A2(_2358_),
    .B1(_2398_),
    .B2(_2427_),
    .C1(_1709_),
    .X(_0219_));
 sky130_fd_sc_hd__xnor2_2 _6135_ (.A(\as2650.pc[4] ),
    .B(_2395_),
    .Y(_2428_));
 sky130_fd_sc_hd__mux4_2 _6136_ (.A0(\as2650.stack[7][4] ),
    .A1(\as2650.stack[4][4] ),
    .A2(\as2650.stack[5][4] ),
    .A3(\as2650.stack[6][4] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_2429_));
 sky130_fd_sc_hd__o22a_1 _6137_ (.A1(\as2650.stack[3][4] ),
    .A2(_3341_),
    .B1(_3345_),
    .B2(\as2650.stack[2][4] ),
    .X(_2430_));
 sky130_fd_sc_hd__o221a_1 _6138_ (.A1(\as2650.stack[0][4] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[1][4] ),
    .C1(_0425_),
    .X(_2431_));
 sky130_fd_sc_hd__a22oi_4 _6139_ (.A1(_3337_),
    .A2(_2429_),
    .B1(_2430_),
    .B2(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__nor2_2 _6140_ (.A(_3119_),
    .B(_2330_),
    .Y(_2433_));
 sky130_fd_sc_hd__xnor2_1 _6141_ (.A(_0672_),
    .B(_2416_),
    .Y(_2434_));
 sky130_fd_sc_hd__nor2_1 _6142_ (.A(_1696_),
    .B(_3121_),
    .Y(_2435_));
 sky130_fd_sc_hd__nand2_1 _6143_ (.A(_3137_),
    .B(_3097_),
    .Y(_2436_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(net5),
    .B(_0409_),
    .Y(_2437_));
 sky130_fd_sc_hd__or2_1 _6145_ (.A(net5),
    .B(_0409_),
    .X(_2438_));
 sky130_fd_sc_hd__o211a_1 _6146_ (.A1(_2405_),
    .A2(_2408_),
    .B1(_2437_),
    .C1(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__a211o_1 _6147_ (.A1(_2437_),
    .A2(_2438_),
    .B1(_2405_),
    .C1(_2408_),
    .X(_2440_));
 sky130_fd_sc_hd__or3b_1 _6148_ (.A(_2439_),
    .B(_0647_),
    .C_N(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(_1490_),
    .A1(_1854_),
    .S(_1090_),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_1 _6150_ (.A0(_3137_),
    .A1(\as2650.addr_buff[4] ),
    .S(_3326_),
    .X(_2443_));
 sky130_fd_sc_hd__inv_2 _6151_ (.A(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__o221a_1 _6152_ (.A1(_1731_),
    .A2(_2428_),
    .B1(_2444_),
    .B2(_3051_),
    .C1(_0646_),
    .X(_2445_));
 sky130_fd_sc_hd__o21a_1 _6153_ (.A1(_3085_),
    .A2(_2442_),
    .B1(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__a31o_1 _6154_ (.A1(_2143_),
    .A2(_2436_),
    .A3(_2441_),
    .B1(_2446_),
    .X(_2447_));
 sky130_fd_sc_hd__o221a_1 _6155_ (.A1(_3228_),
    .A2(_2428_),
    .B1(_2442_),
    .B2(_1690_),
    .C1(_0643_),
    .X(_2448_));
 sky130_fd_sc_hd__a21o_1 _6156_ (.A1(_2435_),
    .A2(_2447_),
    .B1(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__a31o_1 _6157_ (.A1(_2218_),
    .A2(_2366_),
    .A3(_2434_),
    .B1(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__a22o_1 _6158_ (.A1(_2433_),
    .A2(_2428_),
    .B1(_2450_),
    .B2(_2008_),
    .X(_2451_));
 sky130_fd_sc_hd__o21a_1 _6159_ (.A1(_2297_),
    .A2(_2432_),
    .B1(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__a21oi_1 _6160_ (.A1(_1882_),
    .A2(_2428_),
    .B1(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__o21ai_1 _6161_ (.A1(_2296_),
    .A2(_2428_),
    .B1(_2358_),
    .Y(_2454_));
 sky130_fd_sc_hd__o221a_1 _6162_ (.A1(_0672_),
    .A2(_2358_),
    .B1(_2453_),
    .B2(_2454_),
    .C1(_1709_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _6163_ (.A(\as2650.pc[5] ),
    .B(\as2650.pc[4] ),
    .C(_2395_),
    .X(_2455_));
 sky130_fd_sc_hd__a21oi_1 _6164_ (.A1(_0672_),
    .A2(_2395_),
    .B1(\as2650.pc[5] ),
    .Y(_2456_));
 sky130_fd_sc_hd__nor2_2 _6165_ (.A(_2455_),
    .B(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__and2_1 _6166_ (.A(net5),
    .B(_0409_),
    .X(_2458_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_3139_),
    .B(_0455_),
    .Y(_2459_));
 sky130_fd_sc_hd__or2_1 _6168_ (.A(_3139_),
    .B(_0455_),
    .X(_2460_));
 sky130_fd_sc_hd__o211a_1 _6169_ (.A1(_2458_),
    .A2(_2439_),
    .B1(_2459_),
    .C1(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__a211oi_1 _6170_ (.A1(_2459_),
    .A2(_2460_),
    .B1(_2458_),
    .C1(_2439_),
    .Y(_2462_));
 sky130_fd_sc_hd__o21ai_1 _6171_ (.A1(_2461_),
    .A2(_2462_),
    .B1(_1865_),
    .Y(_2463_));
 sky130_fd_sc_hd__o211a_1 _6172_ (.A1(_3140_),
    .A2(_1865_),
    .B1(_2410_),
    .C1(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__and3_1 _6173_ (.A(\as2650.pc[5] ),
    .B(\as2650.pc[4] ),
    .C(_2416_),
    .X(_2465_));
 sky130_fd_sc_hd__a21oi_1 _6174_ (.A1(_0672_),
    .A2(_2416_),
    .B1(\as2650.pc[5] ),
    .Y(_2466_));
 sky130_fd_sc_hd__mux2_1 _6175_ (.A0(\as2650.pc[5] ),
    .A1(_1878_),
    .S(_1090_),
    .X(_2467_));
 sky130_fd_sc_hd__a221o_1 _6176_ (.A1(_3140_),
    .A2(_1601_),
    .B1(_1857_),
    .B2(\as2650.addr_buff[5] ),
    .C1(_3051_),
    .X(_2468_));
 sky130_fd_sc_hd__o211a_1 _6177_ (.A1(_1731_),
    .A2(_2457_),
    .B1(_2468_),
    .C1(_3159_),
    .X(_2469_));
 sky130_fd_sc_hd__o21ai_1 _6178_ (.A1(_3085_),
    .A2(_2467_),
    .B1(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__o31a_1 _6179_ (.A1(_2365_),
    .A2(_2465_),
    .A3(_2466_),
    .B1(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__a2bb2o_1 _6180_ (.A1_N(_2120_),
    .A2_N(_2471_),
    .B1(_2457_),
    .B2(_2433_),
    .X(_2472_));
 sky130_fd_sc_hd__or3_1 _6181_ (.A(_1696_),
    .B(_2464_),
    .C(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__a221o_1 _6182_ (.A1(_1641_),
    .A2(_2457_),
    .B1(_2467_),
    .B2(_1740_),
    .C1(_1871_),
    .X(_2474_));
 sky130_fd_sc_hd__mux4_1 _6183_ (.A0(\as2650.stack[7][5] ),
    .A1(\as2650.stack[4][5] ),
    .A2(\as2650.stack[5][5] ),
    .A3(\as2650.stack[6][5] ),
    .S0(_3339_),
    .S1(_3343_),
    .X(_2475_));
 sky130_fd_sc_hd__and3_1 _6184_ (.A(\as2650.psu[2] ),
    .B(\as2650.stack[3][5] ),
    .C(_3335_),
    .X(_2476_));
 sky130_fd_sc_hd__o22a_1 _6185_ (.A1(\as2650.stack[0][5] ),
    .A2(_3350_),
    .B1(_3353_),
    .B2(\as2650.stack[1][5] ),
    .X(_2477_));
 sky130_fd_sc_hd__o221a_1 _6186_ (.A1(\as2650.stack[2][5] ),
    .A2(_3344_),
    .B1(_2476_),
    .B2(_3334_),
    .C1(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__a21o_1 _6187_ (.A1(_3337_),
    .A2(_2475_),
    .B1(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__a22o_1 _6188_ (.A1(_0991_),
    .A2(_2457_),
    .B1(_2479_),
    .B2(_2226_),
    .X(_2480_));
 sky130_fd_sc_hd__a21oi_1 _6189_ (.A1(_2473_),
    .A2(_2474_),
    .B1(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__nor2_1 _6190_ (.A(_1881_),
    .B(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__a211o_1 _6191_ (.A1(_1882_),
    .A2(_2457_),
    .B1(_2482_),
    .C1(_2393_),
    .X(_2483_));
 sky130_fd_sc_hd__o211a_1 _6192_ (.A1(_0676_),
    .A2(_2294_),
    .B1(_2483_),
    .C1(_1745_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_2 _6193_ (.A(_0680_),
    .B(_2455_),
    .X(_2484_));
 sky130_fd_sc_hd__nor2_1 _6194_ (.A(_0680_),
    .B(_2455_),
    .Y(_2485_));
 sky130_fd_sc_hd__nor2_2 _6195_ (.A(_2484_),
    .B(_2485_),
    .Y(_2486_));
 sky130_fd_sc_hd__mux2_1 _6196_ (.A0(_0680_),
    .A1(_1935_),
    .S(_1091_),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(\as2650.addr_buff[6] ),
    .A1(_3144_),
    .S(_1608_),
    .X(_2488_));
 sky130_fd_sc_hd__a221o_1 _6198_ (.A1(_1692_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(_0973_),
    .C1(_2120_),
    .X(_2489_));
 sky130_fd_sc_hd__a21oi_1 _6199_ (.A1(_1699_),
    .A2(_2487_),
    .B1(_2489_),
    .Y(_2490_));
 sky130_fd_sc_hd__and2_1 _6200_ (.A(_3142_),
    .B(_0500_),
    .X(_2491_));
 sky130_fd_sc_hd__inv_2 _6201_ (.A(_2491_),
    .Y(_2492_));
 sky130_fd_sc_hd__or2_1 _6202_ (.A(_3142_),
    .B(_0500_),
    .X(_2493_));
 sky130_fd_sc_hd__inv_2 _6203_ (.A(_2459_),
    .Y(_2494_));
 sky130_fd_sc_hd__a211oi_1 _6204_ (.A1(_2492_),
    .A2(_2493_),
    .B1(_2494_),
    .C1(_2461_),
    .Y(_2495_));
 sky130_fd_sc_hd__o211a_1 _6205_ (.A1(_2494_),
    .A2(_2461_),
    .B1(_2492_),
    .C1(_2493_),
    .X(_2496_));
 sky130_fd_sc_hd__nand2_1 _6206_ (.A(_3144_),
    .B(_1772_),
    .Y(_2497_));
 sky130_fd_sc_hd__o311a_1 _6207_ (.A1(_1857_),
    .A2(_2495_),
    .A3(_2496_),
    .B1(_2497_),
    .C1(_2143_),
    .X(_2498_));
 sky130_fd_sc_hd__o21ai_1 _6208_ (.A1(_2490_),
    .A2(_2498_),
    .B1(_3330_),
    .Y(_2499_));
 sky130_fd_sc_hd__nand2_1 _6209_ (.A(_0680_),
    .B(_2465_),
    .Y(_2500_));
 sky130_fd_sc_hd__or2_1 _6210_ (.A(_0680_),
    .B(_2465_),
    .X(_2501_));
 sky130_fd_sc_hd__a211o_1 _6211_ (.A1(_2500_),
    .A2(_2501_),
    .B1(_2120_),
    .C1(_2365_),
    .X(_2502_));
 sky130_fd_sc_hd__o211a_1 _6212_ (.A1(_2381_),
    .A2(_2486_),
    .B1(_2502_),
    .C1(_2218_),
    .X(_2503_));
 sky130_fd_sc_hd__o221a_1 _6213_ (.A1(_1690_),
    .A2(_2487_),
    .B1(_2486_),
    .B2(_3228_),
    .C1(_2319_),
    .X(_2504_));
 sky130_fd_sc_hd__a21o_1 _6214_ (.A1(_2499_),
    .A2(_2503_),
    .B1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__o22a_1 _6215_ (.A1(\as2650.stack[7][6] ),
    .A2(_3341_),
    .B1(_3345_),
    .B2(\as2650.stack[6][6] ),
    .X(_2506_));
 sky130_fd_sc_hd__o22a_1 _6216_ (.A1(\as2650.stack[4][6] ),
    .A2(_3351_),
    .B1(_3354_),
    .B2(\as2650.stack[5][6] ),
    .X(_2507_));
 sky130_fd_sc_hd__and3_1 _6217_ (.A(\as2650.psu[2] ),
    .B(\as2650.stack[3][6] ),
    .C(_3335_),
    .X(_2508_));
 sky130_fd_sc_hd__o22a_1 _6218_ (.A1(\as2650.stack[0][6] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[1][6] ),
    .X(_2509_));
 sky130_fd_sc_hd__o221a_1 _6219_ (.A1(\as2650.stack[2][6] ),
    .A2(_3345_),
    .B1(_2508_),
    .B2(_3334_),
    .C1(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__a31o_2 _6220_ (.A1(_3337_),
    .A2(_2506_),
    .A3(_2507_),
    .B1(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__or2_1 _6221_ (.A(_2297_),
    .B(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__o211a_1 _6222_ (.A1(_2296_),
    .A2(_2486_),
    .B1(_2512_),
    .C1(_2008_),
    .X(_2513_));
 sky130_fd_sc_hd__a221o_1 _6223_ (.A1(_1882_),
    .A2(_2486_),
    .B1(_2505_),
    .B2(_2513_),
    .C1(_2393_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_4 _6224_ (.A(_3154_),
    .X(_2515_));
 sky130_fd_sc_hd__o211a_1 _6225_ (.A1(_0681_),
    .A2(_2294_),
    .B1(_2514_),
    .C1(_2515_),
    .X(_0222_));
 sky130_fd_sc_hd__xnor2_2 _6226_ (.A(\as2650.pc[7] ),
    .B(_2484_),
    .Y(_2516_));
 sky130_fd_sc_hd__mux2_1 _6227_ (.A0(\as2650.pc[7] ),
    .A1(_1950_),
    .S(_1090_),
    .X(_2517_));
 sky130_fd_sc_hd__nand2_1 _6228_ (.A(_1740_),
    .B(_2517_),
    .Y(_2518_));
 sky130_fd_sc_hd__or2_1 _6229_ (.A(_3228_),
    .B(_2516_),
    .X(_2519_));
 sky130_fd_sc_hd__and3_1 _6230_ (.A(\as2650.pc[7] ),
    .B(_0680_),
    .C(_2465_),
    .X(_2520_));
 sky130_fd_sc_hd__a21oi_1 _6231_ (.A1(_0680_),
    .A2(_2465_),
    .B1(\as2650.pc[7] ),
    .Y(_2521_));
 sky130_fd_sc_hd__mux2_1 _6232_ (.A0(_3151_),
    .A1(_3146_),
    .S(_1607_),
    .X(_2522_));
 sky130_fd_sc_hd__o2bb2a_1 _6233_ (.A1_N(_1692_),
    .A2_N(_2516_),
    .B1(_2522_),
    .B2(_3051_),
    .X(_2523_));
 sky130_fd_sc_hd__o211ai_1 _6234_ (.A1(_3085_),
    .A2(_2517_),
    .B1(_2523_),
    .C1(_3159_),
    .Y(_2524_));
 sky130_fd_sc_hd__o31a_1 _6235_ (.A1(_2365_),
    .A2(_2520_),
    .A3(_2521_),
    .B1(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__nand2_1 _6236_ (.A(net8),
    .B(_3265_),
    .Y(_2526_));
 sky130_fd_sc_hd__or2_1 _6237_ (.A(net8),
    .B(_3265_),
    .X(_2527_));
 sky130_fd_sc_hd__nand2_1 _6238_ (.A(_2526_),
    .B(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__nor2_1 _6239_ (.A(_2491_),
    .B(_2496_),
    .Y(_2529_));
 sky130_fd_sc_hd__xnor2_1 _6240_ (.A(_2528_),
    .B(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__a21bo_1 _6241_ (.A1(_1865_),
    .A2(_2530_),
    .B1_N(_2410_),
    .X(_2531_));
 sky130_fd_sc_hd__nor2_1 _6242_ (.A(_3148_),
    .B(_1865_),
    .Y(_2532_));
 sky130_fd_sc_hd__o221a_1 _6243_ (.A1(_0641_),
    .A2(_2525_),
    .B1(_2531_),
    .B2(_2532_),
    .C1(_3076_),
    .X(_2533_));
 sky130_fd_sc_hd__o21a_1 _6244_ (.A1(_2381_),
    .A2(_2516_),
    .B1(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__a31o_1 _6245_ (.A1(_2319_),
    .A2(_2518_),
    .A3(_2519_),
    .B1(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__o22a_1 _6246_ (.A1(\as2650.stack[7][7] ),
    .A2(_3341_),
    .B1(_3344_),
    .B2(\as2650.stack[6][7] ),
    .X(_2536_));
 sky130_fd_sc_hd__o221a_1 _6247_ (.A1(\as2650.stack[4][7] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[5][7] ),
    .C1(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__o22a_1 _6248_ (.A1(\as2650.stack[0][7] ),
    .A2(_3350_),
    .B1(_3354_),
    .B2(\as2650.stack[1][7] ),
    .X(_2538_));
 sky130_fd_sc_hd__o221a_1 _6249_ (.A1(\as2650.stack[3][7] ),
    .A2(_3341_),
    .B1(_3345_),
    .B2(\as2650.stack[2][7] ),
    .C1(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_2 _6250_ (.A0(_2537_),
    .A1(_2539_),
    .S(_0425_),
    .X(_2540_));
 sky130_fd_sc_hd__o2bb2a_1 _6251_ (.A1_N(_2226_),
    .A2_N(_2540_),
    .B1(_2516_),
    .B2(_2296_),
    .X(_2541_));
 sky130_fd_sc_hd__a21o_1 _6252_ (.A1(_2535_),
    .A2(_2541_),
    .B1(_1881_),
    .X(_2542_));
 sky130_fd_sc_hd__o211ai_1 _6253_ (.A1(_2323_),
    .A2(_2516_),
    .B1(_2542_),
    .C1(_2358_),
    .Y(_2543_));
 sky130_fd_sc_hd__o211a_1 _6254_ (.A1(_0685_),
    .A2(_2294_),
    .B1(_2543_),
    .C1(_2515_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _6255_ (.A(\as2650.pc[8] ),
    .B(\as2650.pc[7] ),
    .C(_2484_),
    .X(_2544_));
 sky130_fd_sc_hd__a21oi_1 _6256_ (.A1(\as2650.pc[7] ),
    .A2(_2484_),
    .B1(_0689_),
    .Y(_2545_));
 sky130_fd_sc_hd__nor2_2 _6257_ (.A(_2544_),
    .B(_2545_),
    .Y(_2546_));
 sky130_fd_sc_hd__o21a_1 _6258_ (.A1(_2528_),
    .A2(_2529_),
    .B1(_2526_),
    .X(_2547_));
 sky130_fd_sc_hd__nor2_1 _6259_ (.A(_0647_),
    .B(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__a21oi_1 _6260_ (.A1(_3030_),
    .A2(_2548_),
    .B1(_3113_),
    .Y(_2549_));
 sky130_fd_sc_hd__o21ai_1 _6261_ (.A1(_3030_),
    .A2(_2548_),
    .B1(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__mux2_1 _6262_ (.A0(_2005_),
    .A1(_2001_),
    .S(_1091_),
    .X(_2551_));
 sky130_fd_sc_hd__mux2_1 _6263_ (.A0(_3028_),
    .A1(_3030_),
    .S(_1608_),
    .X(_2552_));
 sky130_fd_sc_hd__o221a_1 _6264_ (.A1(_1732_),
    .A2(_2546_),
    .B1(_2552_),
    .B2(_0892_),
    .C1(_2158_),
    .X(_2553_));
 sky130_fd_sc_hd__a21bo_1 _6265_ (.A1(_1699_),
    .A2(_2551_),
    .B1_N(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__a21oi_1 _6266_ (.A1(_2550_),
    .A2(_2554_),
    .B1(_0889_),
    .Y(_2555_));
 sky130_fd_sc_hd__nand2_1 _6267_ (.A(_0689_),
    .B(_2520_),
    .Y(_2556_));
 sky130_fd_sc_hd__or2_1 _6268_ (.A(_0689_),
    .B(_2520_),
    .X(_2557_));
 sky130_fd_sc_hd__a31o_1 _6269_ (.A1(_2366_),
    .A2(_2556_),
    .A3(_2557_),
    .B1(_2319_),
    .X(_2558_));
 sky130_fd_sc_hd__a211o_1 _6270_ (.A1(_2433_),
    .A2(_2546_),
    .B1(_2555_),
    .C1(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__nor2_1 _6271_ (.A(_0888_),
    .B(_2551_),
    .Y(_2560_));
 sky130_fd_sc_hd__a211o_1 _6272_ (.A1(_0888_),
    .A2(_2546_),
    .B1(_2560_),
    .C1(_2218_),
    .X(_2561_));
 sky130_fd_sc_hd__o22a_1 _6273_ (.A1(_3360_),
    .A2(_2297_),
    .B1(_2546_),
    .B2(_2296_),
    .X(_2562_));
 sky130_fd_sc_hd__and3_1 _6274_ (.A(_2008_),
    .B(_2561_),
    .C(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a221o_1 _6275_ (.A1(_1882_),
    .A2(_2546_),
    .B1(_2559_),
    .B2(_2563_),
    .C1(_2393_),
    .X(_2564_));
 sky130_fd_sc_hd__o211a_1 _6276_ (.A1(_0689_),
    .A2(_2294_),
    .B1(_2564_),
    .C1(_2515_),
    .X(_0224_));
 sky130_fd_sc_hd__and2_1 _6277_ (.A(\as2650.pc[9] ),
    .B(_2544_),
    .X(_2565_));
 sky130_fd_sc_hd__nor2_1 _6278_ (.A(_0704_),
    .B(_2544_),
    .Y(_2566_));
 sky130_fd_sc_hd__or2_2 _6279_ (.A(_2565_),
    .B(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__nor2_1 _6280_ (.A(_2323_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__and3_1 _6281_ (.A(_0704_),
    .B(_0689_),
    .C(_2520_),
    .X(_2569_));
 sky130_fd_sc_hd__a21oi_1 _6282_ (.A1(_0689_),
    .A2(_2520_),
    .B1(_0704_),
    .Y(_2570_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(_0704_),
    .A1(_2035_),
    .S(_1090_),
    .X(_2571_));
 sky130_fd_sc_hd__nor2_1 _6284_ (.A(_3084_),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__nand2_1 _6285_ (.A(\as2650.addr_buff[1] ),
    .B(_1601_),
    .Y(_2573_));
 sky130_fd_sc_hd__a32o_1 _6286_ (.A1(_0902_),
    .A2(_2573_),
    .A3(_2339_),
    .B1(_2567_),
    .B2(_1692_),
    .X(_2574_));
 sky130_fd_sc_hd__or3_1 _6287_ (.A(_0690_),
    .B(_2572_),
    .C(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__o31a_1 _6288_ (.A1(_2365_),
    .A2(_2569_),
    .A3(_2570_),
    .B1(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__or2_1 _6289_ (.A(_2120_),
    .B(_2576_),
    .X(_2577_));
 sky130_fd_sc_hd__a21oi_1 _6290_ (.A1(_3030_),
    .A2(_2548_),
    .B1(\as2650.addr_buff[1] ),
    .Y(_2578_));
 sky130_fd_sc_hd__and3b_1 _6291_ (.A_N(_2547_),
    .B(_2018_),
    .C(_1601_),
    .X(_2579_));
 sky130_fd_sc_hd__or3b_1 _6292_ (.A(_2578_),
    .B(_2579_),
    .C_N(_2410_),
    .X(_2580_));
 sky130_fd_sc_hd__o211a_1 _6293_ (.A1(_2381_),
    .A2(_2567_),
    .B1(_2577_),
    .C1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__nor2_1 _6294_ (.A(_0887_),
    .B(_2571_),
    .Y(_2582_));
 sky130_fd_sc_hd__a211o_1 _6295_ (.A1(_0907_),
    .A2(_2567_),
    .B1(_2582_),
    .C1(_2218_),
    .X(_2583_));
 sky130_fd_sc_hd__o221a_1 _6296_ (.A1(_0321_),
    .A2(_2297_),
    .B1(_2567_),
    .B2(_2296_),
    .C1(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__o21ai_1 _6297_ (.A1(_2319_),
    .A2(_2581_),
    .B1(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__a21o_1 _6298_ (.A1(_2323_),
    .A2(_2585_),
    .B1(_2393_),
    .X(_2586_));
 sky130_fd_sc_hd__o221a_1 _6299_ (.A1(_0704_),
    .A2(_2358_),
    .B1(_2568_),
    .B2(_2586_),
    .C1(_1709_),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_2 _6300_ (.A(_0713_),
    .B(_2565_),
    .Y(_2587_));
 sky130_fd_sc_hd__nor2_1 _6301_ (.A(\as2650.addr_buff[2] ),
    .B(_2579_),
    .Y(_2588_));
 sky130_fd_sc_hd__a21o_1 _6302_ (.A1(_2051_),
    .A2(_2548_),
    .B1(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__clkinv_2 _6303_ (.A(\as2650.pc[10] ),
    .Y(_2590_));
 sky130_fd_sc_hd__mux2_1 _6304_ (.A0(_2590_),
    .A1(_2059_),
    .S(_1090_),
    .X(_2591_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(_3131_),
    .A1(\as2650.addr_buff[2] ),
    .S(_1607_),
    .X(_2592_));
 sky130_fd_sc_hd__a21oi_1 _6306_ (.A1(_0973_),
    .A2(_2592_),
    .B1(_0641_),
    .Y(_2593_));
 sky130_fd_sc_hd__o221a_1 _6307_ (.A1(_3085_),
    .A2(_2591_),
    .B1(_2587_),
    .B2(_1732_),
    .C1(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__a21o_1 _6308_ (.A1(_2143_),
    .A2(_2589_),
    .B1(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__xnor2_1 _6309_ (.A(_0713_),
    .B(_2569_),
    .Y(_2596_));
 sky130_fd_sc_hd__a22o_1 _6310_ (.A1(_0767_),
    .A2(_2595_),
    .B1(_2596_),
    .B2(_2366_),
    .X(_2597_));
 sky130_fd_sc_hd__a211o_1 _6311_ (.A1(_2433_),
    .A2(_2587_),
    .B1(_2597_),
    .C1(_1696_),
    .X(_2598_));
 sky130_fd_sc_hd__a221o_1 _6312_ (.A1(_1740_),
    .A2(_2591_),
    .B1(_2587_),
    .B2(_1641_),
    .C1(_1871_),
    .X(_2599_));
 sky130_fd_sc_hd__nand2_1 _6313_ (.A(_2598_),
    .B(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__o2bb2a_1 _6314_ (.A1_N(_0991_),
    .A2_N(_2587_),
    .B1(_2297_),
    .B2(_0332_),
    .X(_2601_));
 sky130_fd_sc_hd__o21ai_1 _6315_ (.A1(_2008_),
    .A2(_2587_),
    .B1(_2293_),
    .Y(_2602_));
 sky130_fd_sc_hd__a31o_1 _6316_ (.A1(_2323_),
    .A2(_2600_),
    .A3(_2601_),
    .B1(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o211a_1 _6317_ (.A1(_0713_),
    .A2(_2294_),
    .B1(_2603_),
    .C1(_2515_),
    .X(_0226_));
 sky130_fd_sc_hd__and3_1 _6318_ (.A(_0719_),
    .B(\as2650.pc[10] ),
    .C(_2565_),
    .X(_2604_));
 sky130_fd_sc_hd__a21oi_1 _6319_ (.A1(_0713_),
    .A2(_2565_),
    .B1(_0719_),
    .Y(_2605_));
 sky130_fd_sc_hd__or2_1 _6320_ (.A(_2604_),
    .B(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__mux2_1 _6321_ (.A0(_0719_),
    .A1(_2071_),
    .S(_1090_),
    .X(_2607_));
 sky130_fd_sc_hd__nor2_1 _6322_ (.A(_0889_),
    .B(_2607_),
    .Y(_2608_));
 sky130_fd_sc_hd__a211o_1 _6323_ (.A1(_0889_),
    .A2(_2606_),
    .B1(_2608_),
    .C1(_2218_),
    .X(_2609_));
 sky130_fd_sc_hd__a21oi_1 _6324_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2579_),
    .B1(\as2650.addr_buff[3] ),
    .Y(_2610_));
 sky130_fd_sc_hd__and2_1 _6325_ (.A(_2094_),
    .B(_2579_),
    .X(_2611_));
 sky130_fd_sc_hd__o21ai_1 _6326_ (.A1(_2610_),
    .A2(_2611_),
    .B1(_2143_),
    .Y(_2612_));
 sky130_fd_sc_hd__mux2_1 _6327_ (.A0(_3135_),
    .A1(\as2650.addr_buff[3] ),
    .S(_1607_),
    .X(_2613_));
 sky130_fd_sc_hd__a2bb2o_1 _6328_ (.A1_N(_1732_),
    .A2_N(_2606_),
    .B1(_2613_),
    .B2(_0973_),
    .X(_2614_));
 sky130_fd_sc_hd__a211o_1 _6329_ (.A1(_1699_),
    .A2(_2607_),
    .B1(_2614_),
    .C1(_0641_),
    .X(_2615_));
 sky130_fd_sc_hd__a21oi_1 _6330_ (.A1(_2612_),
    .A2(_2615_),
    .B1(_0888_),
    .Y(_2616_));
 sky130_fd_sc_hd__and3_1 _6331_ (.A(_0719_),
    .B(\as2650.pc[10] ),
    .C(_2569_),
    .X(_2617_));
 sky130_fd_sc_hd__a21oi_1 _6332_ (.A1(_0713_),
    .A2(_2569_),
    .B1(_0719_),
    .Y(_2618_));
 sky130_fd_sc_hd__o21a_1 _6333_ (.A1(_2617_),
    .A2(_2618_),
    .B1(_2366_),
    .X(_2619_));
 sky130_fd_sc_hd__a2111o_1 _6334_ (.A1(_2433_),
    .A2(_2606_),
    .B1(_2616_),
    .C1(_2619_),
    .D1(_2319_),
    .X(_2620_));
 sky130_fd_sc_hd__o221a_1 _6335_ (.A1(_0430_),
    .A2(_2297_),
    .B1(_2606_),
    .B2(_2296_),
    .C1(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__a21oi_1 _6336_ (.A1(_2609_),
    .A2(_2621_),
    .B1(_1882_),
    .Y(_2622_));
 sky130_fd_sc_hd__o21ai_1 _6337_ (.A1(_2323_),
    .A2(_2606_),
    .B1(_2358_),
    .Y(_2623_));
 sky130_fd_sc_hd__o221a_1 _6338_ (.A1(_0719_),
    .A2(_2358_),
    .B1(_2622_),
    .B2(_2623_),
    .C1(_1709_),
    .X(_0227_));
 sky130_fd_sc_hd__and2_1 _6339_ (.A(_0726_),
    .B(_2604_),
    .X(_2624_));
 sky130_fd_sc_hd__nor2_1 _6340_ (.A(_0726_),
    .B(_2604_),
    .Y(_2625_));
 sky130_fd_sc_hd__nor2_2 _6341_ (.A(_2624_),
    .B(_2625_),
    .Y(_2626_));
 sky130_fd_sc_hd__or2_1 _6342_ (.A(_2008_),
    .B(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__xnor2_1 _6343_ (.A(\as2650.addr_buff[4] ),
    .B(_2611_),
    .Y(_2628_));
 sky130_fd_sc_hd__mux2_1 _6344_ (.A0(_0726_),
    .A1(_2106_),
    .S(_1090_),
    .X(_2629_));
 sky130_fd_sc_hd__o21ai_1 _6345_ (.A1(_2091_),
    .A2(_1857_),
    .B1(_2436_),
    .Y(_2630_));
 sky130_fd_sc_hd__a221o_1 _6346_ (.A1(_1692_),
    .A2(_2626_),
    .B1(_2630_),
    .B2(_0902_),
    .C1(_0641_),
    .X(_2631_));
 sky130_fd_sc_hd__a21oi_1 _6347_ (.A1(_1699_),
    .A2(_2629_),
    .B1(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__a21oi_1 _6348_ (.A1(_2143_),
    .A2(_2628_),
    .B1(_2632_),
    .Y(_2633_));
 sky130_fd_sc_hd__and2_1 _6349_ (.A(_0726_),
    .B(_2617_),
    .X(_2634_));
 sky130_fd_sc_hd__nor2_1 _6350_ (.A(_0726_),
    .B(_2617_),
    .Y(_2635_));
 sky130_fd_sc_hd__o21ai_1 _6351_ (.A1(_2634_),
    .A2(_2635_),
    .B1(_2366_),
    .Y(_2636_));
 sky130_fd_sc_hd__o211a_1 _6352_ (.A1(_0691_),
    .A2(_2633_),
    .B1(_2636_),
    .C1(_1871_),
    .X(_2637_));
 sky130_fd_sc_hd__or2_1 _6353_ (.A(_3160_),
    .B(_2626_),
    .X(_2638_));
 sky130_fd_sc_hd__o211a_1 _6354_ (.A1(_0887_),
    .A2(_2629_),
    .B1(_2638_),
    .C1(_1696_),
    .X(_2639_));
 sky130_fd_sc_hd__o32a_1 _6355_ (.A1(_1881_),
    .A2(_2637_),
    .A3(_2639_),
    .B1(_2381_),
    .B2(_2626_),
    .X(_2640_));
 sky130_fd_sc_hd__a21o_1 _6356_ (.A1(_0488_),
    .A2(_2226_),
    .B1(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__a221o_1 _6357_ (.A1(_0991_),
    .A2(_2626_),
    .B1(_2627_),
    .B2(_2641_),
    .C1(_2393_),
    .X(_2642_));
 sky130_fd_sc_hd__o211a_1 _6358_ (.A1(_0726_),
    .A2(_2294_),
    .B1(_2642_),
    .C1(_2515_),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_1 _6359_ (.A(\as2650.pc[13] ),
    .B(_2624_),
    .Y(_2643_));
 sky130_fd_sc_hd__or2_1 _6360_ (.A(\as2650.pc[13] ),
    .B(_2624_),
    .X(_2644_));
 sky130_fd_sc_hd__nand2_1 _6361_ (.A(_2643_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__nor2_1 _6362_ (.A(_2323_),
    .B(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__or2_1 _6363_ (.A(\as2650.pc[13] ),
    .B(_2634_),
    .X(_2647_));
 sky130_fd_sc_hd__nand2_1 _6364_ (.A(\as2650.pc[13] ),
    .B(_2634_),
    .Y(_2648_));
 sky130_fd_sc_hd__nor2_1 _6365_ (.A(_2208_),
    .B(_2645_),
    .Y(_2649_));
 sky130_fd_sc_hd__a31o_1 _6366_ (.A1(_2208_),
    .A2(_2647_),
    .A3(_2648_),
    .B1(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__inv_2 _6367_ (.A(_2645_),
    .Y(_2651_));
 sky130_fd_sc_hd__a221o_1 _6368_ (.A1(\as2650.addr_buff[5] ),
    .A2(_1865_),
    .B1(_1692_),
    .B2(_2651_),
    .C1(_3110_),
    .X(_2652_));
 sky130_fd_sc_hd__a21o_1 _6369_ (.A1(_0888_),
    .A2(_2650_),
    .B1(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__a31o_1 _6370_ (.A1(\as2650.pc[13] ),
    .A2(_3149_),
    .A3(_1699_),
    .B1(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__a31o_1 _6371_ (.A1(_0887_),
    .A2(_2643_),
    .A3(_2644_),
    .B1(_3076_),
    .X(_2655_));
 sky130_fd_sc_hd__a32o_1 _6372_ (.A1(\as2650.pc[13] ),
    .A2(_3149_),
    .A3(_1740_),
    .B1(_2655_),
    .B2(_1618_),
    .X(_2656_));
 sky130_fd_sc_hd__a22o_1 _6373_ (.A1(\as2650.addr_buff[5] ),
    .A2(_1857_),
    .B1(_2611_),
    .B2(\as2650.addr_buff[4] ),
    .X(_2657_));
 sky130_fd_sc_hd__nor2_1 _6374_ (.A(_0891_),
    .B(_2645_),
    .Y(_2658_));
 sky130_fd_sc_hd__a211o_1 _6375_ (.A1(_0891_),
    .A2(_2657_),
    .B1(_2658_),
    .C1(_2158_),
    .X(_2659_));
 sky130_fd_sc_hd__a22o_1 _6376_ (.A1(_0541_),
    .A2(_2226_),
    .B1(_2651_),
    .B2(_0991_),
    .X(_2660_));
 sky130_fd_sc_hd__a31o_1 _6377_ (.A1(_2654_),
    .A2(_2656_),
    .A3(_2659_),
    .B1(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__a21o_1 _6378_ (.A1(_2323_),
    .A2(_2661_),
    .B1(_2393_),
    .X(_2662_));
 sky130_fd_sc_hd__o221a_1 _6379_ (.A1(\as2650.pc[13] ),
    .A2(_2358_),
    .B1(_2646_),
    .B2(_2662_),
    .C1(_1709_),
    .X(_0229_));
 sky130_fd_sc_hd__xnor2_2 _6380_ (.A(\as2650.pc[14] ),
    .B(_2643_),
    .Y(_2663_));
 sky130_fd_sc_hd__xnor2_1 _6381_ (.A(\as2650.pc[14] ),
    .B(_2648_),
    .Y(_2664_));
 sky130_fd_sc_hd__mux2_1 _6382_ (.A0(_2663_),
    .A1(_2664_),
    .S(_2208_),
    .X(_2665_));
 sky130_fd_sc_hd__and2_1 _6383_ (.A(\as2650.pc[14] ),
    .B(_3147_),
    .X(_2666_));
 sky130_fd_sc_hd__o221a_1 _6384_ (.A1(\as2650.addr_buff[6] ),
    .A2(_0892_),
    .B1(_3085_),
    .B2(_2666_),
    .C1(_3098_),
    .X(_2667_));
 sky130_fd_sc_hd__o21a_1 _6385_ (.A1(_1732_),
    .A2(_2663_),
    .B1(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__a211o_1 _6386_ (.A1(_0908_),
    .A2(_2665_),
    .B1(_2668_),
    .C1(_2120_),
    .X(_2669_));
 sky130_fd_sc_hd__and3_1 _6387_ (.A(\as2650.addr_buff[6] ),
    .B(_1857_),
    .C(_0891_),
    .X(_2670_));
 sky130_fd_sc_hd__a211o_1 _6388_ (.A1(_1609_),
    .A2(_2663_),
    .B1(_2670_),
    .C1(_2158_),
    .X(_2671_));
 sky130_fd_sc_hd__a21o_1 _6389_ (.A1(_2669_),
    .A2(_2671_),
    .B1(_2319_),
    .X(_2672_));
 sky130_fd_sc_hd__a31o_1 _6390_ (.A1(\as2650.pc[14] ),
    .A2(_3149_),
    .A3(_3080_),
    .B1(_3076_),
    .X(_2673_));
 sky130_fd_sc_hd__a21o_1 _6391_ (.A1(_0888_),
    .A2(_2663_),
    .B1(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__o221a_1 _6392_ (.A1(_0550_),
    .A2(_1003_),
    .B1(_2663_),
    .B2(_2295_),
    .C1(_2008_),
    .X(_2675_));
 sky130_fd_sc_hd__and2_1 _6393_ (.A(_2674_),
    .B(_2675_),
    .X(_2676_));
 sky130_fd_sc_hd__a221o_1 _6394_ (.A1(_1882_),
    .A2(_2663_),
    .B1(_2672_),
    .B2(_2676_),
    .C1(_2393_),
    .X(_2677_));
 sky130_fd_sc_hd__o211a_1 _6395_ (.A1(\as2650.pc[14] ),
    .A2(_2294_),
    .B1(_2677_),
    .C1(_2515_),
    .X(_0230_));
 sky130_fd_sc_hd__a31o_1 _6396_ (.A1(\as2650.cycle[7] ),
    .A2(_3049_),
    .A3(_1681_),
    .B1(\as2650.halted ),
    .X(_2678_));
 sky130_fd_sc_hd__or4_1 _6397_ (.A(_3039_),
    .B(_0963_),
    .C(_0974_),
    .D(_1012_),
    .X(_2679_));
 sky130_fd_sc_hd__nor2_1 _6398_ (.A(_3292_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__or3b_1 _6399_ (.A(_2678_),
    .B(_2680_),
    .C_N(_1630_),
    .X(_2681_));
 sky130_fd_sc_hd__a22o_1 _6400_ (.A1(_3186_),
    .A2(_3299_),
    .B1(_3229_),
    .B2(_1607_),
    .X(_2682_));
 sky130_fd_sc_hd__o211a_1 _6401_ (.A1(_3186_),
    .A2(_3210_),
    .B1(_1774_),
    .C1(_3252_),
    .X(_2683_));
 sky130_fd_sc_hd__o21ai_1 _6402_ (.A1(_2682_),
    .A2(_2683_),
    .B1(_0969_),
    .Y(_2684_));
 sky130_fd_sc_hd__o21ai_1 _6403_ (.A1(_3193_),
    .A2(_0988_),
    .B1(_3200_),
    .Y(_2685_));
 sky130_fd_sc_hd__nand2_1 _6404_ (.A(_3186_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__a31o_1 _6405_ (.A1(_3067_),
    .A2(_3120_),
    .A3(_3167_),
    .B1(_0643_),
    .X(_2687_));
 sky130_fd_sc_hd__a21o_1 _6406_ (.A1(_0654_),
    .A2(_2687_),
    .B1(_3049_),
    .X(_2688_));
 sky130_fd_sc_hd__and4_1 _6407_ (.A(_1002_),
    .B(_2684_),
    .C(_2686_),
    .D(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__or3b_1 _6408_ (.A(_2681_),
    .B(_0995_),
    .C_N(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__or4_1 _6409_ (.A(_0647_),
    .B(_3216_),
    .C(_3229_),
    .D(_3230_),
    .X(_2691_));
 sky130_fd_sc_hd__or3_1 _6410_ (.A(_3214_),
    .B(_1673_),
    .C(_1009_),
    .X(_2692_));
 sky130_fd_sc_hd__or3_1 _6411_ (.A(_3101_),
    .B(_1609_),
    .C(_1637_),
    .X(_2693_));
 sky130_fd_sc_hd__or4_1 _6412_ (.A(\as2650.cycle[7] ),
    .B(_3088_),
    .C(_3059_),
    .D(_1686_),
    .X(_2694_));
 sky130_fd_sc_hd__and3_1 _6413_ (.A(_3074_),
    .B(_1003_),
    .C(_2128_),
    .X(_2695_));
 sky130_fd_sc_hd__and3_1 _6414_ (.A(_3064_),
    .B(_2694_),
    .C(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__and4b_1 _6415_ (.A_N(_3054_),
    .B(_1662_),
    .C(_1652_),
    .D(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__o2111a_1 _6416_ (.A1(_1687_),
    .A2(_2691_),
    .B1(_2692_),
    .C1(_2693_),
    .D1(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__or3b_1 _6417_ (.A(_0977_),
    .B(_2690_),
    .C_N(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__buf_2 _6418_ (.A(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__clkbuf_4 _6419_ (.A(_1865_),
    .X(_2701_));
 sky130_fd_sc_hd__mux2_1 _6420_ (.A0(_3260_),
    .A1(_3250_),
    .S(_3090_),
    .X(_2702_));
 sky130_fd_sc_hd__or2_1 _6421_ (.A(_0647_),
    .B(_3325_),
    .X(_2703_));
 sky130_fd_sc_hd__o211a_1 _6422_ (.A1(_2701_),
    .A2(_2702_),
    .B1(_2703_),
    .C1(_3103_),
    .X(_2704_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(_0777_),
    .B(_1026_),
    .Y(_2705_));
 sky130_fd_sc_hd__nand2_1 _6424_ (.A(_1028_),
    .B(_0881_),
    .Y(_2706_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(\as2650.carry ),
    .B(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__a211o_1 _6426_ (.A1(_3339_),
    .A2(_1650_),
    .B1(_2707_),
    .C1(_0761_),
    .X(_2708_));
 sky130_fd_sc_hd__inv_2 _6427_ (.A(_2301_),
    .Y(_2709_));
 sky130_fd_sc_hd__o221a_1 _6428_ (.A1(_0760_),
    .A2(_0696_),
    .B1(_2709_),
    .B2(_3331_),
    .C1(_0988_),
    .X(_2710_));
 sky130_fd_sc_hd__a221o_1 _6429_ (.A1(_0985_),
    .A2(_3280_),
    .B1(_2708_),
    .B2(_2710_),
    .C1(_3198_),
    .X(_2711_));
 sky130_fd_sc_hd__o221a_1 _6430_ (.A1(_3029_),
    .A2(_1037_),
    .B1(_2705_),
    .B2(_2711_),
    .C1(_0981_),
    .X(_2712_));
 sky130_fd_sc_hd__a2111o_1 _6431_ (.A1(_3287_),
    .A2(_2270_),
    .B1(_2704_),
    .C1(_2712_),
    .D1(_2700_),
    .X(_2713_));
 sky130_fd_sc_hd__o21ba_1 _6432_ (.A1(_1098_),
    .A2(_3288_),
    .B1_N(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__a211oi_2 _6433_ (.A1(_3361_),
    .A2(_2700_),
    .B1(_2714_),
    .C1(_0921_),
    .Y(_0231_));
 sky130_fd_sc_hd__o2111a_1 _6434_ (.A1(_1687_),
    .A2(_2691_),
    .B1(_2692_),
    .C1(_2688_),
    .D1(_2693_),
    .X(_2715_));
 sky130_fd_sc_hd__and3_1 _6435_ (.A(_1002_),
    .B(_2684_),
    .C(_2686_),
    .X(_2716_));
 sky130_fd_sc_hd__nor2_1 _6436_ (.A(_0977_),
    .B(_2681_),
    .Y(_2717_));
 sky130_fd_sc_hd__or4_1 _6437_ (.A(_3079_),
    .B(_0875_),
    .C(_0878_),
    .D(_0994_),
    .X(_2718_));
 sky130_fd_sc_hd__o31a_1 _6438_ (.A1(_1617_),
    .A2(_3080_),
    .A3(_3363_),
    .B1(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__and4b_1 _6439_ (.A_N(_3054_),
    .B(_3064_),
    .C(_1006_),
    .D(_2695_),
    .X(_2720_));
 sky130_fd_sc_hd__and4b_1 _6440_ (.A_N(_2124_),
    .B(_2717_),
    .C(_2719_),
    .D(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__and3_1 _6441_ (.A(_2715_),
    .B(_2716_),
    .C(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__clkbuf_2 _6442_ (.A(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__mux2_1 _6443_ (.A0(_0303_),
    .A1(_0307_),
    .S(_3091_),
    .X(_2724_));
 sky130_fd_sc_hd__or2_1 _6444_ (.A(_1772_),
    .B(_3389_),
    .X(_2725_));
 sky130_fd_sc_hd__o211a_1 _6445_ (.A1(_2701_),
    .A2(_2724_),
    .B1(_2725_),
    .C1(_1803_),
    .X(_2726_));
 sky130_fd_sc_hd__nor2_2 _6446_ (.A(_3173_),
    .B(_0883_),
    .Y(_2727_));
 sky130_fd_sc_hd__nor2_1 _6447_ (.A(_0946_),
    .B(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__a21o_1 _6448_ (.A1(_3343_),
    .A2(_1650_),
    .B1(_0761_),
    .X(_2729_));
 sky130_fd_sc_hd__o21a_1 _6449_ (.A1(_0760_),
    .A2(_0707_),
    .B1(_0988_),
    .X(_2730_));
 sky130_fd_sc_hd__o221a_1 _6450_ (.A1(_3331_),
    .A2(_2352_),
    .B1(_2728_),
    .B2(_2729_),
    .C1(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__a221o_1 _6451_ (.A1(_0986_),
    .A2(_3287_),
    .B1(_3397_),
    .B2(_0985_),
    .C1(_1019_),
    .X(_2732_));
 sky130_fd_sc_hd__o221a_1 _6452_ (.A1(_3129_),
    .A2(_1037_),
    .B1(_2731_),
    .B2(_2732_),
    .C1(_0981_),
    .X(_2733_));
 sky130_fd_sc_hd__a211o_1 _6453_ (.A1(_3280_),
    .A2(_2270_),
    .B1(_2700_),
    .C1(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__a211o_1 _6454_ (.A1(_3123_),
    .A2(_3401_),
    .B1(_2726_),
    .C1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__o211a_1 _6455_ (.A1(_0659_),
    .A2(_2723_),
    .B1(_2735_),
    .C1(_2515_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _6456_ (.A0(_0342_),
    .A1(_0340_),
    .S(_3091_),
    .X(_2736_));
 sky130_fd_sc_hd__o21a_1 _6457_ (.A1(_2701_),
    .A2(_2736_),
    .B1(_3103_),
    .X(_2737_));
 sky130_fd_sc_hd__o21a_1 _6458_ (.A1(_1772_),
    .A2(_0377_),
    .B1(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__inv_2 _6459_ (.A(\as2650.overflow ),
    .Y(_2739_));
 sky130_fd_sc_hd__nor2_1 _6460_ (.A(_2739_),
    .B(_2727_),
    .Y(_2740_));
 sky130_fd_sc_hd__a21o_1 _6461_ (.A1(_0317_),
    .A2(_1650_),
    .B1(_0761_),
    .X(_2741_));
 sky130_fd_sc_hd__o21a_1 _6462_ (.A1(_0760_),
    .A2(_0712_),
    .B1(_0988_),
    .X(_2742_));
 sky130_fd_sc_hd__o221a_1 _6463_ (.A1(_3331_),
    .A2(_2391_),
    .B1(_2740_),
    .B2(_2741_),
    .C1(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__a221o_1 _6464_ (.A1(_0986_),
    .A2(_3280_),
    .B1(_0354_),
    .B2(_0985_),
    .C1(_1019_),
    .X(_2744_));
 sky130_fd_sc_hd__o221a_1 _6465_ (.A1(_3132_),
    .A2(_1037_),
    .B1(_2743_),
    .B2(_2744_),
    .C1(_0981_),
    .X(_2745_));
 sky130_fd_sc_hd__inv_2 _6466_ (.A(_0345_),
    .Y(_2746_));
 sky130_fd_sc_hd__a221o_1 _6467_ (.A1(_3123_),
    .A2(_2746_),
    .B1(_2270_),
    .B2(_3397_),
    .C1(_2700_),
    .X(_2747_));
 sky130_fd_sc_hd__or3_1 _6468_ (.A(_2738_),
    .B(_2745_),
    .C(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__o211a_1 _6469_ (.A1(_0664_),
    .A2(_2723_),
    .B1(_2748_),
    .C1(_2515_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6470_ (.A0(_0420_),
    .A1(_0403_),
    .S(_3091_),
    .X(_2749_));
 sky130_fd_sc_hd__nand2_1 _6471_ (.A(_2701_),
    .B(_0397_),
    .Y(_2750_));
 sky130_fd_sc_hd__o211a_1 _6472_ (.A1(_2701_),
    .A2(_2749_),
    .B1(_2750_),
    .C1(_1803_),
    .X(_2751_));
 sky130_fd_sc_hd__a21o_1 _6473_ (.A1(\as2650.psl[3] ),
    .A2(_2706_),
    .B1(_0761_),
    .X(_2752_));
 sky130_fd_sc_hd__a21o_1 _6474_ (.A1(\as2650.psu[3] ),
    .A2(_1650_),
    .B1(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__o221a_1 _6475_ (.A1(_0760_),
    .A2(_0718_),
    .B1(_2403_),
    .B2(_3331_),
    .C1(_0988_),
    .X(_2754_));
 sky130_fd_sc_hd__a221o_1 _6476_ (.A1(_0986_),
    .A2(_3397_),
    .B1(_0439_),
    .B2(_0985_),
    .C1(_3198_),
    .X(_2755_));
 sky130_fd_sc_hd__a21o_1 _6477_ (.A1(_2753_),
    .A2(_2754_),
    .B1(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__o211a_1 _6478_ (.A1(_3135_),
    .A2(_1037_),
    .B1(_0981_),
    .C1(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__a221o_1 _6479_ (.A1(_3123_),
    .A2(_0406_),
    .B1(_2270_),
    .B2(_0354_),
    .C1(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__or3_1 _6480_ (.A(_2700_),
    .B(_2751_),
    .C(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__o211a_1 _6481_ (.A1(_0667_),
    .A2(_2723_),
    .B1(_2759_),
    .C1(_2515_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6482_ (.A0(_0477_),
    .A1(_0480_),
    .S(_3091_),
    .X(_2760_));
 sky130_fd_sc_hd__or2_1 _6483_ (.A(_2701_),
    .B(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__o211a_1 _6484_ (.A1(_1772_),
    .A2(_0454_),
    .B1(_2761_),
    .C1(_1803_),
    .X(_2762_));
 sky130_fd_sc_hd__nor2_1 _6485_ (.A(\as2650.psu[4] ),
    .B(_2706_),
    .Y(_2763_));
 sky130_fd_sc_hd__a211o_1 _6486_ (.A1(_3184_),
    .A2(_2706_),
    .B1(_2763_),
    .C1(_0313_),
    .X(_2764_));
 sky130_fd_sc_hd__o211a_1 _6487_ (.A1(_3331_),
    .A2(_2432_),
    .B1(_2764_),
    .C1(_0760_),
    .X(_2765_));
 sky130_fd_sc_hd__o21ai_1 _6488_ (.A1(_0760_),
    .A2(_0724_),
    .B1(_0777_),
    .Y(_2766_));
 sky130_fd_sc_hd__a2bb2o_1 _6489_ (.A1_N(_2765_),
    .A2_N(_2766_),
    .B1(_0986_),
    .B2(_0354_),
    .X(_2767_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(_0461_),
    .A1(_2767_),
    .S(_0876_),
    .X(_2768_));
 sky130_fd_sc_hd__or2_1 _6491_ (.A(_1019_),
    .B(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__a21oi_1 _6492_ (.A1(_0465_),
    .A2(_1019_),
    .B1(_0898_),
    .Y(_2770_));
 sky130_fd_sc_hd__a221o_1 _6493_ (.A1(_3123_),
    .A2(_0463_),
    .B1(_2769_),
    .B2(_2770_),
    .C1(_2700_),
    .X(_2771_));
 sky130_fd_sc_hd__a211o_1 _6494_ (.A1(_0439_),
    .A2(_2270_),
    .B1(_2762_),
    .C1(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__o211a_1 _6495_ (.A1(_0671_),
    .A2(_2723_),
    .B1(_2772_),
    .C1(_2515_),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _6496_ (.A(_3091_),
    .B(_0499_),
    .X(_2773_));
 sky130_fd_sc_hd__a211o_1 _6497_ (.A1(_1710_),
    .A2(_0516_),
    .B1(_2773_),
    .C1(_2701_),
    .X(_2774_));
 sky130_fd_sc_hd__o211a_1 _6498_ (.A1(_1772_),
    .A2(_0535_),
    .B1(_2774_),
    .C1(_1803_),
    .X(_2775_));
 sky130_fd_sc_hd__mux2_1 _6499_ (.A0(\as2650.psl[5] ),
    .A1(\as2650.psu[5] ),
    .S(_2727_),
    .X(_2776_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(_2479_),
    .A1(_2776_),
    .S(_3174_),
    .X(_2777_));
 sky130_fd_sc_hd__mux2_1 _6501_ (.A0(_0731_),
    .A1(_2777_),
    .S(_3181_),
    .X(_2778_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_0777_),
    .B(_0414_),
    .Y(_2779_));
 sky130_fd_sc_hd__a21o_1 _6503_ (.A1(_0777_),
    .A2(_2778_),
    .B1(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__mux2_1 _6504_ (.A0(_0566_),
    .A1(_2780_),
    .S(_0876_),
    .X(_2781_));
 sky130_fd_sc_hd__or2_1 _6505_ (.A(_1019_),
    .B(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__nand2_1 _6506_ (.A(_1046_),
    .B(_1019_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor2_1 _6507_ (.A(_1098_),
    .B(_0507_),
    .Y(_2784_));
 sky130_fd_sc_hd__a311o_1 _6508_ (.A1(_0981_),
    .A2(_2782_),
    .A3(_2783_),
    .B1(_2700_),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a211o_1 _6509_ (.A1(_0461_),
    .A2(_2270_),
    .B1(_2775_),
    .C1(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__buf_4 _6510_ (.A(_3154_),
    .X(_2787_));
 sky130_fd_sc_hd__o211a_1 _6511_ (.A1(_0675_),
    .A2(_2723_),
    .B1(_2786_),
    .C1(_2787_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(_0579_),
    .A1(_0577_),
    .S(_3091_),
    .X(_2788_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(_2701_),
    .B(_0571_),
    .Y(_2789_));
 sky130_fd_sc_hd__o211a_1 _6514_ (.A1(_2701_),
    .A2(_2788_),
    .B1(_2789_),
    .C1(_1803_),
    .X(_2790_));
 sky130_fd_sc_hd__nor2_1 _6515_ (.A(_1098_),
    .B(_0584_),
    .Y(_2791_));
 sky130_fd_sc_hd__mux2_1 _6516_ (.A0(\as2650.psl[6] ),
    .A1(io_out[26]),
    .S(_2727_),
    .X(_2792_));
 sky130_fd_sc_hd__o221a_1 _6517_ (.A1(_0760_),
    .A2(_0736_),
    .B1(_2511_),
    .B2(_3331_),
    .C1(_0988_),
    .X(_2793_));
 sky130_fd_sc_hd__o21ai_1 _6518_ (.A1(_0761_),
    .A2(_2792_),
    .B1(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__o221a_1 _6519_ (.A1(_0876_),
    .A2(_0596_),
    .B1(_0491_),
    .B2(_0777_),
    .C1(_1037_),
    .X(_2795_));
 sky130_fd_sc_hd__nand2_1 _6520_ (.A(_2794_),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__a32o_1 _6521_ (.A1(_0981_),
    .A2(_1023_),
    .A3(_2796_),
    .B1(_0566_),
    .B2(_2270_),
    .X(_2797_));
 sky130_fd_sc_hd__or4_1 _6522_ (.A(_2700_),
    .B(_2790_),
    .C(_2791_),
    .D(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__o211a_1 _6523_ (.A1(_0679_),
    .A2(_2723_),
    .B1(_2798_),
    .C1(_2787_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(_0628_),
    .A1(_0616_),
    .S(_3091_),
    .X(_2799_));
 sky130_fd_sc_hd__or2_1 _6525_ (.A(_1772_),
    .B(_0611_),
    .X(_2800_));
 sky130_fd_sc_hd__o211a_1 _6526_ (.A1(_2701_),
    .A2(_2799_),
    .B1(_2800_),
    .C1(_1803_),
    .X(_2801_));
 sky130_fd_sc_hd__nor2_1 _6527_ (.A(_1098_),
    .B(_0621_),
    .Y(_2802_));
 sky130_fd_sc_hd__mux2_1 _6528_ (.A0(\as2650.psl[7] ),
    .A1(\as2650.psu[7] ),
    .S(_2727_),
    .X(_2803_));
 sky130_fd_sc_hd__or2_1 _6529_ (.A(_3331_),
    .B(_2540_),
    .X(_2804_));
 sky130_fd_sc_hd__o221a_1 _6530_ (.A1(_0760_),
    .A2(_1315_),
    .B1(_2803_),
    .B2(_0761_),
    .C1(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__o21ai_1 _6531_ (.A1(_0878_),
    .A2(_2805_),
    .B1(_1043_),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_1 _6532_ (.A(_1020_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__a221o_1 _6533_ (.A1(_3271_),
    .A2(_2270_),
    .B1(_2807_),
    .B2(_0981_),
    .C1(_2700_),
    .X(_2808_));
 sky130_fd_sc_hd__or3_1 _6534_ (.A(_2801_),
    .B(_2802_),
    .C(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__o211a_1 _6535_ (.A1(_0684_),
    .A2(_2723_),
    .B1(_2809_),
    .C1(_2787_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6536_ (.A0(_0636_),
    .A1(\as2650.stack[6][0] ),
    .S(_0701_),
    .X(_2810_));
 sky130_fd_sc_hd__or3_4 _6537_ (.A(_0700_),
    .B(_0316_),
    .C(_0725_),
    .X(_2811_));
 sky130_fd_sc_hd__mux2_1 _6538_ (.A0(_0634_),
    .A1(_2810_),
    .S(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__clkbuf_1 _6539_ (.A(_2812_),
    .X(_0239_));
 sky130_fd_sc_hd__nor3_4 _6540_ (.A(_0700_),
    .B(_0316_),
    .C(_0697_),
    .Y(_2813_));
 sky130_fd_sc_hd__nor3_4 _6541_ (.A(_0700_),
    .B(_0329_),
    .C(_0932_),
    .Y(_2814_));
 sky130_fd_sc_hd__or2_1 _6542_ (.A(\as2650.stack[6][1] ),
    .B(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__o21a_1 _6543_ (.A1(_0661_),
    .A2(_0701_),
    .B1(_2811_),
    .X(_2816_));
 sky130_fd_sc_hd__a22o_1 _6544_ (.A1(_0659_),
    .A2(_2813_),
    .B1(_2815_),
    .B2(_2816_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _6545_ (.A(\as2650.stack[6][2] ),
    .B(_2814_),
    .X(_2817_));
 sky130_fd_sc_hd__a21oi_1 _6546_ (.A1(_1484_),
    .A2(_2814_),
    .B1(_2813_),
    .Y(_2818_));
 sky130_fd_sc_hd__a22o_1 _6547_ (.A1(_0664_),
    .A2(_2813_),
    .B1(_2817_),
    .B2(_2818_),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _6548_ (.A(\as2650.stack[6][3] ),
    .B(_2814_),
    .X(_2819_));
 sky130_fd_sc_hd__a21oi_1 _6549_ (.A1(_1487_),
    .A2(_2814_),
    .B1(_2813_),
    .Y(_2820_));
 sky130_fd_sc_hd__a22o_1 _6550_ (.A1(_0667_),
    .A2(_2813_),
    .B1(_2819_),
    .B2(_2820_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _6551_ (.A(\as2650.stack[6][4] ),
    .B(_2814_),
    .X(_2821_));
 sky130_fd_sc_hd__a21oi_1 _6552_ (.A1(_1490_),
    .A2(_2814_),
    .B1(_2813_),
    .Y(_2822_));
 sky130_fd_sc_hd__a22o_1 _6553_ (.A1(_0671_),
    .A2(_2813_),
    .B1(_2821_),
    .B2(_2822_),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _6554_ (.A(\as2650.stack[6][5] ),
    .B(_2814_),
    .X(_2823_));
 sky130_fd_sc_hd__o21a_1 _6555_ (.A1(_0676_),
    .A2(_0701_),
    .B1(_2811_),
    .X(_2824_));
 sky130_fd_sc_hd__a22o_1 _6556_ (.A1(_0675_),
    .A2(_2813_),
    .B1(_2823_),
    .B2(_2824_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6557_ (.A0(_0681_),
    .A1(\as2650.stack[6][6] ),
    .S(_0701_),
    .X(_2825_));
 sky130_fd_sc_hd__mux2_1 _6558_ (.A0(_0679_),
    .A1(_2825_),
    .S(_2811_),
    .X(_2826_));
 sky130_fd_sc_hd__clkbuf_1 _6559_ (.A(_2826_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _6560_ (.A(\as2650.stack[6][7] ),
    .B(_2814_),
    .X(_2827_));
 sky130_fd_sc_hd__o21a_1 _6561_ (.A1(_0685_),
    .A2(_0701_),
    .B1(_2811_),
    .X(_2828_));
 sky130_fd_sc_hd__a22o_1 _6562_ (.A1(_0684_),
    .A2(_2813_),
    .B1(_2827_),
    .B2(_2828_),
    .X(_0246_));
 sky130_fd_sc_hd__or3_4 _6563_ (.A(_0700_),
    .B(_0316_),
    .C(_0649_),
    .X(_2829_));
 sky130_fd_sc_hd__mux2_1 _6564_ (.A0(_0636_),
    .A1(\as2650.stack[7][0] ),
    .S(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _6565_ (.A0(_0634_),
    .A1(_2830_),
    .S(_1283_),
    .X(_2831_));
 sky130_fd_sc_hd__clkbuf_1 _6566_ (.A(_2831_),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_4 _6567_ (.A(_0697_),
    .B(_1281_),
    .Y(_2832_));
 sky130_fd_sc_hd__nor3_4 _6568_ (.A(_0700_),
    .B(_0316_),
    .C(_0932_),
    .Y(_2833_));
 sky130_fd_sc_hd__or2_1 _6569_ (.A(\as2650.stack[7][1] ),
    .B(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__o21a_1 _6570_ (.A1(_0661_),
    .A2(_2829_),
    .B1(_1283_),
    .X(_2835_));
 sky130_fd_sc_hd__a22o_1 _6571_ (.A1(_0659_),
    .A2(_2832_),
    .B1(_2834_),
    .B2(_2835_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _6572_ (.A(\as2650.stack[7][2] ),
    .B(_2833_),
    .X(_2836_));
 sky130_fd_sc_hd__a21oi_1 _6573_ (.A1(_1484_),
    .A2(_2833_),
    .B1(_2832_),
    .Y(_2837_));
 sky130_fd_sc_hd__a22o_1 _6574_ (.A1(_0664_),
    .A2(_2832_),
    .B1(_2836_),
    .B2(_2837_),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _6575_ (.A(\as2650.stack[7][3] ),
    .B(_2833_),
    .X(_2838_));
 sky130_fd_sc_hd__a21oi_1 _6576_ (.A1(_1487_),
    .A2(_2833_),
    .B1(_2832_),
    .Y(_2839_));
 sky130_fd_sc_hd__a22o_1 _6577_ (.A1(_0667_),
    .A2(_2832_),
    .B1(_2838_),
    .B2(_2839_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _6578_ (.A(\as2650.stack[7][4] ),
    .B(_2833_),
    .X(_2840_));
 sky130_fd_sc_hd__a21oi_1 _6579_ (.A1(_1490_),
    .A2(_2833_),
    .B1(_2832_),
    .Y(_2841_));
 sky130_fd_sc_hd__a22o_1 _6580_ (.A1(_0671_),
    .A2(_2832_),
    .B1(_2840_),
    .B2(_2841_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _6581_ (.A(\as2650.stack[7][5] ),
    .B(_2833_),
    .X(_2842_));
 sky130_fd_sc_hd__o21a_1 _6582_ (.A1(_0676_),
    .A2(_2829_),
    .B1(_1283_),
    .X(_2843_));
 sky130_fd_sc_hd__a22o_1 _6583_ (.A1(_0675_),
    .A2(_2832_),
    .B1(_2842_),
    .B2(_2843_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _6584_ (.A(\as2650.stack[7][6] ),
    .B(_2833_),
    .X(_2844_));
 sky130_fd_sc_hd__o21a_1 _6585_ (.A1(_0681_),
    .A2(_2829_),
    .B1(_1283_),
    .X(_2845_));
 sky130_fd_sc_hd__a22o_1 _6586_ (.A1(_0679_),
    .A2(_2832_),
    .B1(_2844_),
    .B2(_2845_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _6587_ (.A(\as2650.stack[7][7] ),
    .B(_2833_),
    .X(_2846_));
 sky130_fd_sc_hd__o21a_1 _6588_ (.A1(_0685_),
    .A2(_2829_),
    .B1(_1283_),
    .X(_2847_));
 sky130_fd_sc_hd__a22o_1 _6589_ (.A1(_0684_),
    .A2(_2832_),
    .B1(_2846_),
    .B2(_2847_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_4 _6590_ (.A(_2811_),
    .B(_2829_),
    .Y(_2848_));
 sky130_fd_sc_hd__mux2_1 _6591_ (.A0(\as2650.stack[7][8] ),
    .A1(_0699_),
    .S(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__clkbuf_1 _6592_ (.A(_2849_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _6593_ (.A0(\as2650.stack[7][9] ),
    .A1(_0709_),
    .S(_2848_),
    .X(_2850_));
 sky130_fd_sc_hd__clkbuf_1 _6594_ (.A(_2850_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _6595_ (.A0(\as2650.stack[7][10] ),
    .A1(_0715_),
    .S(_2848_),
    .X(_2851_));
 sky130_fd_sc_hd__clkbuf_1 _6596_ (.A(_2851_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _6597_ (.A0(\as2650.stack[7][11] ),
    .A1(_0721_),
    .S(_2848_),
    .X(_2852_));
 sky130_fd_sc_hd__clkbuf_1 _6598_ (.A(_2852_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _6599_ (.A0(\as2650.stack[7][12] ),
    .A1(_0728_),
    .S(_2848_),
    .X(_2853_));
 sky130_fd_sc_hd__clkbuf_1 _6600_ (.A(_2853_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _6601_ (.A0(\as2650.stack[7][13] ),
    .A1(_0733_),
    .S(_2848_),
    .X(_2854_));
 sky130_fd_sc_hd__clkbuf_1 _6602_ (.A(_2854_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _6603_ (.A0(\as2650.stack[7][14] ),
    .A1(_0738_),
    .S(_2848_),
    .X(_2855_));
 sky130_fd_sc_hd__clkbuf_1 _6604_ (.A(_2855_),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_2 _6605_ (.A(_3153_),
    .B(_3364_),
    .Y(_2856_));
 sky130_fd_sc_hd__nor2_4 _6606_ (.A(_1010_),
    .B(_3234_),
    .Y(_2857_));
 sky130_fd_sc_hd__nor2_4 _6607_ (.A(_2856_),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__nor3_4 _6608_ (.A(_3330_),
    .B(_3165_),
    .C(_3363_),
    .Y(_2859_));
 sky130_fd_sc_hd__a32o_1 _6609_ (.A1(_0634_),
    .A2(_2859_),
    .A3(_0696_),
    .B1(_2857_),
    .B2(_3329_),
    .X(_2860_));
 sky130_fd_sc_hd__a21o_1 _6610_ (.A1(\as2650.r123[1][0] ),
    .A2(_2858_),
    .B1(_2860_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_4 _6611_ (.A(_2859_),
    .X(_2861_));
 sky130_fd_sc_hd__a22o_1 _6612_ (.A1(_0312_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][1] ),
    .X(_2862_));
 sky130_fd_sc_hd__a21o_1 _6613_ (.A1(_2861_),
    .A2(_1125_),
    .B1(_2862_),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _6614_ (.A1(_0378_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][2] ),
    .X(_2863_));
 sky130_fd_sc_hd__a21o_1 _6615_ (.A1(_2861_),
    .A2(_1135_),
    .B1(_2863_),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _6616_ (.A1(_0424_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][3] ),
    .X(_2864_));
 sky130_fd_sc_hd__a21o_1 _6617_ (.A1(_2861_),
    .A2(_1147_),
    .B1(_2864_),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _6618_ (.A1(_0483_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][4] ),
    .X(_2865_));
 sky130_fd_sc_hd__a21o_1 _6619_ (.A1(_2861_),
    .A2(_1170_),
    .B1(_2865_),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _6620_ (.A1(_0536_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][5] ),
    .X(_2866_));
 sky130_fd_sc_hd__a21o_1 _6621_ (.A1(_2861_),
    .A2(_1196_),
    .B1(_2866_),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _6622_ (.A1(_0592_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][6] ),
    .X(_2867_));
 sky130_fd_sc_hd__a21o_1 _6623_ (.A1(_2861_),
    .A2(_1230_),
    .B1(_2867_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _6624_ (.A1(_0631_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(\as2650.r123[1][7] ),
    .X(_2868_));
 sky130_fd_sc_hd__a21o_1 _6625_ (.A1(_2861_),
    .A2(_1268_),
    .B1(_2868_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_4 _6626_ (.A(_3073_),
    .B(_3234_),
    .Y(_2869_));
 sky130_fd_sc_hd__nor2_2 _6627_ (.A(_2856_),
    .B(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__a22o_1 _6628_ (.A1(_2861_),
    .A2(_1337_),
    .B1(_2870_),
    .B2(\as2650.r123[2][0] ),
    .X(_2871_));
 sky130_fd_sc_hd__a21o_1 _6629_ (.A1(_3329_),
    .A2(_2869_),
    .B1(_2871_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _6630_ (.A1(_2859_),
    .A2(_1369_),
    .B1(_2870_),
    .B2(\as2650.r123[2][1] ),
    .X(_2872_));
 sky130_fd_sc_hd__a21o_1 _6631_ (.A1(_0312_),
    .A2(_2869_),
    .B1(_2872_),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _6632_ (.A1(_2859_),
    .A2(_1402_),
    .B1(_2870_),
    .B2(\as2650.r123[2][2] ),
    .X(_2873_));
 sky130_fd_sc_hd__a21o_1 _6633_ (.A1(_0378_),
    .A2(_2869_),
    .B1(_2873_),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _6634_ (.A1(_2859_),
    .A2(_1427_),
    .B1(_2870_),
    .B2(\as2650.r123[2][3] ),
    .X(_2874_));
 sky130_fd_sc_hd__a21o_1 _6635_ (.A1(_0424_),
    .A2(_2869_),
    .B1(_2874_),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _6636_ (.A1(_2859_),
    .A2(_1446_),
    .B1(_2870_),
    .B2(\as2650.r123[2][4] ),
    .X(_2875_));
 sky130_fd_sc_hd__a21o_1 _6637_ (.A1(_0483_),
    .A2(_2869_),
    .B1(_2875_),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _6638_ (.A1(_2859_),
    .A2(_1460_),
    .B1(_2870_),
    .B2(\as2650.r123[2][5] ),
    .X(_2876_));
 sky130_fd_sc_hd__a21o_1 _6639_ (.A1(_0536_),
    .A2(_2869_),
    .B1(_2876_),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _6640_ (.A1(_0592_),
    .A2(_2869_),
    .B1(_2870_),
    .B2(\as2650.r123[2][6] ),
    .X(_2877_));
 sky130_fd_sc_hd__a21o_1 _6641_ (.A1(_2861_),
    .A2(_1471_),
    .B1(_2877_),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _6642_ (.A1(_0631_),
    .A2(_2869_),
    .B1(_2870_),
    .B2(\as2650.r123[2][7] ),
    .X(_2878_));
 sky130_fd_sc_hd__a21o_1 _6643_ (.A1(_2861_),
    .A2(_1475_),
    .B1(_2878_),
    .X(_0277_));
 sky130_fd_sc_hd__o211a_1 _6644_ (.A1(_3206_),
    .A2(_0980_),
    .B1(_1003_),
    .C1(_2128_),
    .X(_2879_));
 sky130_fd_sc_hd__o2111a_1 _6645_ (.A1(_0691_),
    .A2(_1000_),
    .B1(_1612_),
    .C1(_2879_),
    .D1(_1653_),
    .X(_2880_));
 sky130_fd_sc_hd__nor2_1 _6646_ (.A(_2126_),
    .B(_2678_),
    .Y(_2881_));
 sky130_fd_sc_hd__and4_1 _6647_ (.A(_1603_),
    .B(_2693_),
    .C(_2880_),
    .D(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__buf_4 _6648_ (.A(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__buf_2 _6649_ (.A(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__nor2_1 _6650_ (.A(_0983_),
    .B(_3210_),
    .Y(_2885_));
 sky130_fd_sc_hd__buf_4 _6651_ (.A(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__mux2_2 _6652_ (.A0(_3244_),
    .A1(_3361_),
    .S(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__o21ai_1 _6653_ (.A1(io_out[0]),
    .A2(_2883_),
    .B1(_1562_),
    .Y(_2888_));
 sky130_fd_sc_hd__a21oi_1 _6654_ (.A1(_2884_),
    .A2(_2887_),
    .B1(_2888_),
    .Y(_0278_));
 sky130_fd_sc_hd__mux2_1 _6655_ (.A0(_3280_),
    .A1(_3391_),
    .S(_2886_),
    .X(_2889_));
 sky130_fd_sc_hd__inv_2 _6656_ (.A(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__nand2_1 _6657_ (.A(_2884_),
    .B(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__o211a_1 _6658_ (.A1(io_out[1]),
    .A2(_2884_),
    .B1(_2891_),
    .C1(_2787_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _6659_ (.A0(_3397_),
    .A1(_0326_),
    .S(_2886_),
    .X(_2892_));
 sky130_fd_sc_hd__inv_2 _6660_ (.A(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__nand2_1 _6661_ (.A(_2884_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__o211a_1 _6662_ (.A1(io_out[2]),
    .A2(_2884_),
    .B1(_2894_),
    .C1(_2787_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _6663_ (.A0(_0354_),
    .A1(_0417_),
    .S(_2885_),
    .X(_2895_));
 sky130_fd_sc_hd__inv_2 _6664_ (.A(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__nand2_1 _6665_ (.A(_2883_),
    .B(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__o211a_1 _6666_ (.A1(io_out[3]),
    .A2(_2884_),
    .B1(_2897_),
    .C1(_2787_),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _6667_ (.A(_0671_),
    .B(_2886_),
    .Y(_2898_));
 sky130_fd_sc_hd__o211ai_4 _6668_ (.A1(_0414_),
    .A2(_2886_),
    .B1(_2898_),
    .C1(_2883_),
    .Y(_2899_));
 sky130_fd_sc_hd__o211a_1 _6669_ (.A1(io_out[4]),
    .A2(_2884_),
    .B1(_2899_),
    .C1(_2787_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _6670_ (.A(_0675_),
    .B(_2886_),
    .Y(_2900_));
 sky130_fd_sc_hd__o211ai_4 _6671_ (.A1(_0491_),
    .A2(_2886_),
    .B1(_2900_),
    .C1(_2883_),
    .Y(_2901_));
 sky130_fd_sc_hd__o211a_1 _6672_ (.A1(io_out[5]),
    .A2(_2884_),
    .B1(_2901_),
    .C1(_2787_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _6673_ (.A(_0679_),
    .B(_2886_),
    .Y(_2902_));
 sky130_fd_sc_hd__o211ai_4 _6674_ (.A1(_0504_),
    .A2(_2886_),
    .B1(_2902_),
    .C1(_2883_),
    .Y(_2903_));
 sky130_fd_sc_hd__o211a_1 _6675_ (.A1(io_out[6]),
    .A2(_2884_),
    .B1(_2903_),
    .C1(_2787_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_2 _6676_ (.A0(_0596_),
    .A1(_0866_),
    .S(_2886_),
    .X(_2904_));
 sky130_fd_sc_hd__o21ai_1 _6677_ (.A1(io_out[7]),
    .A2(_2883_),
    .B1(_1562_),
    .Y(_2905_));
 sky130_fd_sc_hd__a21oi_1 _6678_ (.A1(_2884_),
    .A2(_2904_),
    .B1(_2905_),
    .Y(_0285_));
 sky130_fd_sc_hd__mux2_1 _6679_ (.A0(_1618_),
    .A1(_3135_),
    .S(_1097_),
    .X(_2906_));
 sky130_fd_sc_hd__clkbuf_1 _6680_ (.A(_2906_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _6681_ (.A0(_1018_),
    .A1(_3137_),
    .S(_1097_),
    .X(_2907_));
 sky130_fd_sc_hd__clkbuf_1 _6682_ (.A(_2907_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _6683_ (.A(_0983_),
    .B(_3079_),
    .Y(_2908_));
 sky130_fd_sc_hd__or3b_1 _6684_ (.A(_0902_),
    .B(_1630_),
    .C_N(_0895_),
    .X(_2909_));
 sky130_fd_sc_hd__and4_1 _6685_ (.A(_1657_),
    .B(_1652_),
    .C(_1705_),
    .D(_2909_),
    .X(_2910_));
 sky130_fd_sc_hd__o211a_1 _6686_ (.A1(_3227_),
    .A2(_3197_),
    .B1(_1003_),
    .C1(_1011_),
    .X(_2911_));
 sky130_fd_sc_hd__and3_1 _6687_ (.A(_1093_),
    .B(_3052_),
    .C(_1009_),
    .X(_2912_));
 sky130_fd_sc_hd__o211a_1 _6688_ (.A1(_3107_),
    .A2(_1602_),
    .B1(_2911_),
    .C1(_2912_),
    .X(_2913_));
 sky130_fd_sc_hd__and3_1 _6689_ (.A(_0999_),
    .B(_2910_),
    .C(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a211o_1 _6690_ (.A1(\as2650.psl[3] ),
    .A2(_0690_),
    .B1(_0876_),
    .C1(_1617_),
    .X(_2915_));
 sky130_fd_sc_hd__and3_1 _6691_ (.A(_1605_),
    .B(_1646_),
    .C(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__a21o_1 _6692_ (.A1(\as2650.psl[3] ),
    .A2(_2908_),
    .B1(_3263_),
    .X(_2917_));
 sky130_fd_sc_hd__and4_1 _6693_ (.A(_2151_),
    .B(_2914_),
    .C(_2916_),
    .D(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__o31a_1 _6694_ (.A1(_3140_),
    .A2(_0878_),
    .A3(_2908_),
    .B1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__a21o_1 _6695_ (.A1(_0513_),
    .A2(_0691_),
    .B1(_1044_),
    .X(_2920_));
 sky130_fd_sc_hd__a31o_1 _6696_ (.A1(_0777_),
    .A2(_2194_),
    .A3(_2920_),
    .B1(_2779_),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _6697_ (.A0(_0566_),
    .A1(_2921_),
    .S(_0876_),
    .X(_2922_));
 sky130_fd_sc_hd__and2_1 _6698_ (.A(_1018_),
    .B(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__a21bo_1 _6699_ (.A1(_0970_),
    .A2(_0454_),
    .B1_N(_2919_),
    .X(_2924_));
 sky130_fd_sc_hd__o221a_1 _6700_ (.A1(\as2650.psl[5] ),
    .A2(_2919_),
    .B1(_2923_),
    .B2(_2924_),
    .C1(_1786_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _6701_ (.A0(_0595_),
    .A1(_0596_),
    .S(_3292_),
    .X(_2925_));
 sky130_fd_sc_hd__o21ai_1 _6702_ (.A1(_3202_),
    .A2(_0461_),
    .B1(_0529_),
    .Y(_2926_));
 sky130_fd_sc_hd__nand2_1 _6703_ (.A(_2926_),
    .B(_0535_),
    .Y(_2927_));
 sky130_fd_sc_hd__or2_1 _6704_ (.A(_3308_),
    .B(_3325_),
    .X(_2928_));
 sky130_fd_sc_hd__o21a_1 _6705_ (.A1(_3385_),
    .A2(_2928_),
    .B1(_3387_),
    .X(_2929_));
 sky130_fd_sc_hd__a21oi_1 _6706_ (.A1(_3389_),
    .A2(_2928_),
    .B1(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__mux2_1 _6707_ (.A0(\as2650.holding_reg[2] ),
    .A1(_3397_),
    .S(_3292_),
    .X(_2931_));
 sky130_fd_sc_hd__o21ba_1 _6708_ (.A1(_2931_),
    .A2(_2930_),
    .B1_N(_0377_),
    .X(_2932_));
 sky130_fd_sc_hd__a221o_1 _6709_ (.A1(_0391_),
    .A2(_0397_),
    .B1(_2930_),
    .B2(_2931_),
    .C1(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__o22a_1 _6710_ (.A1(_0391_),
    .A2(_0397_),
    .B1(_0449_),
    .B2(_0453_),
    .X(_2934_));
 sky130_fd_sc_hd__a2bb2o_1 _6711_ (.A1_N(_0435_),
    .A2_N(_0454_),
    .B1(_2933_),
    .B2(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__nor2_1 _6712_ (.A(_2926_),
    .B(_0535_),
    .Y(_2936_));
 sky130_fd_sc_hd__a21oi_1 _6713_ (.A1(_2927_),
    .A2(_2935_),
    .B1(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__nor2_1 _6714_ (.A(_0565_),
    .B(_0571_),
    .Y(_2938_));
 sky130_fd_sc_hd__nand2_1 _6715_ (.A(_0565_),
    .B(_0571_),
    .Y(_2939_));
 sky130_fd_sc_hd__o221a_1 _6716_ (.A1(_0611_),
    .A2(_2925_),
    .B1(_2937_),
    .B2(_2938_),
    .C1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__and2_1 _6717_ (.A(_0611_),
    .B(_2925_),
    .X(_2941_));
 sky130_fd_sc_hd__o31a_1 _6718_ (.A1(_3029_),
    .A2(_0878_),
    .A3(_2908_),
    .B1(_2918_),
    .X(_2942_));
 sky130_fd_sc_hd__a21o_1 _6719_ (.A1(_3262_),
    .A2(_0907_),
    .B1(_1044_),
    .X(_2943_));
 sky130_fd_sc_hd__nand3_1 _6720_ (.A(_0777_),
    .B(_2173_),
    .C(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21oi_1 _6721_ (.A1(_0986_),
    .A2(_3271_),
    .B1(_0985_),
    .Y(_2945_));
 sky130_fd_sc_hd__a221o_1 _6722_ (.A1(_0985_),
    .A2(_3244_),
    .B1(_2944_),
    .B2(_2945_),
    .C1(_0970_),
    .X(_2946_));
 sky130_fd_sc_hd__o311a_1 _6723_ (.A1(_1018_),
    .A2(_2940_),
    .A3(_2941_),
    .B1(_2942_),
    .C1(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__o21ai_1 _6724_ (.A1(\as2650.carry ),
    .A2(_2942_),
    .B1(_1786_),
    .Y(_2948_));
 sky130_fd_sc_hd__nor2_1 _6725_ (.A(_2947_),
    .B(_2948_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _6726_ (.A(_0317_),
    .B(_3346_),
    .Y(_2949_));
 sky130_fd_sc_hd__nand2_1 _6727_ (.A(_1079_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__mux2_1 _6728_ (.A0(_0326_),
    .A1(_2950_),
    .S(_0653_),
    .X(_2951_));
 sky130_fd_sc_hd__a21o_1 _6729_ (.A1(_3132_),
    .A2(_0916_),
    .B1(_0691_),
    .X(_2952_));
 sky130_fd_sc_hd__o31a_1 _6730_ (.A1(_3330_),
    .A2(_0313_),
    .A3(_2951_),
    .B1(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__nor2_1 _6731_ (.A(_2144_),
    .B(_0990_),
    .Y(_2954_));
 sky130_fd_sc_hd__o221a_1 _6732_ (.A1(_0990_),
    .A2(_2953_),
    .B1(_2954_),
    .B2(_3338_),
    .C1(_0972_),
    .X(_2955_));
 sky130_fd_sc_hd__a21oi_1 _6733_ (.A1(_1618_),
    .A2(_2950_),
    .B1(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__nand2_1 _6734_ (.A(_3079_),
    .B(_0991_),
    .Y(_2957_));
 sky130_fd_sc_hd__nor2_1 _6735_ (.A(_0992_),
    .B(_2226_),
    .Y(_2958_));
 sky130_fd_sc_hd__inv_2 _6736_ (.A(_2141_),
    .Y(_2959_));
 sky130_fd_sc_hd__o221a_1 _6737_ (.A1(_1872_),
    .A2(_2285_),
    .B1(_2958_),
    .B2(_0887_),
    .C1(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__or4_1 _6738_ (.A(_1617_),
    .B(_0875_),
    .C(_0878_),
    .D(_0886_),
    .X(_2961_));
 sky130_fd_sc_hd__o22a_1 _6739_ (.A1(_1640_),
    .A2(_2435_),
    .B1(_0904_),
    .B2(_2957_),
    .X(_2962_));
 sky130_fd_sc_hd__a31o_1 _6740_ (.A1(_0972_),
    .A2(_3181_),
    .A3(_1649_),
    .B1(_3158_),
    .X(_2963_));
 sky130_fd_sc_hd__o221a_1 _6741_ (.A1(_3040_),
    .A2(_3045_),
    .B1(_3292_),
    .B2(_3196_),
    .C1(_0759_),
    .X(_2964_));
 sky130_fd_sc_hd__a21oi_1 _6742_ (.A1(_3323_),
    .A2(_1008_),
    .B1(_0646_),
    .Y(_2965_));
 sky130_fd_sc_hd__a31oi_1 _6743_ (.A1(_3227_),
    .A2(_0646_),
    .A3(_0644_),
    .B1(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__o221a_1 _6744_ (.A1(_3227_),
    .A2(_0987_),
    .B1(_1695_),
    .B2(_2131_),
    .C1(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__o211a_1 _6745_ (.A1(_0902_),
    .A2(_1044_),
    .B1(_2964_),
    .C1(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__and3_1 _6746_ (.A(_1652_),
    .B(_2963_),
    .C(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__and4bb_1 _6747_ (.A_N(_2287_),
    .B_N(_2280_),
    .C(_2962_),
    .D(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__and3_1 _6748_ (.A(_2960_),
    .B(_2961_),
    .C(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__o21a_1 _6749_ (.A1(_3132_),
    .A2(_2957_),
    .B1(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__mux2_1 _6750_ (.A0(_0700_),
    .A1(_2956_),
    .S(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__nor2_1 _6751_ (.A(_1629_),
    .B(_2973_),
    .Y(_0290_));
 sky130_fd_sc_hd__and2_1 _6752_ (.A(_3341_),
    .B(_3344_),
    .X(_2974_));
 sky130_fd_sc_hd__nand2_1 _6753_ (.A(_3342_),
    .B(_0316_),
    .Y(_2975_));
 sky130_fd_sc_hd__mux2_1 _6754_ (.A0(_3391_),
    .A1(_2974_),
    .S(_0653_),
    .X(_2976_));
 sky130_fd_sc_hd__or3_1 _6755_ (.A(_3159_),
    .B(_0313_),
    .C(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__o211a_1 _6756_ (.A1(_0690_),
    .A2(_0916_),
    .B1(_2180_),
    .C1(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__o221a_1 _6757_ (.A1(_2975_),
    .A2(_2954_),
    .B1(_2978_),
    .B2(_0990_),
    .C1(_0972_),
    .X(_2979_));
 sky130_fd_sc_hd__a21o_1 _6758_ (.A1(_1618_),
    .A2(_2974_),
    .B1(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__o21a_1 _6759_ (.A1(_3129_),
    .A2(_2957_),
    .B1(_2971_),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _6760_ (.A0(_3343_),
    .A1(_2980_),
    .S(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__and2_1 _6761_ (.A(_3154_),
    .B(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__clkbuf_1 _6762_ (.A(_2983_),
    .X(_0291_));
 sky130_fd_sc_hd__or3_1 _6763_ (.A(_0313_),
    .B(_0653_),
    .C(_2295_),
    .X(_2984_));
 sky130_fd_sc_hd__o311a_1 _6764_ (.A1(_3071_),
    .A2(_3292_),
    .A3(_3173_),
    .B1(_0691_),
    .C1(_3262_),
    .X(_2985_));
 sky130_fd_sc_hd__a31o_1 _6765_ (.A1(_3029_),
    .A2(_3080_),
    .A3(_0916_),
    .B1(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__a32o_1 _6766_ (.A1(_3348_),
    .A2(_2957_),
    .A3(_2984_),
    .B1(_2986_),
    .B2(_0991_),
    .X(_2987_));
 sky130_fd_sc_hd__o21a_1 _6767_ (.A1(_3029_),
    .A2(_2957_),
    .B1(_2971_),
    .X(_2988_));
 sky130_fd_sc_hd__mux2_1 _6768_ (.A0(_3339_),
    .A1(_2987_),
    .S(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__and2_1 _6769_ (.A(_3154_),
    .B(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__clkbuf_1 _6770_ (.A(_2990_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_1 _6771_ (.A(_0611_),
    .B(_2925_),
    .Y(_2991_));
 sky130_fd_sc_hd__or2_1 _6772_ (.A(_2991_),
    .B(_2941_),
    .X(_2992_));
 sky130_fd_sc_hd__a21o_1 _6773_ (.A1(_0326_),
    .A2(_0907_),
    .B1(_1044_),
    .X(_2993_));
 sky130_fd_sc_hd__o221a_1 _6774_ (.A1(_1617_),
    .A2(_0988_),
    .B1(_2908_),
    .B2(_3132_),
    .C1(_1605_),
    .X(_2994_));
 sky130_fd_sc_hd__nand3_1 _6775_ (.A(_0885_),
    .B(_2914_),
    .C(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__a31o_1 _6776_ (.A1(_0983_),
    .A2(_2184_),
    .A3(_2993_),
    .B1(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__a31o_1 _6777_ (.A1(_0970_),
    .A2(_0603_),
    .A3(_2992_),
    .B1(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__nand2_1 _6778_ (.A(_2739_),
    .B(_2995_),
    .Y(_2998_));
 sky130_fd_sc_hd__and3_1 _6779_ (.A(_3154_),
    .B(_2997_),
    .C(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__clkbuf_1 _6780_ (.A(_2999_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _6781_ (.A(_3137_),
    .B(_0908_),
    .Y(_3000_));
 sky130_fd_sc_hd__nor3_1 _6782_ (.A(_3079_),
    .B(_3173_),
    .C(_0880_),
    .Y(_3001_));
 sky130_fd_sc_hd__nor2_1 _6783_ (.A(_1010_),
    .B(_0691_),
    .Y(_3002_));
 sky130_fd_sc_hd__a211o_1 _6784_ (.A1(_0892_),
    .A2(_0895_),
    .B1(_3119_),
    .C1(\as2650.halted ),
    .X(_3003_));
 sky130_fd_sc_hd__or4_1 _6785_ (.A(_3001_),
    .B(_0979_),
    .C(_3002_),
    .D(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__a21o_2 _6786_ (.A1(_0908_),
    .A2(_0998_),
    .B1(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__o21ai_1 _6787_ (.A1(_3000_),
    .A2(_3005_),
    .B1(_3163_),
    .Y(_3006_));
 sky130_fd_sc_hd__o31a_1 _6788_ (.A1(_0465_),
    .A2(_0908_),
    .A3(_0896_),
    .B1(_2190_),
    .X(_3007_));
 sky130_fd_sc_hd__or2_1 _6789_ (.A(_3005_),
    .B(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__a21oi_1 _6790_ (.A1(_3006_),
    .A2(_3008_),
    .B1(_1629_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _6791_ (.A(_3135_),
    .B(_0908_),
    .Y(_3009_));
 sky130_fd_sc_hd__o21ai_1 _6792_ (.A1(_3009_),
    .A2(_3005_),
    .B1(\as2650.psl[3] ),
    .Y(_3010_));
 sky130_fd_sc_hd__o31a_1 _6793_ (.A1(_0818_),
    .A2(_0908_),
    .A3(_0896_),
    .B1(_2186_),
    .X(_3011_));
 sky130_fd_sc_hd__or2_1 _6794_ (.A(_3005_),
    .B(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__a21oi_1 _6795_ (.A1(_3010_),
    .A2(_3012_),
    .B1(_1629_),
    .Y(_0295_));
 sky130_fd_sc_hd__o31a_1 _6796_ (.A1(_1047_),
    .A2(_0908_),
    .A3(_1044_),
    .B1(_2181_),
    .X(_3013_));
 sky130_fd_sc_hd__inv_2 _6797_ (.A(_3005_),
    .Y(_3014_));
 sky130_fd_sc_hd__a21o_1 _6798_ (.A1(_2180_),
    .A2(_3014_),
    .B1(\as2650.psl[1] ),
    .X(_3015_));
 sky130_fd_sc_hd__o211a_1 _6799_ (.A1(_3005_),
    .A2(_3013_),
    .B1(_3015_),
    .C1(_2787_),
    .X(_0296_));
 sky130_fd_sc_hd__a211o_1 _6800_ (.A1(_0892_),
    .A2(_0895_),
    .B1(_0891_),
    .C1(\as2650.halted ),
    .X(_3016_));
 sky130_fd_sc_hd__nor2_1 _6801_ (.A(_3330_),
    .B(_0996_),
    .Y(_3017_));
 sky130_fd_sc_hd__o21ai_1 _6802_ (.A1(_3330_),
    .A2(_2706_),
    .B1(_3169_),
    .Y(_3018_));
 sky130_fd_sc_hd__or4_2 _6803_ (.A(_1010_),
    .B(_3016_),
    .C(_3017_),
    .D(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__nor2_1 _6804_ (.A(_0908_),
    .B(_0916_),
    .Y(_3020_));
 sky130_fd_sc_hd__o2bb2a_1 _6805_ (.A1_N(_3144_),
    .A2_N(_3020_),
    .B1(_3330_),
    .B2(_0545_),
    .X(_3021_));
 sky130_fd_sc_hd__a21oi_1 _6806_ (.A1(_1022_),
    .A2(_3330_),
    .B1(_3019_),
    .Y(_3022_));
 sky130_fd_sc_hd__or2_1 _6807_ (.A(io_out[26]),
    .B(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__o211a_1 _6808_ (.A1(_3019_),
    .A2(_3021_),
    .B1(_3023_),
    .C1(_1709_),
    .X(_0297_));
 sky130_fd_sc_hd__o21ai_1 _6809_ (.A1(_3000_),
    .A2(_3019_),
    .B1(\as2650.psu[4] ),
    .Y(_3024_));
 sky130_fd_sc_hd__or3_1 _6810_ (.A(_2191_),
    .B(_3020_),
    .C(_3019_),
    .X(_3025_));
 sky130_fd_sc_hd__a21oi_1 _6811_ (.A1(_3024_),
    .A2(_3025_),
    .B1(_1629_),
    .Y(_0298_));
 sky130_fd_sc_hd__o21ai_1 _6812_ (.A1(_3009_),
    .A2(_3019_),
    .B1(\as2650.psu[3] ),
    .Y(_3026_));
 sky130_fd_sc_hd__or3_1 _6813_ (.A(_2187_),
    .B(_3020_),
    .C(_3019_),
    .X(_3027_));
 sky130_fd_sc_hd__a21oi_1 _6814_ (.A1(_3026_),
    .A2(_3027_),
    .B1(_1629_),
    .Y(_0299_));
 sky130_fd_sc_hd__dfxtp_1 _6815_ (.CLK(clknet_leaf_7_clk),
    .D(_0000_),
    .Q(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6816_ (.CLK(clknet_leaf_7_clk),
    .D(_0001_),
    .Q(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6817_ (.CLK(clknet_leaf_7_clk),
    .D(_0002_),
    .Q(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6818_ (.CLK(clknet_leaf_7_clk),
    .D(_0003_),
    .Q(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6819_ (.CLK(clknet_leaf_7_clk),
    .D(_0004_),
    .Q(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6820_ (.CLK(clknet_leaf_7_clk),
    .D(_0005_),
    .Q(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6821_ (.CLK(clknet_leaf_7_clk),
    .D(_0006_),
    .Q(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6822_ (.CLK(clknet_leaf_8_clk),
    .D(_0007_),
    .Q(\as2650.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6823_ (.CLK(clknet_leaf_28_clk),
    .D(_0008_),
    .Q(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(clknet_leaf_28_clk),
    .D(_0009_),
    .Q(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(clknet_leaf_19_clk),
    .D(_0010_),
    .Q(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6826_ (.CLK(clknet_leaf_19_clk),
    .D(_0011_),
    .Q(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6827_ (.CLK(clknet_leaf_27_clk),
    .D(_0012_),
    .Q(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6828_ (.CLK(clknet_leaf_27_clk),
    .D(_0013_),
    .Q(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6829_ (.CLK(clknet_leaf_19_clk),
    .D(_0014_),
    .Q(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6830_ (.CLK(clknet_leaf_19_clk),
    .D(_0015_),
    .Q(\as2650.r123[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6831_ (.CLK(clknet_leaf_33_clk),
    .D(_0016_),
    .Q(\as2650.stack[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6832_ (.CLK(clknet_leaf_32_clk),
    .D(_0017_),
    .Q(\as2650.stack[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6833_ (.CLK(clknet_leaf_29_clk),
    .D(_0018_),
    .Q(\as2650.stack[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6834_ (.CLK(clknet_leaf_2_clk),
    .D(_0019_),
    .Q(\as2650.stack[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6835_ (.CLK(clknet_leaf_2_clk),
    .D(_0020_),
    .Q(\as2650.stack[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(clknet_leaf_31_clk),
    .D(_0021_),
    .Q(\as2650.stack[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(clknet_leaf_33_clk),
    .D(_0022_),
    .Q(\as2650.stack[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6838_ (.CLK(clknet_leaf_33_clk),
    .D(_0023_),
    .Q(\as2650.stack[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(clknet_leaf_32_clk),
    .D(_0024_),
    .Q(\as2650.stack[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6840_ (.CLK(clknet_leaf_26_clk),
    .D(_0025_),
    .Q(\as2650.stack[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6841_ (.CLK(clknet_leaf_24_clk),
    .D(_0026_),
    .Q(\as2650.stack[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6842_ (.CLK(clknet_leaf_31_clk),
    .D(_0027_),
    .Q(\as2650.stack[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6843_ (.CLK(clknet_leaf_25_clk),
    .D(_0028_),
    .Q(\as2650.stack[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(clknet_leaf_25_clk),
    .D(_0029_),
    .Q(\as2650.stack[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6845_ (.CLK(clknet_leaf_32_clk),
    .D(_0030_),
    .Q(\as2650.stack[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6846_ (.CLK(clknet_leaf_19_clk),
    .D(_0031_),
    .Q(\as2650.r123_2[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6847_ (.CLK(clknet_leaf_19_clk),
    .D(_0032_),
    .Q(\as2650.r123_2[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6848_ (.CLK(clknet_leaf_19_clk),
    .D(_0033_),
    .Q(\as2650.r123_2[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6849_ (.CLK(clknet_leaf_19_clk),
    .D(_0034_),
    .Q(\as2650.r123_2[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(clknet_leaf_19_clk),
    .D(_0035_),
    .Q(\as2650.r123_2[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6851_ (.CLK(clknet_leaf_19_clk),
    .D(_0036_),
    .Q(\as2650.r123_2[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(clknet_leaf_19_clk),
    .D(_0037_),
    .Q(\as2650.r123_2[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6853_ (.CLK(clknet_leaf_18_clk),
    .D(_0038_),
    .Q(\as2650.r123_2[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(clknet_leaf_28_clk),
    .D(_0039_),
    .Q(\as2650.psu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(clknet_leaf_32_clk),
    .D(_0040_),
    .Q(\as2650.stack[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6856_ (.CLK(clknet_leaf_25_clk),
    .D(_0041_),
    .Q(\as2650.stack[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(clknet_leaf_24_clk),
    .D(_0042_),
    .Q(\as2650.stack[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(clknet_leaf_31_clk),
    .D(_0043_),
    .Q(\as2650.stack[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(clknet_leaf_25_clk),
    .D(_0044_),
    .Q(\as2650.stack[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6860_ (.CLK(clknet_leaf_25_clk),
    .D(_0045_),
    .Q(\as2650.stack[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6861_ (.CLK(clknet_leaf_32_clk),
    .D(_0046_),
    .Q(\as2650.stack[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6862_ (.CLK(clknet_leaf_32_clk),
    .D(_0047_),
    .Q(\as2650.stack[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6863_ (.CLK(clknet_leaf_26_clk),
    .D(_0048_),
    .Q(\as2650.stack[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6864_ (.CLK(clknet_leaf_24_clk),
    .D(_0049_),
    .Q(\as2650.stack[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6865_ (.CLK(clknet_leaf_31_clk),
    .D(_0050_),
    .Q(\as2650.stack[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6866_ (.CLK(clknet_leaf_24_clk),
    .D(_0051_),
    .Q(\as2650.stack[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6867_ (.CLK(clknet_leaf_24_clk),
    .D(_0052_),
    .Q(\as2650.stack[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6868_ (.CLK(clknet_leaf_32_clk),
    .D(_0053_),
    .Q(\as2650.stack[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6869_ (.CLK(clknet_leaf_17_clk),
    .D(_0054_),
    .Q(\as2650.psl[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(clknet_leaf_17_clk),
    .D(_0055_),
    .Q(\as2650.psl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(clknet_leaf_31_clk),
    .D(_0056_),
    .Q(\as2650.stack[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(clknet_leaf_28_clk),
    .D(_0057_),
    .Q(\as2650.stack[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(clknet_leaf_28_clk),
    .D(_0058_),
    .Q(\as2650.stack[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6874_ (.CLK(clknet_leaf_29_clk),
    .D(_0059_),
    .Q(\as2650.stack[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(clknet_leaf_26_clk),
    .D(_0060_),
    .Q(\as2650.stack[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6876_ (.CLK(clknet_leaf_26_clk),
    .D(_0061_),
    .Q(\as2650.stack[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(clknet_leaf_31_clk),
    .D(_0062_),
    .Q(\as2650.stack[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6878_ (.CLK(clknet_leaf_20_clk),
    .D(_0063_),
    .Q(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6879_ (.CLK(clknet_leaf_17_clk),
    .D(_0064_),
    .Q(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6880_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0065_),
    .Q(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6881_ (.CLK(clknet_leaf_11_clk),
    .D(_0066_),
    .Q(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6882_ (.CLK(clknet_leaf_11_clk),
    .D(_0067_),
    .Q(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(clknet_leaf_11_clk),
    .D(_0068_),
    .Q(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6884_ (.CLK(clknet_leaf_31_clk),
    .D(_0069_),
    .Q(\as2650.stack[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(clknet_leaf_27_clk),
    .D(_0070_),
    .Q(\as2650.stack[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6886_ (.CLK(clknet_leaf_27_clk),
    .D(_0071_),
    .Q(\as2650.stack[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6887_ (.CLK(clknet_leaf_31_clk),
    .D(_0072_),
    .Q(\as2650.stack[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6888_ (.CLK(clknet_leaf_26_clk),
    .D(_0073_),
    .Q(\as2650.stack[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6889_ (.CLK(clknet_leaf_26_clk),
    .D(_0074_),
    .Q(\as2650.stack[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6890_ (.CLK(clknet_leaf_31_clk),
    .D(_0075_),
    .Q(\as2650.stack[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(clknet_leaf_19_clk),
    .D(_0076_),
    .Q(\as2650.r123_2[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6892_ (.CLK(clknet_leaf_20_clk),
    .D(_0077_),
    .Q(\as2650.r123_2[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(clknet_leaf_20_clk),
    .D(_0078_),
    .Q(\as2650.r123_2[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6894_ (.CLK(clknet_leaf_20_clk),
    .D(_0079_),
    .Q(\as2650.r123_2[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(clknet_leaf_20_clk),
    .D(_0080_),
    .Q(\as2650.r123_2[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0081_),
    .Q(\as2650.r123_2[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(clknet_leaf_20_clk),
    .D(_0082_),
    .Q(\as2650.r123_2[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(clknet_leaf_19_clk),
    .D(_0083_),
    .Q(\as2650.r123_2[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(clknet_leaf_32_clk),
    .D(_0084_),
    .Q(\as2650.stack[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(clknet_leaf_29_clk),
    .D(_0085_),
    .Q(\as2650.stack[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(clknet_leaf_27_clk),
    .D(_0086_),
    .Q(\as2650.stack[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_leaf_29_clk),
    .D(_0087_),
    .Q(\as2650.stack[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(clknet_leaf_26_clk),
    .D(_0088_),
    .Q(\as2650.stack[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(clknet_leaf_25_clk),
    .D(_0089_),
    .Q(\as2650.stack[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(clknet_leaf_32_clk),
    .D(_0090_),
    .Q(\as2650.stack[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(clknet_leaf_25_clk),
    .D(_0091_),
    .Q(\as2650.stack[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(clknet_leaf_26_clk),
    .D(_0092_),
    .Q(\as2650.stack[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(clknet_leaf_27_clk),
    .D(_0093_),
    .Q(\as2650.stack[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(clknet_leaf_31_clk),
    .D(_0094_),
    .Q(\as2650.stack[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(clknet_leaf_26_clk),
    .D(_0095_),
    .Q(\as2650.stack[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(clknet_leaf_26_clk),
    .D(_0096_),
    .Q(\as2650.stack[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6912_ (.CLK(clknet_leaf_31_clk),
    .D(_0097_),
    .Q(\as2650.stack[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6913_ (.CLK(clknet_leaf_0_clk),
    .D(_0098_),
    .Q(\as2650.r123_2[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6914_ (.CLK(clknet_leaf_36_clk),
    .D(_0099_),
    .Q(\as2650.r123_2[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(clknet_leaf_22_clk),
    .D(_0100_),
    .Q(\as2650.r123_2[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(clknet_leaf_1_clk),
    .D(_0101_),
    .Q(\as2650.r123_2[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6917_ (.CLK(clknet_leaf_22_clk),
    .D(_0102_),
    .Q(\as2650.r123_2[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6918_ (.CLK(clknet_leaf_23_clk),
    .D(_0103_),
    .Q(\as2650.r123_2[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6919_ (.CLK(clknet_leaf_36_clk),
    .D(_0104_),
    .Q(\as2650.r123_2[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(clknet_leaf_22_clk),
    .D(_0105_),
    .Q(\as2650.r123_2[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6921_ (.CLK(clknet_leaf_16_clk),
    .D(_0106_),
    .Q(\as2650.r123_2[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(clknet_leaf_15_clk),
    .D(_0107_),
    .Q(\as2650.r123_2[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(clknet_leaf_15_clk),
    .D(_0108_),
    .Q(\as2650.r123_2[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(clknet_leaf_15_clk),
    .D(_0109_),
    .Q(\as2650.r123_2[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(clknet_leaf_15_clk),
    .D(_0110_),
    .Q(\as2650.r123_2[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6926_ (.CLK(clknet_leaf_15_clk),
    .D(_0111_),
    .Q(\as2650.r123_2[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(clknet_leaf_17_clk),
    .D(_0112_),
    .Q(\as2650.r123_2[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(clknet_leaf_18_clk),
    .D(_0113_),
    .Q(\as2650.r123_2[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(clknet_leaf_33_clk),
    .D(_0114_),
    .Q(\as2650.stack[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(clknet_leaf_32_clk),
    .D(_0115_),
    .Q(\as2650.stack[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(clknet_leaf_29_clk),
    .D(_0116_),
    .Q(\as2650.stack[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(clknet_leaf_30_clk),
    .D(_0117_),
    .Q(\as2650.stack[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(clknet_leaf_29_clk),
    .D(_0118_),
    .Q(\as2650.stack[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(clknet_leaf_31_clk),
    .D(_0119_),
    .Q(\as2650.stack[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(clknet_leaf_33_clk),
    .D(_0120_),
    .Q(\as2650.stack[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(clknet_leaf_33_clk),
    .D(_0121_),
    .Q(\as2650.stack[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(clknet_leaf_35_clk),
    .D(_0122_),
    .Q(\as2650.stack[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(clknet_leaf_35_clk),
    .D(_0123_),
    .Q(\as2650.stack[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(clknet_leaf_29_clk),
    .D(_0124_),
    .Q(\as2650.stack[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(clknet_leaf_37_clk),
    .D(_0125_),
    .Q(\as2650.stack[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(clknet_leaf_2_clk),
    .D(_0126_),
    .Q(\as2650.stack[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(clknet_leaf_34_clk),
    .D(_0127_),
    .Q(\as2650.stack[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(clknet_leaf_34_clk),
    .D(_0128_),
    .Q(\as2650.stack[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(clknet_leaf_34_clk),
    .D(_0129_),
    .Q(\as2650.stack[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(clknet_leaf_36_clk),
    .D(_0130_),
    .Q(\as2650.stack[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(clknet_leaf_34_clk),
    .D(_0131_),
    .Q(\as2650.stack[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(clknet_leaf_2_clk),
    .D(_0132_),
    .Q(\as2650.stack[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(clknet_leaf_37_clk),
    .D(_0133_),
    .Q(\as2650.stack[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(clknet_leaf_37_clk),
    .D(_0134_),
    .Q(\as2650.stack[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(clknet_leaf_37_clk),
    .D(_0135_),
    .Q(\as2650.stack[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6951_ (.CLK(clknet_leaf_34_clk),
    .D(_0136_),
    .Q(\as2650.stack[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(clknet_leaf_34_clk),
    .D(_0137_),
    .Q(\as2650.stack[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6953_ (.CLK(clknet_leaf_22_clk),
    .D(_0138_),
    .Q(\as2650.r123[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(clknet_leaf_1_clk),
    .D(_0139_),
    .Q(\as2650.r123[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(clknet_leaf_23_clk),
    .D(_0140_),
    .Q(\as2650.r123[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6956_ (.CLK(clknet_leaf_22_clk),
    .D(_0141_),
    .Q(\as2650.r123[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6957_ (.CLK(clknet_leaf_22_clk),
    .D(_0142_),
    .Q(\as2650.r123[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6958_ (.CLK(clknet_leaf_0_clk),
    .D(_0143_),
    .Q(\as2650.r123[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6959_ (.CLK(clknet_leaf_22_clk),
    .D(_0144_),
    .Q(\as2650.r123[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6960_ (.CLK(clknet_leaf_36_clk),
    .D(_0145_),
    .Q(\as2650.r123[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6961_ (.CLK(clknet_leaf_35_clk),
    .D(_0146_),
    .Q(\as2650.stack[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6962_ (.CLK(clknet_leaf_35_clk),
    .D(_0147_),
    .Q(\as2650.stack[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(clknet_leaf_30_clk),
    .D(_0148_),
    .Q(\as2650.stack[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6964_ (.CLK(clknet_leaf_37_clk),
    .D(_0149_),
    .Q(\as2650.stack[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(clknet_leaf_37_clk),
    .D(_0150_),
    .Q(\as2650.stack[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(clknet_leaf_34_clk),
    .D(_0151_),
    .Q(\as2650.stack[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(clknet_leaf_34_clk),
    .D(_0152_),
    .Q(\as2650.stack[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(clknet_leaf_34_clk),
    .D(_0153_),
    .Q(\as2650.stack[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(clknet_leaf_24_clk),
    .D(_0154_),
    .Q(\lfsr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(clknet_leaf_24_clk),
    .D(_0155_),
    .Q(\lfsr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(clknet_leaf_26_clk),
    .D(_0156_),
    .Q(\lfsr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(clknet_leaf_26_clk),
    .D(_0157_),
    .Q(\lfsr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(clknet_leaf_26_clk),
    .D(_0158_),
    .Q(\lfsr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(clknet_leaf_27_clk),
    .D(_0159_),
    .Q(\as2650.sense ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_leaf_26_clk),
    .D(_0160_),
    .Q(\lfsr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_leaf_26_clk),
    .D(_0161_),
    .Q(\lfsr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_leaf_24_clk),
    .D(_0162_),
    .Q(\lfsr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_leaf_24_clk),
    .D(_0163_),
    .Q(\lfsr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_leaf_24_clk),
    .D(_0164_),
    .Q(\lfsr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(clknet_leaf_24_clk),
    .D(_0165_),
    .Q(\lfsr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_leaf_24_clk),
    .D(_0166_),
    .Q(\lfsr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_leaf_24_clk),
    .D(_0167_),
    .Q(\lfsr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_leaf_24_clk),
    .D(_0168_),
    .Q(\lfsr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_leaf_24_clk),
    .D(_0169_),
    .Q(\lfsr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_leaf_36_clk),
    .D(_0170_),
    .Q(\as2650.stack[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_leaf_36_clk),
    .D(_0171_),
    .Q(\as2650.stack[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_leaf_37_clk),
    .D(_0172_),
    .Q(\as2650.stack[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(clknet_leaf_37_clk),
    .D(_0173_),
    .Q(\as2650.stack[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_leaf_37_clk),
    .D(_0174_),
    .Q(\as2650.stack[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(clknet_leaf_37_clk),
    .D(_0175_),
    .Q(\as2650.stack[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(clknet_leaf_34_clk),
    .D(_0176_),
    .Q(\as2650.stack[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(clknet_leaf_34_clk),
    .D(_0177_),
    .Q(\as2650.stack[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _6993_ (.CLK(clknet_leaf_6_clk),
    .D(_0178_),
    .Q(io_out[23]));
 sky130_fd_sc_hd__dfxtp_2 _6994_ (.CLK(clknet_leaf_7_clk),
    .D(_0179_),
    .Q(io_out[25]));
 sky130_fd_sc_hd__dfxtp_2 _6995_ (.CLK(clknet_leaf_10_clk),
    .D(_0180_),
    .Q(io_out[24]));
 sky130_fd_sc_hd__dfxtp_4 _6996_ (.CLK(clknet_leaf_4_clk),
    .D(_0181_),
    .Q(io_out[8]));
 sky130_fd_sc_hd__dfxtp_4 _6997_ (.CLK(clknet_leaf_4_clk),
    .D(_0182_),
    .Q(io_out[9]));
 sky130_fd_sc_hd__dfxtp_4 _6998_ (.CLK(clknet_leaf_6_clk),
    .D(_0183_),
    .Q(io_out[10]));
 sky130_fd_sc_hd__dfxtp_4 _6999_ (.CLK(clknet_leaf_6_clk),
    .D(_0184_),
    .Q(io_out[11]));
 sky130_fd_sc_hd__dfxtp_4 _7000_ (.CLK(clknet_leaf_6_clk),
    .D(_0185_),
    .Q(io_out[12]));
 sky130_fd_sc_hd__dfxtp_4 _7001_ (.CLK(clknet_leaf_4_clk),
    .D(_0186_),
    .Q(io_out[13]));
 sky130_fd_sc_hd__dfxtp_4 _7002_ (.CLK(clknet_leaf_6_clk),
    .D(_0187_),
    .Q(io_out[14]));
 sky130_fd_sc_hd__dfxtp_4 _7003_ (.CLK(clknet_leaf_4_clk),
    .D(_0188_),
    .Q(io_out[15]));
 sky130_fd_sc_hd__dfxtp_4 _7004_ (.CLK(clknet_leaf_4_clk),
    .D(_0189_),
    .Q(io_out[16]));
 sky130_fd_sc_hd__dfxtp_4 _7005_ (.CLK(clknet_leaf_4_clk),
    .D(_0190_),
    .Q(io_out[17]));
 sky130_fd_sc_hd__dfxtp_4 _7006_ (.CLK(clknet_leaf_4_clk),
    .D(_0191_),
    .Q(io_out[18]));
 sky130_fd_sc_hd__dfxtp_4 _7007_ (.CLK(clknet_leaf_4_clk),
    .D(_0192_),
    .Q(io_out[19]));
 sky130_fd_sc_hd__dfxtp_4 _7008_ (.CLK(clknet_leaf_4_clk),
    .D(_0193_),
    .Q(io_out[20]));
 sky130_fd_sc_hd__dfxtp_4 _7009_ (.CLK(clknet_leaf_3_clk),
    .D(_0194_),
    .Q(io_out[21]));
 sky130_fd_sc_hd__dfxtp_4 _7010_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0195_),
    .Q(io_out[22]));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(clknet_leaf_13_clk),
    .D(_0196_),
    .Q(\as2650.idx_ctrl[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7012_ (.CLK(clknet_leaf_13_clk),
    .D(_0197_),
    .Q(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7013_ (.CLK(clknet_leaf_16_clk),
    .D(_0198_),
    .Q(\as2650.holding_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7014_ (.CLK(clknet_leaf_15_clk),
    .D(_0199_),
    .Q(\as2650.holding_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7015_ (.CLK(clknet_leaf_15_clk),
    .D(_0200_),
    .Q(\as2650.holding_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7016_ (.CLK(clknet_leaf_14_clk),
    .D(_0201_),
    .Q(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7017_ (.CLK(clknet_leaf_14_clk),
    .D(_0202_),
    .Q(\as2650.holding_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7018_ (.CLK(clknet_leaf_14_clk),
    .D(_0203_),
    .Q(\as2650.holding_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7019_ (.CLK(clknet_leaf_17_clk),
    .D(_0204_),
    .Q(\as2650.holding_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7020_ (.CLK(clknet_leaf_16_clk),
    .D(_0205_),
    .Q(\as2650.holding_reg[7] ));
 sky130_fd_sc_hd__dfxtp_4 _7021_ (.CLK(clknet_leaf_10_clk),
    .D(_0206_),
    .Q(\as2650.halted ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(clknet_leaf_8_clk),
    .D(_0207_),
    .Q(\as2650.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(clknet_leaf_8_clk),
    .D(_0208_),
    .Q(\as2650.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(clknet_leaf_8_clk),
    .D(_0209_),
    .Q(\as2650.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(clknet_leaf_8_clk),
    .D(_0210_),
    .Q(\as2650.cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(clknet_leaf_8_clk),
    .D(_0211_),
    .Q(\as2650.cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(clknet_leaf_9_clk),
    .D(_0212_),
    .Q(\as2650.cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(clknet_leaf_9_clk),
    .D(_0213_),
    .Q(\as2650.cycle[6] ));
 sky130_fd_sc_hd__dfxtp_4 _7029_ (.CLK(clknet_leaf_9_clk),
    .D(_0214_),
    .Q(\as2650.cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7030_ (.CLK(clknet_leaf_3_clk),
    .D(_0215_),
    .Q(\as2650.psu[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(clknet_leaf_3_clk),
    .D(_0216_),
    .Q(\as2650.pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7032_ (.CLK(clknet_leaf_3_clk),
    .D(_0217_),
    .Q(\as2650.pc[1] ));
 sky130_fd_sc_hd__dfxtp_4 _7033_ (.CLK(clknet_leaf_2_clk),
    .D(_0218_),
    .Q(\as2650.pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7034_ (.CLK(clknet_leaf_2_clk),
    .D(_0219_),
    .Q(\as2650.pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7035_ (.CLK(clknet_leaf_2_clk),
    .D(_0220_),
    .Q(\as2650.pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7036_ (.CLK(clknet_leaf_2_clk),
    .D(_0221_),
    .Q(\as2650.pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(clknet_leaf_1_clk),
    .D(_0222_),
    .Q(\as2650.pc[6] ));
 sky130_fd_sc_hd__dfxtp_4 _7038_ (.CLK(clknet_leaf_0_clk),
    .D(_0223_),
    .Q(\as2650.pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7039_ (.CLK(clknet_leaf_0_clk),
    .D(_0224_),
    .Q(\as2650.pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_leaf_0_clk),
    .D(_0225_),
    .Q(\as2650.pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _7041_ (.CLK(clknet_leaf_0_clk),
    .D(_0226_),
    .Q(\as2650.pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_leaf_1_clk),
    .D(_0227_),
    .Q(\as2650.pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(clknet_leaf_1_clk),
    .D(_0228_),
    .Q(\as2650.pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7044_ (.CLK(clknet_leaf_2_clk),
    .D(_0229_),
    .Q(\as2650.pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _7045_ (.CLK(clknet_leaf_3_clk),
    .D(_0230_),
    .Q(\as2650.pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(clknet_leaf_16_clk),
    .D(_0231_),
    .Q(\as2650.r0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7047_ (.CLK(clknet_leaf_27_clk),
    .D(_0232_),
    .Q(\as2650.r0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7048_ (.CLK(clknet_leaf_27_clk),
    .D(_0233_),
    .Q(\as2650.r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7049_ (.CLK(clknet_leaf_27_clk),
    .D(_0234_),
    .Q(\as2650.r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(clknet_leaf_27_clk),
    .D(_0235_),
    .Q(\as2650.r0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7051_ (.CLK(clknet_leaf_27_clk),
    .D(_0236_),
    .Q(\as2650.r0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7052_ (.CLK(clknet_leaf_27_clk),
    .D(_0237_),
    .Q(\as2650.r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(clknet_leaf_27_clk),
    .D(_0238_),
    .Q(\as2650.r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(clknet_leaf_33_clk),
    .D(_0239_),
    .Q(\as2650.stack[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(clknet_leaf_31_clk),
    .D(_0240_),
    .Q(\as2650.stack[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(clknet_leaf_29_clk),
    .D(_0241_),
    .Q(\as2650.stack[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(clknet_leaf_30_clk),
    .D(_0242_),
    .Q(\as2650.stack[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(clknet_leaf_29_clk),
    .D(_0243_),
    .Q(\as2650.stack[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7059_ (.CLK(clknet_leaf_31_clk),
    .D(_0244_),
    .Q(\as2650.stack[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(clknet_leaf_32_clk),
    .D(_0245_),
    .Q(\as2650.stack[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7061_ (.CLK(clknet_leaf_33_clk),
    .D(_0246_),
    .Q(\as2650.stack[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7062_ (.CLK(clknet_leaf_32_clk),
    .D(_0247_),
    .Q(\as2650.stack[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(clknet_leaf_32_clk),
    .D(_0248_),
    .Q(\as2650.stack[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7064_ (.CLK(clknet_leaf_29_clk),
    .D(_0249_),
    .Q(\as2650.stack[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7065_ (.CLK(clknet_leaf_30_clk),
    .D(_0250_),
    .Q(\as2650.stack[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7066_ (.CLK(clknet_leaf_29_clk),
    .D(_0251_),
    .Q(\as2650.stack[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7067_ (.CLK(clknet_leaf_31_clk),
    .D(_0252_),
    .Q(\as2650.stack[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7068_ (.CLK(clknet_leaf_32_clk),
    .D(_0253_),
    .Q(\as2650.stack[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7069_ (.CLK(clknet_leaf_31_clk),
    .D(_0254_),
    .Q(\as2650.stack[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(clknet_leaf_32_clk),
    .D(_0255_),
    .Q(\as2650.stack[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(clknet_leaf_26_clk),
    .D(_0256_),
    .Q(\as2650.stack[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7072_ (.CLK(clknet_leaf_24_clk),
    .D(_0257_),
    .Q(\as2650.stack[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(clknet_leaf_26_clk),
    .D(_0258_),
    .Q(\as2650.stack[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(clknet_leaf_24_clk),
    .D(_0259_),
    .Q(\as2650.stack[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(clknet_leaf_25_clk),
    .D(_0260_),
    .Q(\as2650.stack[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7076_ (.CLK(clknet_leaf_32_clk),
    .D(_0261_),
    .Q(\as2650.stack[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7077_ (.CLK(clknet_leaf_19_clk),
    .D(_0262_),
    .Q(\as2650.r123[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7078_ (.CLK(clknet_leaf_20_clk),
    .D(_0263_),
    .Q(\as2650.r123[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(clknet_leaf_20_clk),
    .D(_0264_),
    .Q(\as2650.r123[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(clknet_leaf_20_clk),
    .D(_0265_),
    .Q(\as2650.r123[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(clknet_leaf_20_clk),
    .D(_0266_),
    .Q(\as2650.r123[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(clknet_leaf_20_clk),
    .D(_0267_),
    .Q(\as2650.r123[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(clknet_leaf_19_clk),
    .D(_0268_),
    .Q(\as2650.r123[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7084_ (.CLK(clknet_leaf_18_clk),
    .D(_0269_),
    .Q(\as2650.r123[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(clknet_leaf_15_clk),
    .D(_0270_),
    .Q(\as2650.r123[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(clknet_leaf_15_clk),
    .D(_0271_),
    .Q(\as2650.r123[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(clknet_leaf_15_clk),
    .D(_0272_),
    .Q(\as2650.r123[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(clknet_leaf_15_clk),
    .D(_0273_),
    .Q(\as2650.r123[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(clknet_leaf_15_clk),
    .D(_0274_),
    .Q(\as2650.r123[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(clknet_leaf_15_clk),
    .D(_0275_),
    .Q(\as2650.r123[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(clknet_leaf_16_clk),
    .D(_0276_),
    .Q(\as2650.r123[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(clknet_leaf_18_clk),
    .D(_0277_),
    .Q(\as2650.r123[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _7093_ (.CLK(clknet_leaf_0_clk),
    .D(_0278_),
    .Q(io_out[0]));
 sky130_fd_sc_hd__dfxtp_2 _7094_ (.CLK(clknet_leaf_0_clk),
    .D(_0279_),
    .Q(io_out[1]));
 sky130_fd_sc_hd__dfxtp_2 _7095_ (.CLK(clknet_leaf_0_clk),
    .D(_0280_),
    .Q(io_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _7096_ (.CLK(clknet_leaf_0_clk),
    .D(_0281_),
    .Q(io_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _7097_ (.CLK(clknet_leaf_0_clk),
    .D(_0282_),
    .Q(io_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _7098_ (.CLK(clknet_leaf_0_clk),
    .D(_0283_),
    .Q(io_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _7099_ (.CLK(clknet_leaf_0_clk),
    .D(_0284_),
    .Q(io_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _7100_ (.CLK(clknet_leaf_0_clk),
    .D(_0285_),
    .Q(io_out[7]));
 sky130_fd_sc_hd__dfxtp_2 _7101_ (.CLK(clknet_leaf_10_clk),
    .D(_0286_),
    .Q(\as2650.ins_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(clknet_leaf_11_clk),
    .D(_0287_),
    .Q(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(clknet_leaf_17_clk),
    .D(_0288_),
    .Q(\as2650.psl[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7104_ (.CLK(clknet_leaf_17_clk),
    .D(_0289_),
    .Q(\as2650.carry ));
 sky130_fd_sc_hd__dfxtp_4 _7105_ (.CLK(clknet_leaf_29_clk),
    .D(_0290_),
    .Q(\as2650.psu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7106_ (.CLK(clknet_leaf_29_clk),
    .D(_0291_),
    .Q(\as2650.psu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7107_ (.CLK(clknet_leaf_29_clk),
    .D(_0292_),
    .Q(\as2650.psu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7108_ (.CLK(clknet_leaf_18_clk),
    .D(_0293_),
    .Q(\as2650.overflow ));
 sky130_fd_sc_hd__dfxtp_1 _7109_ (.CLK(clknet_leaf_20_clk),
    .D(_0294_),
    .Q(\as2650.psl[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7110_ (.CLK(clknet_leaf_18_clk),
    .D(_0295_),
    .Q(\as2650.psl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7111_ (.CLK(clknet_leaf_18_clk),
    .D(_0296_),
    .Q(\as2650.psl[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7112_ (.CLK(clknet_leaf_28_clk),
    .D(_0297_),
    .Q(io_out[26]));
 sky130_fd_sc_hd__dfxtp_1 _7113_ (.CLK(clknet_leaf_18_clk),
    .D(_0298_),
    .Q(\as2650.psu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7114_ (.CLK(clknet_leaf_18_clk),
    .D(_0299_),
    .Q(\as2650.psu[3] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(rst),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__D (.DIODE(_0063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A0 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A1 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A1 (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A1 (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A2 (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A1 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__C1 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A2 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A2 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A2 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A2 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B1 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B1 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A2 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A1 (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A1 (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A1 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A0 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A1 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A0 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A1 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A1 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__B2 (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__B1 (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B2 (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A2 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A2 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A0 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(_0345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B (.DIODE(_0345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A (.DIODE(_0345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B (.DIODE(_0345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A1 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A1 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A3 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__C (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__D (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__B (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A0 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__B2 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B2 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__B1 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A2 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A0 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A0 (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__B (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__B1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__C1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__B1_N (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A2 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__C (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A1 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__B (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A0 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A0 (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A2 (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B (.DIODE(_0406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__B (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__B (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B1 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__B (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__D (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A0 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A1 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A1 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__S (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__C1 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__C1 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__C1 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__C1 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A1 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__D (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A2_N (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__D (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__B (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A0 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A0 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A2 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A_N (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A0 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__B1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B2 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A2 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__C (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A0 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A1 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A1 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B1 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__B2 (.DIODE(_0488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A1 (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B1 (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B1 (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A1 (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A0 (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__C (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A2 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A2 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A0 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A0 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A2 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A2 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B2 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A1 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B2 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A0 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A3 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__C (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A0 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A0 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A2 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A0 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A2 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__C (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A0 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A2 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A1 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__B (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A2 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B1 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A0 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__B (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A0 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A0 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A0 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__C1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__C1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__B1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__C1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__B2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__B1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__C1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A1 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B1 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A2 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__C (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__C (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__C (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__C (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__C (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A1 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B1 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__C (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__D1 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__S (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A0 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A0 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A0 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A0 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A1_N (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A0 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A0 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A0 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A0 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A0 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A0 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A0 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A0 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A0 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A0 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A0 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1_N (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A0 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A0 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A1 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A0 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A0 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A0 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A0 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A0 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A0 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A0 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__B1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A2 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A1 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A2 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__C1 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__B (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A2 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__C1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A3 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__C (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__C (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__C (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__C (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A0 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A3 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__C1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__D (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__B2 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__C (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__C (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A0 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1_N (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B2 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B1 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__B (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__D (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__B1 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B1 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__D (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B1 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__C (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__C (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__C (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A0 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B2 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A0 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A1 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A2 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A2 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__D (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__C (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__B (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__B (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__B (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__C1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__C1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__S (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__S (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__C1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__D (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__B1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A2 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__B (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A1_N (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A1_N (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__B (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A1_N (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__B (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A1_N (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1 (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1_N (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__B (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A1_N (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1_N (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__B (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A0 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__B (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__B (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__B1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__B (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__S (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__S (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__S (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B2 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__C (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__C (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__C (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__B1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__C1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__D_N (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__C1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__C1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__B1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__C1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__C1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__C1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1_N (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__C1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__B1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__C (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__C1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__B (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__B2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__C1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__B (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__C (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__D (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__C_N (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__C_N (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__D (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A3 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__C (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__B (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__B (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__C1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B2 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__C (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A2 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A2 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__B (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__B (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__C1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A2 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B2 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__B (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A1 (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__B (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__C1 (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B2 (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(_0907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__B (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__S (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__S (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__S (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__B (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__C (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A3 (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__C (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A3 (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A1_N (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__C1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__C1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__C1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B2 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1_N (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__C1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__C1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__C1 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__C1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__C1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__D1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__B2 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__B2 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__C1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__C1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__C1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__C1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__C (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A3 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__C1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__C1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__C1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A2 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A2 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A3 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__C (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A1 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__B (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__D (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B1 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__C (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__B (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__B2 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__B2 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A1_N (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__D (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A_N (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A2_N (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A3 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__B (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B1 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__B1 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B1 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A1 (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A0 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__D1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B2 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__C1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__C1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__C1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__C1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A3 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A3 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A2 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A3 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A0 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A0 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B1 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B2 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__B1 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A2 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A1 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A2 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B1 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B1 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__C (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__B (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__B (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__S (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(_1080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__S (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__B1 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__B1 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B2 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__C (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B1 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B1 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B1 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__C1 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B2 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__B1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A2 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__C (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A3 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B2 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A2 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A2 (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A2 (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A2_N (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A2 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__C (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A2 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A2 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__C (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A2 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A2 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A2 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B1 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A2 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A2 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B1 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A2 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A2 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A2 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A2 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A0 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1_N (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__S (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A1 (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B1 (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__B1 (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__C (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B2 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__B1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__C1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__B1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__C1 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A0 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__B2 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__B1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__C (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B2 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__C1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__C1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__B (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__B2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A1 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A3 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__D (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__S (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__C (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1_N (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B2 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__C1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__B1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A3 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__C1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__C1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__B1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B2 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__B1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A2 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__D1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B2 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A1_N (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A3 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__C1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__C1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__C1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A3 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B1 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__C (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A2_N (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B2 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2_N (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__B (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__B1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__C1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B2 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B2 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__B2 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(_1721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A1 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1_N (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__B2 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A1 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A1_N (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__B1 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A2 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A3 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__B2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__B2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__C1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B1 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__B (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A1 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__B1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__C1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__B1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__C1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B2 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__C1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A2 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A2 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A1 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B1 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__S (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A2 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__S (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A1_N (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1_N (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A2 (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1 (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A2 (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B1 (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A (.DIODE(_1865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A1 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__C1 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B1 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__C1 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B2 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A1 (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B1 (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__C (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__C1 (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(_1882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A2 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__C1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__C1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__C1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__B2 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__C1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__C1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__B (.DIODE(_2018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__C_N (.DIODE(_2018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A1 (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A3 (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A2 (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B2 (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__C1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__B1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__C1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1_N (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__C1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__C1 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A2 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__B1 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B1 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__S (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A0 (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A2 (.DIODE(_2184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A0 (.DIODE(_2184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__C1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__C1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__C1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__C1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__C1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A2 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__B1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A2 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A2 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A1_N (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B2 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A2 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B1 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__B1 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A2 (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A (.DIODE(_2270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A1 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A1 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A1 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__B2 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__D1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__C1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__C1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__C1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__S (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A2 (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A2 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B1 (.DIODE(_2391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__B1 (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A2 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A2 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A0 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__B1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__C1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__B (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A2_N (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__C1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__B1 (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B1 (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A2 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__B1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__C1 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__B1 (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__B1 (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A2 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A2 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__C1 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__C1 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__C1 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A2 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__S (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__B (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__B (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__B (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__S (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__S (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__S (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A (.DIODE(_2889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A (.DIODE(_2892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__B1 (.DIODE(_2901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__B1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A2 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B (.DIODE(_2997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A0 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__B1 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A1 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A1 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__B1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B2 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A0 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__B2 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B2 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__C (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A2 (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__B (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A (.DIODE(_3037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__B (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__B (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A (.DIODE(_3039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A1 (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A1 (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A2_N (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__C (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B1 (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A2 (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__B2 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__C1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B2 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__B (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__B (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__C (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__B (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__B1 (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B (.DIODE(_3056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B2 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__C_N (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__C1 (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__C1 (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_3061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__B (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A0 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__B (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A_N (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A_N (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__C (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__B (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__B2 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B2 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B2 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B2 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__C (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__C (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A1 (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__C (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__B1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__C1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__C (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A3 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__B (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A2 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A3 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A1 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__S (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__S (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__S (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A3 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A1 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A1 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__B (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A3 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__S (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1_N (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__S (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__C1 (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B1 (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_3091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A2 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A1 (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__B (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A2 (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__B1 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__C1 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B2 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B1 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B1 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A3 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A1 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__C (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__B2 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B2 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B2 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__B (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__C1 (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B (.DIODE(_3107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__C (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__B1 (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__B1 (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__B (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__C1 (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A1 (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__C (.DIODE(_3121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B2 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A0 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A0 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A0 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A0 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A0 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A0 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A0 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A0 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A0 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A1 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A0 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A1 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A1 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A0 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B1 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B2 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A0 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A0 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A0 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__C (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A0 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A0 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(_3139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B2 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__D (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A0 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B1 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B1 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A1 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1_N (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A1 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B2 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B2 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A1 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A0 (.DIODE(_3144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A1 (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A (.DIODE(_3146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__S (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__S (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__B (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B2 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__S (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__B (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A2 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A2 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A2 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B1 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A2 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A2 (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(_3149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__S (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__B2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A0 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A0 (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A1 (.DIODE(_3151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__B1 (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__C1 (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__C1 (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A1 (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A2 (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A1 (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B2 (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B1 (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__B (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A (.DIODE(_3160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S1 (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__S (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B1 (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A1 (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__S1 (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__S1 (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__S (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A (.DIODE(_3163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__D (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A3 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A2 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A2 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A2 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A2 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__S (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__S (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__B (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__C (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__C (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__C (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__B (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__B (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__S (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__S (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__B (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__S0 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__S0 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A1 (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__B (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__C (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__C (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__B (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__B (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B1 (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A1 (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__S (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__S (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__S (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A1 (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__S (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__S (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A (.DIODE(_3202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A2 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A2 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__B (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A2 (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B1 (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B2 (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B1 (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__C (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__D (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A3 (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A2 (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__B (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__B (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__C (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__C (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A1 (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A1 (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A1 (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B2 (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__B (.DIODE(_3220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__B (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A1 (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__C1 (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A1 (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B2 (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__C (.DIODE(_3221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A1 (.DIODE(_3226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A1 (.DIODE(_3226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A2 (.DIODE(_3226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B2 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B2 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A2 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A2 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A3 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__C (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B1 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A1 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__C (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A2 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A0 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__S (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A1 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A1 (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A2 (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__C (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A2 (.DIODE(_3250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__C1 (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A2 (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A1 (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A (.DIODE(_3252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__B1 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__S (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__S (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__S (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__S (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__C (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__D (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A0 (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A3 (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A2 (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A2 (.DIODE(_3260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__C1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A0 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__C (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__B (.DIODE(_3265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__B (.DIODE(_3265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B1 (.DIODE(_3265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A1 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A3 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A2 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__B1 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__B (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A2 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A0 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A2 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A1 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A2 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A2 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__B2 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A2 (.DIODE(_3280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A2 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A1 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A0 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B (.DIODE(_3287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__B1 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__S (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__S (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__B (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__B1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B1 (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(_3318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__C (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A2 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__C1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__C1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__C1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__C1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__C1 (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A1 (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A0 (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A1 (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A1 (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A (.DIODE(_3323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__S (.DIODE(_3326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A (.DIODE(_3326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(_3326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(_3329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B2 (.DIODE(_3329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(_3329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A2 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__B1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A2 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A_N (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B2 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A1 (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(_3334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__C (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B (.DIODE(_3335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__B2 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B2 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__C1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A1 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A1 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__S0 (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(_3339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A0 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__S1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__B1 (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A2 (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__B1 (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A2 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A2 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B1 (.DIODE(_3346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A2 (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B1 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A2 (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(_3351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__B (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B1 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__B1 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__B1 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A2 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A1 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B1 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A2 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__C (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A3 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A2 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__D_N (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__B (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__C (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A1 (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A0 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B2 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A0 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__B (.DIODE(_3392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B (.DIODE(_3392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B1 (.DIODE(_3392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A1 (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A3 (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__C (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A (.DIODE(_3395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A1 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__B (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A0 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A2 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__B2 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B1 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A0 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A2 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A2 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A1 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B2 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A1 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A1 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A1 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A0 (.DIODE(_3398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B2 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B2 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A2 (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A1 (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__B (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B2 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B2 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1_N (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__C (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__B1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__B1_N (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__D1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B2 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__B2 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__B2 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B2 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A_N (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A0 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__B (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A_N (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A1 (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A1 (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__C1 (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__C1 (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B1 (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B1 (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__B (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A_N (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A (.DIODE(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__D1 (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B (.DIODE(\as2650.pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A (.DIODE(\as2650.pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(\as2650.pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__B2 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__B1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A0 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A0 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__B (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A (.DIODE(\as2650.pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A0 (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B1 (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B1 (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A (.DIODE(\as2650.pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(\as2650.pc[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(\as2650.pc[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A1 (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B1 (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A0 (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A (.DIODE(\as2650.pc[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__B1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B2 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__B_N (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A1 (.DIODE(\as2650.psl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A0 (.DIODE(\as2650.psl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__B2 (.DIODE(\as2650.psl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B2 (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B2 (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__B2 (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A1 (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1 (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A1 (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(\as2650.r0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A (.DIODE(\as2650.r0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A (.DIODE(\as2650.r0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A (.DIODE(\as2650.r0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(\as2650.r0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A1 (.DIODE(\as2650.r0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(\as2650.r0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A (.DIODE(\as2650.r0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(\as2650.r0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A1 (.DIODE(\as2650.r0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A0 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A0 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A0 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A1 (.DIODE(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A0 (.DIODE(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A1 (.DIODE(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A0 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A0 (.DIODE(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A1 (.DIODE(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A1 (.DIODE(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A0 (.DIODE(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A1 (.DIODE(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B2 (.DIODE(\as2650.sense ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B (.DIODE(\as2650.sense ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A1 (.DIODE(io_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A1 (.DIODE(io_out[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(io_out[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(io_out[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A1 (.DIODE(io_out[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B1 (.DIODE(io_out[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(io_out[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A (.DIODE(io_out[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A1 (.DIODE(io_out[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A (.DIODE(io_out[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A (.DIODE(io_out[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A0 (.DIODE(io_out[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__B (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B2 (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(io_out[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(io_out[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A (.DIODE(io_out[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A1 (.DIODE(io_out[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B1 (.DIODE(io_out[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A (.DIODE(io_out[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(io_out[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A0 (.DIODE(io_out[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A1 (.DIODE(io_out[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A (.DIODE(io_out[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(io_out[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(io_out[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(io_out[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(io_out[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(io_out[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__B1 (.DIODE(io_out[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A (.DIODE(io_out[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A (.DIODE(io_out[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(io_out[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A1 (.DIODE(io_out[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A (.DIODE(io_out[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A (.DIODE(io_out[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A1 (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A (.DIODE(io_out[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(io_out[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(io_out[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B1 (.DIODE(io_out[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(io_out[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A0 (.DIODE(io_out[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A1 (.DIODE(io_out[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A (.DIODE(io_out[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(io_out[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A0 (.DIODE(io_out[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(io_out[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A0 (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A1 (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A1 (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(io_out[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1 (.DIODE(io_out[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(io_out[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(io_out[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B1_N (.DIODE(io_out[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(io_out[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A (.DIODE(io_out[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A1 (.DIODE(io_out[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B2 (.DIODE(io_out[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A1 (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A1 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A1 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A2 (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__C (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A0 (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(io_out[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A1 (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A0 (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A0 (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A (.DIODE(io_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_895 ();
endmodule

