magic
tech sky130B
magscale 1 2
timestamp 1674823762
<< viali >>
rect 1869 15521 1903 15555
rect 2329 15521 2363 15555
rect 8585 15521 8619 15555
rect 9505 15521 9539 15555
rect 2605 15453 2639 15487
rect 4261 15453 4295 15487
rect 4813 15453 4847 15487
rect 5365 15453 5399 15487
rect 6837 15453 6871 15487
rect 8309 15453 8343 15487
rect 9781 15453 9815 15487
rect 5549 15385 5583 15419
rect 4077 15317 4111 15351
rect 6929 15317 6963 15351
rect 4629 15113 4663 15147
rect 5641 15113 5675 15147
rect 6653 15113 6687 15147
rect 8677 15113 8711 15147
rect 1593 14977 1627 15011
rect 4169 14977 4203 15011
rect 5733 14977 5767 15011
rect 5825 14977 5859 15011
rect 10333 14977 10367 15011
rect 1869 14909 1903 14943
rect 5457 14909 5491 14943
rect 10057 14909 10091 14943
rect 3985 14773 4019 14807
rect 5549 14773 5583 14807
rect 1593 14569 1627 14603
rect 4077 14569 4111 14603
rect 9689 14569 9723 14603
rect 10333 14569 10367 14603
rect 7113 14433 7147 14467
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 3985 14365 4019 14399
rect 4261 14365 4295 14399
rect 4445 14365 4479 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 6101 14365 6135 14399
rect 7225 14365 7259 14399
rect 7757 14365 7791 14399
rect 7941 14365 7975 14399
rect 4721 14297 4755 14331
rect 5917 14297 5951 14331
rect 6837 14297 6871 14331
rect 7021 14297 7055 14331
rect 7113 14297 7147 14331
rect 3249 14229 3283 14263
rect 4353 14229 4387 14263
rect 5549 14229 5583 14263
rect 7849 14229 7883 14263
rect 5549 14025 5583 14059
rect 7205 14025 7239 14059
rect 8217 14025 8251 14059
rect 3893 13957 3927 13991
rect 4629 13957 4663 13991
rect 7665 13957 7699 13991
rect 2145 13889 2179 13923
rect 2329 13889 2363 13923
rect 2881 13889 2915 13923
rect 3709 13889 3743 13923
rect 3801 13889 3835 13923
rect 4077 13889 4111 13923
rect 4537 13889 4571 13923
rect 4721 13889 4755 13923
rect 5365 13889 5399 13923
rect 5641 13889 5675 13923
rect 6561 13889 6595 13923
rect 6654 13889 6688 13923
rect 6837 13889 6871 13923
rect 6929 13889 6963 13923
rect 7067 13889 7101 13923
rect 7849 13889 7883 13923
rect 7941 13889 7975 13923
rect 8033 13889 8067 13923
rect 2237 13821 2271 13855
rect 5181 13821 5215 13855
rect 2881 13753 2915 13787
rect 3525 13685 3559 13719
rect 8033 13481 8067 13515
rect 6101 13345 6135 13379
rect 6285 13345 6319 13379
rect 7297 13345 7331 13379
rect 8125 13345 8159 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 2973 13277 3007 13311
rect 3249 13277 3283 13311
rect 4537 13277 4571 13311
rect 4813 13277 4847 13311
rect 4905 13277 4939 13311
rect 6561 13277 6595 13311
rect 7205 13277 7239 13311
rect 8033 13277 8067 13311
rect 3065 13209 3099 13243
rect 4721 13209 4755 13243
rect 2513 13141 2547 13175
rect 3433 13141 3467 13175
rect 5089 13141 5123 13175
rect 6469 13141 6503 13175
rect 7573 13141 7607 13175
rect 8401 13141 8435 13175
rect 3617 12869 3651 12903
rect 5549 12869 5583 12903
rect 6561 12869 6595 12903
rect 6745 12869 6779 12903
rect 2881 12801 2915 12835
rect 3893 12801 3927 12835
rect 4629 12801 4663 12835
rect 4813 12801 4847 12835
rect 5273 12801 5307 12835
rect 5365 12801 5399 12835
rect 6837 12801 6871 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 3157 12733 3191 12767
rect 3709 12733 3743 12767
rect 3065 12665 3099 12699
rect 2697 12597 2731 12631
rect 3617 12597 3651 12631
rect 4077 12597 4111 12631
rect 4721 12597 4755 12631
rect 5273 12597 5307 12631
rect 6653 12597 6687 12631
rect 7389 12597 7423 12631
rect 8033 12597 8067 12631
rect 7849 12325 7883 12359
rect 8585 12325 8619 12359
rect 3157 12189 3191 12223
rect 4629 12189 4663 12223
rect 4813 12189 4847 12223
rect 7573 12189 7607 12223
rect 7665 12189 7699 12223
rect 7849 12189 7883 12223
rect 8309 12189 8343 12223
rect 8401 12189 8435 12223
rect 8585 12121 8619 12155
rect 3065 12053 3099 12087
rect 4629 12053 4663 12087
rect 4169 11849 4203 11883
rect 6837 11849 6871 11883
rect 5181 11781 5215 11815
rect 4077 11713 4111 11747
rect 4353 11713 4387 11747
rect 4997 11713 5031 11747
rect 6745 11713 6779 11747
rect 7021 11713 7055 11747
rect 4353 11509 4387 11543
rect 4813 11509 4847 11543
rect 7021 11509 7055 11543
rect 6745 11305 6779 11339
rect 4445 11237 4479 11271
rect 4169 11169 4203 11203
rect 5273 11169 5307 11203
rect 5457 11169 5491 11203
rect 6101 11169 6135 11203
rect 7113 11169 7147 11203
rect 4445 11101 4479 11135
rect 4537 11101 4571 11135
rect 5181 11101 5215 11135
rect 5365 11101 5399 11135
rect 6009 11101 6043 11135
rect 6193 11101 6227 11135
rect 7021 11101 7055 11135
rect 7665 11101 7699 11135
rect 7849 11101 7883 11135
rect 4353 10965 4387 10999
rect 4997 10965 5031 10999
rect 7757 10965 7791 10999
rect 4185 10761 4219 10795
rect 6929 10761 6963 10795
rect 3985 10693 4019 10727
rect 5089 10693 5123 10727
rect 5181 10693 5215 10727
rect 4997 10625 5031 10659
rect 5365 10625 5399 10659
rect 6745 10625 6779 10659
rect 7021 10625 7055 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 7757 10625 7791 10659
rect 8401 10625 8435 10659
rect 8493 10557 8527 10591
rect 4169 10421 4203 10455
rect 4353 10421 4387 10455
rect 4813 10421 4847 10455
rect 6561 10421 6595 10455
rect 7941 10421 7975 10455
rect 8401 10421 8435 10455
rect 8769 10421 8803 10455
rect 5089 10217 5123 10251
rect 6837 10217 6871 10251
rect 7481 10217 7515 10251
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 7481 10013 7515 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8217 10013 8251 10047
rect 4905 9945 4939 9979
rect 5105 9945 5139 9979
rect 6101 9945 6135 9979
rect 6653 9945 6687 9979
rect 4261 9877 4295 9911
rect 5273 9877 5307 9911
rect 5733 9877 5767 9911
rect 6853 9877 6887 9911
rect 7021 9877 7055 9911
rect 8309 9877 8343 9911
rect 4813 9673 4847 9707
rect 6653 9673 6687 9707
rect 6009 9605 6043 9639
rect 7941 9605 7975 9639
rect 8861 9605 8895 9639
rect 4721 9537 4755 9571
rect 4997 9537 5031 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7849 9537 7883 9571
rect 8125 9537 8159 9571
rect 8769 9537 8803 9571
rect 9045 9537 9079 9571
rect 5733 9401 5767 9435
rect 7021 9401 7055 9435
rect 4997 9333 5031 9367
rect 5549 9333 5583 9367
rect 8309 9333 8343 9367
rect 9229 9333 9263 9367
rect 5733 8993 5767 9027
rect 6193 8993 6227 9027
rect 7481 8993 7515 9027
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 5825 8925 5859 8959
rect 7573 8925 7607 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 8493 8857 8527 8891
rect 5089 8789 5123 8823
rect 7941 8789 7975 8823
rect 8401 8449 8435 8483
rect 8493 8381 8527 8415
rect 8769 8313 8803 8347
rect 10057 3009 10091 3043
rect 10241 2805 10275 2839
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 4261 2397 4295 2431
rect 5273 2397 5307 2431
rect 6745 2397 6779 2431
rect 8217 2397 8251 2431
rect 9689 2397 9723 2431
rect 1685 2261 1719 2295
rect 2421 2261 2455 2295
rect 4077 2261 4111 2295
rect 5457 2261 5491 2295
rect 6929 2261 6963 2295
rect 8401 2261 8435 2295
rect 9873 2261 9907 2295
<< metal1 >>
rect 1104 15802 10856 15824
rect 1104 15750 2169 15802
rect 2221 15750 2233 15802
rect 2285 15750 2297 15802
rect 2349 15750 2361 15802
rect 2413 15750 2425 15802
rect 2477 15750 4607 15802
rect 4659 15750 4671 15802
rect 4723 15750 4735 15802
rect 4787 15750 4799 15802
rect 4851 15750 4863 15802
rect 4915 15750 7045 15802
rect 7097 15750 7109 15802
rect 7161 15750 7173 15802
rect 7225 15750 7237 15802
rect 7289 15750 7301 15802
rect 7353 15750 9483 15802
rect 9535 15750 9547 15802
rect 9599 15750 9611 15802
rect 9663 15750 9675 15802
rect 9727 15750 9739 15802
rect 9791 15750 10856 15802
rect 1104 15728 10856 15750
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 2317 15555 2375 15561
rect 2317 15552 2329 15555
rect 1903 15524 2329 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 2317 15521 2329 15524
rect 2363 15552 2375 15555
rect 2498 15552 2504 15564
rect 2363 15524 2504 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8168 15524 8585 15552
rect 8168 15512 8174 15524
rect 8573 15521 8585 15524
rect 8619 15552 8631 15555
rect 8662 15552 8668 15564
rect 8619 15524 8668 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9456 15524 9505 15552
rect 9456 15512 9462 15524
rect 9493 15521 9505 15524
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2593 15487 2651 15493
rect 2593 15484 2605 15487
rect 2096 15456 2605 15484
rect 2096 15444 2102 15456
rect 2593 15453 2605 15456
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 5350 15484 5356 15496
rect 4847 15456 5356 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6696 15456 6837 15484
rect 6696 15444 6702 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 8297 15487 8355 15493
rect 8297 15484 8309 15487
rect 6825 15447 6883 15453
rect 6932 15456 8309 15484
rect 5537 15419 5595 15425
rect 5537 15385 5549 15419
rect 5583 15416 5595 15419
rect 5718 15416 5724 15428
rect 5583 15388 5724 15416
rect 5583 15385 5595 15388
rect 5537 15379 5595 15385
rect 5718 15376 5724 15388
rect 5776 15376 5782 15428
rect 6178 15376 6184 15428
rect 6236 15416 6242 15428
rect 6932 15416 6960 15456
rect 8297 15453 8309 15456
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 6236 15388 6960 15416
rect 6236 15376 6242 15388
rect 7650 15376 7656 15428
rect 7708 15416 7714 15428
rect 9784 15416 9812 15447
rect 7708 15388 9812 15416
rect 7708 15376 7714 15388
rect 4062 15348 4068 15360
rect 4023 15320 4068 15348
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 1104 15258 11016 15280
rect 1104 15206 3388 15258
rect 3440 15206 3452 15258
rect 3504 15206 3516 15258
rect 3568 15206 3580 15258
rect 3632 15206 3644 15258
rect 3696 15206 5826 15258
rect 5878 15206 5890 15258
rect 5942 15206 5954 15258
rect 6006 15206 6018 15258
rect 6070 15206 6082 15258
rect 6134 15206 8264 15258
rect 8316 15206 8328 15258
rect 8380 15206 8392 15258
rect 8444 15206 8456 15258
rect 8508 15206 8520 15258
rect 8572 15206 10702 15258
rect 10754 15206 10766 15258
rect 10818 15206 10830 15258
rect 10882 15206 10894 15258
rect 10946 15206 10958 15258
rect 11010 15206 11016 15258
rect 1104 15184 11016 15206
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4212 15116 4629 15144
rect 4212 15104 4218 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 4617 15107 4675 15113
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 6178 15144 6184 15156
rect 5675 15116 6184 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 6638 15144 6644 15156
rect 6599 15116 6644 15144
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 1026 14968 1032 15020
rect 1084 15008 1090 15020
rect 1578 15008 1584 15020
rect 1084 14980 1584 15008
rect 1084 14968 1090 14980
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 1854 14940 1860 14952
rect 1815 14912 1860 14940
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 4172 14940 4200 14971
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 5592 14980 5733 15008
rect 5592 14968 5598 14980
rect 5721 14977 5733 14980
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 10318 15008 10324 15020
rect 5868 14980 5913 15008
rect 10231 14980 10324 15008
rect 5868 14968 5874 14980
rect 10318 14968 10324 14980
rect 10376 15008 10382 15020
rect 11054 15008 11060 15020
rect 10376 14980 11060 15008
rect 10376 14968 10382 14980
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 4338 14940 4344 14952
rect 4172 14912 4344 14940
rect 4338 14900 4344 14912
rect 4396 14940 4402 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 4396 14912 5457 14940
rect 4396 14900 4402 14912
rect 5445 14909 5457 14912
rect 5491 14940 5503 14943
rect 6914 14940 6920 14952
rect 5491 14912 6920 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 8168 14912 10057 14940
rect 8168 14900 8174 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3936 14776 3985 14804
rect 3936 14764 3942 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 5626 14804 5632 14816
rect 5583 14776 5632 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 1104 14714 10856 14736
rect 1104 14662 2169 14714
rect 2221 14662 2233 14714
rect 2285 14662 2297 14714
rect 2349 14662 2361 14714
rect 2413 14662 2425 14714
rect 2477 14662 4607 14714
rect 4659 14662 4671 14714
rect 4723 14662 4735 14714
rect 4787 14662 4799 14714
rect 4851 14662 4863 14714
rect 4915 14662 7045 14714
rect 7097 14662 7109 14714
rect 7161 14662 7173 14714
rect 7225 14662 7237 14714
rect 7289 14662 7301 14714
rect 7353 14662 9483 14714
rect 9535 14662 9547 14714
rect 9599 14662 9611 14714
rect 9663 14662 9675 14714
rect 9727 14662 9739 14714
rect 9791 14662 10856 14714
rect 1104 14640 10856 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 4062 14600 4068 14612
rect 3975 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14600 4126 14612
rect 5718 14600 5724 14612
rect 4120 14572 5724 14600
rect 4120 14560 4126 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 9398 14560 9404 14612
rect 9456 14600 9462 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9456 14572 9689 14600
rect 9456 14560 9462 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 10318 14600 10324 14612
rect 10279 14572 10324 14600
rect 9677 14563 9735 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 4080 14464 4108 14560
rect 7650 14532 7656 14544
rect 6840 14504 7656 14532
rect 4522 14464 4528 14476
rect 3108 14436 4108 14464
rect 4264 14436 4528 14464
rect 3108 14424 3114 14436
rect 3142 14356 3148 14408
rect 3200 14396 3206 14408
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 3200 14368 3249 14396
rect 3200 14356 3206 14368
rect 3237 14365 3249 14368
rect 3283 14396 3295 14399
rect 3326 14396 3332 14408
rect 3283 14368 3332 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 3436 14405 3464 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3421 14359 3479 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4264 14405 4292 14436
rect 4522 14424 4528 14436
rect 4580 14464 4586 14476
rect 6178 14464 6184 14476
rect 4580 14436 6184 14464
rect 4580 14424 4586 14436
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4080 14368 4261 14396
rect 2314 14288 2320 14340
rect 2372 14328 2378 14340
rect 3786 14328 3792 14340
rect 2372 14300 3792 14328
rect 2372 14288 2378 14300
rect 3786 14288 3792 14300
rect 3844 14328 3850 14340
rect 4080 14328 4108 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4430 14396 4436 14408
rect 4391 14368 4436 14396
rect 4249 14359 4307 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 5718 14396 5724 14408
rect 5679 14368 5724 14396
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 5828 14405 5856 14436
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6730 14396 6736 14408
rect 6135 14368 6736 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 3844 14300 4108 14328
rect 3844 14288 3850 14300
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4709 14331 4767 14337
rect 4709 14328 4721 14331
rect 4212 14300 4721 14328
rect 4212 14288 4218 14300
rect 4709 14297 4721 14300
rect 4755 14297 4767 14331
rect 4709 14291 4767 14297
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 6840 14337 6868 14504
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 7147 14436 7788 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 7760 14408 7788 14436
rect 7213 14399 7271 14405
rect 7213 14365 7225 14399
rect 7259 14396 7271 14399
rect 7742 14396 7748 14408
rect 7259 14368 7328 14396
rect 7703 14368 7748 14396
rect 7259 14365 7271 14368
rect 7213 14359 7271 14365
rect 5905 14331 5963 14337
rect 5905 14328 5917 14331
rect 4856 14300 5917 14328
rect 4856 14288 4862 14300
rect 5905 14297 5917 14300
rect 5951 14297 5963 14331
rect 5905 14291 5963 14297
rect 6825 14331 6883 14337
rect 6825 14297 6837 14331
rect 6871 14297 6883 14331
rect 6825 14291 6883 14297
rect 7009 14331 7067 14337
rect 7009 14297 7021 14331
rect 7055 14297 7067 14331
rect 7009 14291 7067 14297
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 3016 14232 3249 14260
rect 3016 14220 3022 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 3237 14223 3295 14229
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 4338 14260 4344 14272
rect 3384 14232 4344 14260
rect 3384 14220 3390 14232
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 5920 14260 5948 14291
rect 7024 14260 7052 14291
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 7300 14328 7328 14368
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 7926 14396 7932 14408
rect 7887 14368 7932 14396
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8110 14328 8116 14340
rect 7156 14300 7201 14328
rect 7300 14300 8116 14328
rect 7156 14288 7162 14300
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 7190 14260 7196 14272
rect 5868 14232 7196 14260
rect 5868 14220 5874 14232
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7834 14260 7840 14272
rect 7795 14232 7840 14260
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 1104 14170 11016 14192
rect 1104 14118 3388 14170
rect 3440 14118 3452 14170
rect 3504 14118 3516 14170
rect 3568 14118 3580 14170
rect 3632 14118 3644 14170
rect 3696 14118 5826 14170
rect 5878 14118 5890 14170
rect 5942 14118 5954 14170
rect 6006 14118 6018 14170
rect 6070 14118 6082 14170
rect 6134 14118 8264 14170
rect 8316 14118 8328 14170
rect 8380 14118 8392 14170
rect 8444 14118 8456 14170
rect 8508 14118 8520 14170
rect 8572 14118 10702 14170
rect 10754 14118 10766 14170
rect 10818 14118 10830 14170
rect 10882 14118 10894 14170
rect 10946 14118 10958 14170
rect 11010 14118 11016 14170
rect 1104 14096 11016 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 4430 14056 4436 14068
rect 2096 14028 4436 14056
rect 2096 14016 2102 14028
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 3896 13997 3924 14028
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5534 14056 5540 14068
rect 5495 14028 5540 14056
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 6822 14016 6828 14068
rect 6880 14016 6886 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6972 14028 7205 14056
rect 6972 14016 6978 14028
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 7984 14028 8217 14056
rect 7984 14016 7990 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 3881 13991 3939 13997
rect 1912 13960 3832 13988
rect 1912 13948 1918 13960
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 2096 13892 2145 13920
rect 2096 13880 2102 13892
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2133 13883 2191 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 3694 13920 3700 13932
rect 3655 13892 3700 13920
rect 2869 13883 2927 13889
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2774 13852 2780 13864
rect 2271 13824 2780 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 2884 13852 2912 13883
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 3804 13929 3832 13960
rect 3881 13957 3893 13991
rect 3927 13957 3939 13991
rect 3881 13951 3939 13957
rect 4617 13991 4675 13997
rect 4617 13957 4629 13991
rect 4663 13988 4675 13991
rect 5552 13988 5580 14016
rect 6840 13988 6868 14016
rect 7650 13988 7656 14000
rect 4663 13960 5488 13988
rect 5552 13960 6684 13988
rect 6840 13960 6960 13988
rect 7611 13960 7656 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 3970 13920 3976 13932
rect 3835 13892 3976 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 3050 13852 3056 13864
rect 2884 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13784 2927 13787
rect 3234 13784 3240 13796
rect 2915 13756 3240 13784
rect 2915 13753 2927 13756
rect 2869 13747 2927 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 3804 13784 3832 13883
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13920 4123 13923
rect 4338 13920 4344 13932
rect 4111 13892 4344 13920
rect 4111 13889 4123 13892
rect 4065 13883 4123 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4522 13920 4528 13932
rect 4483 13892 4528 13920
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 4798 13920 4804 13932
rect 4755 13892 4804 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 5092 13892 5365 13920
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 5092 13852 5120 13892
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 4212 13824 5120 13852
rect 5169 13855 5227 13861
rect 4212 13812 4218 13824
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5258 13852 5264 13864
rect 5215 13824 5264 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5460 13852 5488 13960
rect 6656 13932 6684 13960
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 6549 13923 6607 13929
rect 5684 13892 5729 13920
rect 5684 13880 5690 13892
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6564 13852 6592 13883
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 6932 13929 6960 13960
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 8110 13988 8116 14000
rect 7944 13960 8116 13988
rect 7098 13929 7104 13932
rect 6825 13923 6883 13929
rect 6696 13892 6789 13920
rect 6696 13880 6702 13892
rect 6825 13889 6837 13923
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 7055 13923 7104 13929
rect 7055 13889 7067 13923
rect 7101 13889 7104 13923
rect 7055 13883 7104 13889
rect 6730 13852 6736 13864
rect 5460 13824 6736 13852
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 4522 13784 4528 13796
rect 3804 13756 4528 13784
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 6840 13784 6868 13883
rect 7098 13880 7104 13883
rect 7156 13920 7162 13932
rect 7466 13920 7472 13932
rect 7156 13892 7472 13920
rect 7156 13880 7162 13892
rect 7466 13880 7472 13892
rect 7524 13920 7530 13932
rect 7944 13929 7972 13960
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7524 13892 7849 13920
rect 7524 13880 7530 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 8036 13852 8064 13883
rect 7248 13824 8064 13852
rect 7248 13812 7254 13824
rect 6512 13756 6868 13784
rect 6512 13744 6518 13756
rect 7944 13728 7972 13824
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3108 13688 3525 13716
rect 3108 13676 3114 13688
rect 3513 13685 3525 13688
rect 3559 13685 3571 13719
rect 3513 13679 3571 13685
rect 7926 13676 7932 13728
rect 7984 13676 7990 13728
rect 1104 13626 10856 13648
rect 1104 13574 2169 13626
rect 2221 13574 2233 13626
rect 2285 13574 2297 13626
rect 2349 13574 2361 13626
rect 2413 13574 2425 13626
rect 2477 13574 4607 13626
rect 4659 13574 4671 13626
rect 4723 13574 4735 13626
rect 4787 13574 4799 13626
rect 4851 13574 4863 13626
rect 4915 13574 7045 13626
rect 7097 13574 7109 13626
rect 7161 13574 7173 13626
rect 7225 13574 7237 13626
rect 7289 13574 7301 13626
rect 7353 13574 9483 13626
rect 9535 13574 9547 13626
rect 9599 13574 9611 13626
rect 9663 13574 9675 13626
rect 9727 13574 9739 13626
rect 9791 13574 10856 13626
rect 1104 13552 10856 13574
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7800 13484 8033 13512
rect 7800 13472 7806 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8021 13475 8079 13481
rect 7650 13444 7656 13456
rect 4908 13416 7656 13444
rect 3142 13376 3148 13388
rect 2516 13348 3148 13376
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2516 13317 2544 13348
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 4430 13336 4436 13388
rect 4488 13376 4494 13388
rect 4488 13348 4844 13376
rect 4488 13336 4494 13348
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 1912 13280 2329 13308
rect 1912 13268 1918 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13277 2559 13311
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2501 13271 2559 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 4154 13308 4160 13320
rect 3283 13280 4160 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4522 13308 4528 13320
rect 4483 13280 4528 13308
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4816 13317 4844 13348
rect 4908 13317 4936 13416
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5684 13348 6101 13376
rect 5684 13336 5690 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 7285 13379 7343 13385
rect 6319 13348 7236 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 4982 13308 4988 13320
rect 4939 13280 4988 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 7208 13317 7236 13348
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7834 13376 7840 13388
rect 7331 13348 7840 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7944 13348 8125 13376
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6512 13280 6561 13308
rect 6512 13268 6518 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7944 13308 7972 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 7239 13280 7972 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8076 13280 8121 13308
rect 8076 13268 8082 13280
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 3053 13243 3111 13249
rect 3053 13240 3065 13243
rect 2832 13212 3065 13240
rect 2832 13200 2838 13212
rect 3053 13209 3065 13212
rect 3099 13209 3111 13243
rect 4706 13240 4712 13252
rect 4667 13212 4712 13240
rect 3053 13203 3111 13209
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 7926 13240 7932 13252
rect 6472 13212 7932 13240
rect 2501 13175 2559 13181
rect 2501 13141 2513 13175
rect 2547 13172 2559 13175
rect 2958 13172 2964 13184
rect 2547 13144 2964 13172
rect 2547 13141 2559 13144
rect 2501 13135 2559 13141
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 3421 13175 3479 13181
rect 3421 13141 3433 13175
rect 3467 13172 3479 13175
rect 4062 13172 4068 13184
rect 3467 13144 4068 13172
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 6472 13181 6500 13212
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13141 6515 13175
rect 6457 13135 6515 13141
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 7834 13172 7840 13184
rect 7607 13144 7840 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 8389 13175 8447 13181
rect 8389 13141 8401 13175
rect 8435 13172 8447 13175
rect 8662 13172 8668 13184
rect 8435 13144 8668 13172
rect 8435 13141 8447 13144
rect 8389 13135 8447 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 1104 13082 11016 13104
rect 1104 13030 3388 13082
rect 3440 13030 3452 13082
rect 3504 13030 3516 13082
rect 3568 13030 3580 13082
rect 3632 13030 3644 13082
rect 3696 13030 5826 13082
rect 5878 13030 5890 13082
rect 5942 13030 5954 13082
rect 6006 13030 6018 13082
rect 6070 13030 6082 13082
rect 6134 13030 8264 13082
rect 8316 13030 8328 13082
rect 8380 13030 8392 13082
rect 8444 13030 8456 13082
rect 8508 13030 8520 13082
rect 8572 13030 10702 13082
rect 10754 13030 10766 13082
rect 10818 13030 10830 13082
rect 10882 13030 10894 13082
rect 10946 13030 10958 13082
rect 11010 13030 11016 13082
rect 1104 13008 11016 13030
rect 6454 12968 6460 12980
rect 5276 12940 6460 12968
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3605 12903 3663 12909
rect 3605 12900 3617 12903
rect 2832 12872 3617 12900
rect 2832 12860 2838 12872
rect 3605 12869 3617 12872
rect 3651 12869 3663 12903
rect 3605 12863 3663 12869
rect 4154 12860 4160 12912
rect 4212 12900 4218 12912
rect 5276 12900 5304 12940
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 4212 12872 5304 12900
rect 4212 12860 4218 12872
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3050 12832 3056 12844
rect 2915 12804 3056 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3878 12832 3884 12844
rect 3839 12804 3884 12832
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 4488 12804 4629 12832
rect 4488 12792 4494 12804
rect 4617 12801 4629 12804
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5276 12841 5304 12872
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 5626 12900 5632 12912
rect 5583 12872 5632 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 6549 12903 6607 12909
rect 6549 12869 6561 12903
rect 6595 12900 6607 12903
rect 6638 12900 6644 12912
rect 6595 12872 6644 12900
rect 6595 12869 6607 12872
rect 6549 12863 6607 12869
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 4764 12804 4813 12832
rect 4764 12792 4770 12804
rect 4801 12801 4813 12804
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 6564 12832 6592 12863
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 7650 12900 7656 12912
rect 6788 12872 6833 12900
rect 7300 12872 7656 12900
rect 6788 12860 6794 12872
rect 7300 12841 7328 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 5399 12804 6592 12832
rect 6825 12835 6883 12841
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 6825 12801 6837 12835
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7285 12795 7343 12801
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 3016 12736 3157 12764
rect 3016 12724 3022 12736
rect 3145 12733 3157 12736
rect 3191 12764 3203 12767
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3191 12736 3709 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 3053 12699 3111 12705
rect 3053 12696 3065 12699
rect 2832 12668 3065 12696
rect 2832 12656 2838 12668
rect 3053 12665 3065 12668
rect 3099 12665 3111 12699
rect 4816 12696 4844 12795
rect 6454 12724 6460 12776
rect 6512 12764 6518 12776
rect 6840 12764 6868 12795
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 6512 12736 6868 12764
rect 6512 12724 6518 12736
rect 8128 12696 8156 12792
rect 4816 12668 8156 12696
rect 3053 12659 3111 12665
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2648 12600 2697 12628
rect 2648 12588 2654 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 3234 12588 3240 12640
rect 3292 12628 3298 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3292 12600 3617 12628
rect 3292 12588 3298 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 3605 12591 3663 12597
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4154 12628 4160 12640
rect 4111 12600 4160 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4709 12631 4767 12637
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 5166 12628 5172 12640
rect 4755 12600 5172 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5350 12628 5356 12640
rect 5307 12600 5356 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 6641 12631 6699 12637
rect 6641 12597 6653 12631
rect 6687 12628 6699 12631
rect 6730 12628 6736 12640
rect 6687 12600 6736 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7650 12628 7656 12640
rect 7423 12600 7656 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8018 12628 8024 12640
rect 7979 12600 8024 12628
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 1104 12538 10856 12560
rect 1104 12486 2169 12538
rect 2221 12486 2233 12538
rect 2285 12486 2297 12538
rect 2349 12486 2361 12538
rect 2413 12486 2425 12538
rect 2477 12486 4607 12538
rect 4659 12486 4671 12538
rect 4723 12486 4735 12538
rect 4787 12486 4799 12538
rect 4851 12486 4863 12538
rect 4915 12486 7045 12538
rect 7097 12486 7109 12538
rect 7161 12486 7173 12538
rect 7225 12486 7237 12538
rect 7289 12486 7301 12538
rect 7353 12486 9483 12538
rect 9535 12486 9547 12538
rect 9599 12486 9611 12538
rect 9663 12486 9675 12538
rect 9727 12486 9739 12538
rect 9791 12486 10856 12538
rect 1104 12464 10856 12486
rect 7837 12359 7895 12365
rect 7837 12325 7849 12359
rect 7883 12356 7895 12359
rect 8573 12359 8631 12365
rect 7883 12328 8524 12356
rect 7883 12325 7895 12328
rect 7837 12319 7895 12325
rect 8496 12288 8524 12328
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 8846 12356 8852 12368
rect 8619 12328 8852 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 7576 12260 8432 12288
rect 8496 12260 8800 12288
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 3016 12192 3157 12220
rect 3016 12180 3022 12192
rect 3145 12189 3157 12192
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4580 12192 4629 12220
rect 4580 12180 4586 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4982 12220 4988 12232
rect 4847 12192 4988 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 7576 12229 7604 12260
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7837 12223 7895 12229
rect 7708 12192 7753 12220
rect 7708 12180 7714 12192
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8018 12220 8024 12232
rect 7883 12192 8024 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8018 12180 8024 12192
rect 8076 12220 8082 12232
rect 8404 12229 8432 12260
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8076 12192 8309 12220
rect 8076 12180 8082 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8662 12220 8668 12232
rect 8435 12192 8668 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8573 12155 8631 12161
rect 8573 12121 8585 12155
rect 8619 12152 8631 12155
rect 8772 12152 8800 12260
rect 9030 12152 9036 12164
rect 8619 12124 9036 12152
rect 8619 12121 8631 12124
rect 8573 12115 8631 12121
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 3050 12084 3056 12096
rect 3011 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4580 12056 4629 12084
rect 4580 12044 4586 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4617 12047 4675 12053
rect 1104 11994 11016 12016
rect 1104 11942 3388 11994
rect 3440 11942 3452 11994
rect 3504 11942 3516 11994
rect 3568 11942 3580 11994
rect 3632 11942 3644 11994
rect 3696 11942 5826 11994
rect 5878 11942 5890 11994
rect 5942 11942 5954 11994
rect 6006 11942 6018 11994
rect 6070 11942 6082 11994
rect 6134 11942 8264 11994
rect 8316 11942 8328 11994
rect 8380 11942 8392 11994
rect 8444 11942 8456 11994
rect 8508 11942 8520 11994
rect 8572 11942 10702 11994
rect 10754 11942 10766 11994
rect 10818 11942 10830 11994
rect 10882 11942 10894 11994
rect 10946 11942 10958 11994
rect 11010 11942 11016 11994
rect 1104 11920 11016 11942
rect 4154 11880 4160 11892
rect 4115 11852 4160 11880
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 6914 11880 6920 11892
rect 6871 11852 6920 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 5166 11812 5172 11824
rect 5127 11784 5172 11812
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 4062 11744 4068 11756
rect 4023 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4522 11744 4528 11756
rect 4387 11716 4528 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4522 11704 4528 11716
rect 4580 11744 4586 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4580 11716 4997 11744
rect 4580 11704 4586 11716
rect 4985 11713 4997 11716
rect 5031 11744 5043 11747
rect 5442 11744 5448 11756
rect 5031 11716 5448 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6730 11744 6736 11756
rect 6691 11716 6736 11744
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6886 11716 7021 11744
rect 6886 11688 6914 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 6822 11636 6828 11688
rect 6880 11648 6914 11688
rect 6880 11636 6886 11648
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4304 11512 4353 11540
rect 4304 11500 4310 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4488 11512 4813 11540
rect 4488 11500 4494 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7558 11540 7564 11552
rect 7055 11512 7564 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 1104 11450 10856 11472
rect 1104 11398 2169 11450
rect 2221 11398 2233 11450
rect 2285 11398 2297 11450
rect 2349 11398 2361 11450
rect 2413 11398 2425 11450
rect 2477 11398 4607 11450
rect 4659 11398 4671 11450
rect 4723 11398 4735 11450
rect 4787 11398 4799 11450
rect 4851 11398 4863 11450
rect 4915 11398 7045 11450
rect 7097 11398 7109 11450
rect 7161 11398 7173 11450
rect 7225 11398 7237 11450
rect 7289 11398 7301 11450
rect 7353 11398 9483 11450
rect 9535 11398 9547 11450
rect 9599 11398 9611 11450
rect 9663 11398 9675 11450
rect 9727 11398 9739 11450
rect 9791 11398 10856 11450
rect 1104 11376 10856 11398
rect 5350 11336 5356 11348
rect 4172 11308 5356 11336
rect 4172 11209 4200 11308
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 6822 11336 6828 11348
rect 6779 11308 6828 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 4433 11271 4491 11277
rect 4433 11237 4445 11271
rect 4479 11268 4491 11271
rect 4982 11268 4988 11280
rect 4479 11240 4988 11268
rect 4479 11237 4491 11240
rect 4433 11231 4491 11237
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 5166 11228 5172 11280
rect 5224 11268 5230 11280
rect 5224 11240 6224 11268
rect 5224 11228 5230 11240
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11169 4215 11203
rect 5074 11200 5080 11212
rect 4157 11163 4215 11169
rect 4448 11172 5080 11200
rect 4448 11141 4476 11172
rect 5074 11160 5080 11172
rect 5132 11200 5138 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 5132 11172 5273 11200
rect 5132 11160 5138 11172
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 5491 11172 6101 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6196 11200 6224 11240
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6196 11172 7113 11200
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 5166 11132 5172 11144
rect 4571 11104 5172 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5350 11132 5356 11144
rect 5311 11104 5356 11132
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 6196 11141 6224 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5592 11104 6009 11132
rect 5592 11092 5598 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7116 11132 7144 11163
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 7116 11104 7665 11132
rect 7009 11095 7067 11101
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 5718 11064 5724 11076
rect 5000 11036 5724 11064
rect 4338 10996 4344 11008
rect 4299 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 5000 11005 5028 11036
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 7024 11064 7052 11095
rect 7742 11092 7748 11144
rect 7800 11132 7806 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7800 11104 7849 11132
rect 7800 11092 7806 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7760 11064 7788 11092
rect 7024 11036 7788 11064
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10965 5043 10999
rect 4985 10959 5043 10965
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7524 10968 7757 10996
rect 7524 10956 7530 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 1104 10906 11016 10928
rect 1104 10854 3388 10906
rect 3440 10854 3452 10906
rect 3504 10854 3516 10906
rect 3568 10854 3580 10906
rect 3632 10854 3644 10906
rect 3696 10854 5826 10906
rect 5878 10854 5890 10906
rect 5942 10854 5954 10906
rect 6006 10854 6018 10906
rect 6070 10854 6082 10906
rect 6134 10854 8264 10906
rect 8316 10854 8328 10906
rect 8380 10854 8392 10906
rect 8444 10854 8456 10906
rect 8508 10854 8520 10906
rect 8572 10854 10702 10906
rect 10754 10854 10766 10906
rect 10818 10854 10830 10906
rect 10882 10854 10894 10906
rect 10946 10854 10958 10906
rect 11010 10854 11016 10906
rect 1104 10832 11016 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4173 10795 4231 10801
rect 4173 10792 4185 10795
rect 4120 10764 4185 10792
rect 4120 10752 4126 10764
rect 4173 10761 4185 10764
rect 4219 10761 4231 10795
rect 4522 10792 4528 10804
rect 4173 10755 4231 10761
rect 4264 10764 4528 10792
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10724 4031 10727
rect 4264 10724 4292 10764
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7650 10792 7656 10804
rect 6972 10764 7656 10792
rect 6972 10752 6978 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 4019 10696 4292 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 4338 10684 4344 10736
rect 4396 10724 4402 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4396 10696 5089 10724
rect 4396 10684 4402 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 6822 10724 6828 10736
rect 5224 10696 5269 10724
rect 6748 10696 6828 10724
rect 5224 10684 5230 10696
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 5350 10656 5356 10668
rect 5311 10628 5356 10656
rect 4985 10619 5043 10625
rect 5000 10588 5028 10619
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 6748 10665 6776 10696
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7009 10619 7067 10625
rect 5074 10588 5080 10600
rect 5000 10560 5080 10588
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7024 10520 7052 10619
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7745 10659 7803 10665
rect 7616 10628 7661 10656
rect 7616 10616 7622 10628
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 7834 10656 7840 10668
rect 7791 10628 7840 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 7834 10616 7840 10628
rect 7892 10656 7898 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 7892 10628 8401 10656
rect 7892 10616 7898 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 7484 10588 7512 10616
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 7484 10560 8493 10588
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 6788 10492 7052 10520
rect 6788 10480 6794 10492
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 7616 10492 8432 10520
rect 7616 10480 7622 10492
rect 4154 10452 4160 10464
rect 4115 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4338 10452 4344 10464
rect 4299 10424 4344 10452
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5074 10452 5080 10464
rect 4847 10424 5080 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6638 10452 6644 10464
rect 6595 10424 6644 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 8202 10452 8208 10464
rect 7975 10424 8208 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8404 10461 8432 10492
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10421 8447 10455
rect 8754 10452 8760 10464
rect 8715 10424 8760 10452
rect 8389 10415 8447 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 1104 10362 10856 10384
rect 1104 10310 2169 10362
rect 2221 10310 2233 10362
rect 2285 10310 2297 10362
rect 2349 10310 2361 10362
rect 2413 10310 2425 10362
rect 2477 10310 4607 10362
rect 4659 10310 4671 10362
rect 4723 10310 4735 10362
rect 4787 10310 4799 10362
rect 4851 10310 4863 10362
rect 4915 10310 7045 10362
rect 7097 10310 7109 10362
rect 7161 10310 7173 10362
rect 7225 10310 7237 10362
rect 7289 10310 7301 10362
rect 7353 10310 9483 10362
rect 9535 10310 9547 10362
rect 9599 10310 9611 10362
rect 9663 10310 9675 10362
rect 9727 10310 9739 10362
rect 9791 10310 10856 10362
rect 1104 10288 10856 10310
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 5040 10220 5089 10248
rect 5040 10208 5046 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 5077 10211 5135 10217
rect 6196 10220 6837 10248
rect 4246 10112 4252 10124
rect 4172 10084 4252 10112
rect 4172 10053 4200 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4157 10007 4215 10013
rect 4172 9976 4200 10007
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 6196 10053 6224 10220
rect 6825 10217 6837 10220
rect 6871 10248 6883 10251
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 6871 10220 7481 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 6822 10072 6828 10124
rect 6880 10072 6886 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 6972 10084 7788 10112
rect 6972 10072 6978 10084
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5776 10016 5917 10044
rect 5776 10004 5782 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 4890 9976 4896 9988
rect 4172 9948 4896 9976
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 5074 9936 5080 9988
rect 5132 9985 5138 9988
rect 5132 9979 5151 9985
rect 5139 9945 5151 9979
rect 5132 9939 5151 9945
rect 5132 9936 5138 9939
rect 4246 9908 4252 9920
rect 4207 9880 4252 9908
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5718 9908 5724 9920
rect 5679 9880 5724 9908
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 5920 9908 5948 10007
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 6638 9976 6644 9988
rect 6135 9948 6644 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 6840 9976 6868 10072
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 7650 10044 7656 10056
rect 7607 10016 7656 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 7484 9976 7512 10007
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7760 10053 7788 10084
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 7745 10007 7803 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 6840 9948 7512 9976
rect 6841 9911 6899 9917
rect 6841 9908 6853 9911
rect 5920 9880 6853 9908
rect 6841 9877 6853 9880
rect 6887 9877 6899 9911
rect 7006 9908 7012 9920
rect 6967 9880 7012 9908
rect 6841 9871 6899 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8662 9908 8668 9920
rect 8343 9880 8668 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 4801 9707 4859 9713
rect 4801 9673 4813 9707
rect 4847 9704 4859 9707
rect 4982 9704 4988 9716
rect 4847 9676 4988 9704
rect 4847 9673 4859 9676
rect 4801 9667 4859 9673
rect 4982 9664 4988 9676
rect 5040 9664 5046 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 5776 9676 6653 9704
rect 5776 9664 5782 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 8754 9664 8760 9716
rect 8812 9664 8818 9716
rect 5074 9636 5080 9648
rect 4724 9608 5080 9636
rect 4724 9577 4752 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5997 9639 6055 9645
rect 5997 9605 6009 9639
rect 6043 9636 6055 9639
rect 7929 9639 7987 9645
rect 6043 9608 6868 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4948 9540 4997 9568
rect 4948 9528 4954 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 6840 9577 6868 9608
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8570 9636 8576 9648
rect 7975 9608 8576 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8570 9596 8576 9608
rect 8628 9636 8634 9648
rect 8772 9636 8800 9664
rect 8628 9608 8800 9636
rect 8628 9596 8634 9608
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 8904 9608 8949 9636
rect 8904 9596 8910 9608
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5316 9540 6561 9568
rect 5316 9528 5322 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7006 9568 7012 9580
rect 6871 9540 7012 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 8110 9568 8116 9580
rect 8071 9540 8116 9568
rect 7837 9531 7895 9537
rect 7466 9500 7472 9512
rect 7024 9472 7472 9500
rect 5718 9432 5724 9444
rect 5679 9404 5724 9432
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 7024 9441 7052 9472
rect 7466 9460 7472 9472
rect 7524 9500 7530 9512
rect 7852 9500 7880 9531
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 9030 9568 9036 9580
rect 8991 9540 9036 9568
rect 8757 9531 8815 9537
rect 7524 9472 7880 9500
rect 7524 9460 7530 9472
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 8772 9376 8800 9531
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 4982 9364 4988 9376
rect 4943 9336 4988 9364
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8754 9364 8760 9376
rect 8343 9336 8760 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 10042 9364 10048 9376
rect 9263 9336 10048 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5276 8996 5733 9024
rect 5276 8968 5304 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6730 9024 6736 9036
rect 6227 8996 6736 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7466 9024 7472 9036
rect 7427 8996 7472 9024
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 8662 9024 8668 9036
rect 8404 8996 8668 9024
rect 4982 8956 4988 8968
rect 4943 8928 4988 8956
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 8404 8965 8432 8996
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 8389 8919 8447 8925
rect 7576 8888 7604 8919
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 7576 8860 8493 8888
rect 8481 8857 8493 8860
rect 8527 8857 8539 8891
rect 8481 8851 8539 8857
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 5258 8820 5264 8832
rect 5123 8792 5264 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 7926 8820 7932 8832
rect 7887 8792 7932 8820
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 8846 8548 8852 8560
rect 8404 8520 8852 8548
rect 8404 8489 8432 8520
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8772 8412 8800 8440
rect 8527 8384 8800 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9950 8344 9956 8356
rect 8803 8316 9956 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 10042 3040 10048 3052
rect 10003 3012 10048 3040
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 11054 2836 11060 2848
rect 10275 2808 11060 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 3050 2496 3056 2508
rect 1872 2468 3056 2496
rect 1872 2437 1900 2468
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 1857 2391 1915 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7984 2400 8217 2428
rect 7984 2388 7990 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9950 2428 9956 2440
rect 9723 2400 9956 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 750 2252 756 2304
rect 808 2292 814 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 808 2264 1685 2292
rect 808 2252 814 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 2222 2252 2228 2304
rect 2280 2292 2286 2304
rect 2409 2295 2467 2301
rect 2409 2292 2421 2295
rect 2280 2264 2421 2292
rect 2280 2252 2286 2264
rect 2409 2261 2421 2264
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3844 2264 4077 2292
rect 3844 2252 3850 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6696 2264 6929 2292
rect 6696 2252 6702 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 6917 2255 6975 2261
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 8389 2295 8447 2301
rect 8389 2292 8401 2295
rect 8168 2264 8401 2292
rect 8168 2252 8174 2264
rect 8389 2261 8401 2264
rect 8435 2261 8447 2295
rect 8389 2255 8447 2261
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9640 2264 9873 2292
rect 9640 2252 9646 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
<< via1 >>
rect 2169 15750 2221 15802
rect 2233 15750 2285 15802
rect 2297 15750 2349 15802
rect 2361 15750 2413 15802
rect 2425 15750 2477 15802
rect 4607 15750 4659 15802
rect 4671 15750 4723 15802
rect 4735 15750 4787 15802
rect 4799 15750 4851 15802
rect 4863 15750 4915 15802
rect 7045 15750 7097 15802
rect 7109 15750 7161 15802
rect 7173 15750 7225 15802
rect 7237 15750 7289 15802
rect 7301 15750 7353 15802
rect 9483 15750 9535 15802
rect 9547 15750 9599 15802
rect 9611 15750 9663 15802
rect 9675 15750 9727 15802
rect 9739 15750 9791 15802
rect 2504 15512 2556 15564
rect 8116 15512 8168 15564
rect 8668 15512 8720 15564
rect 9404 15512 9456 15564
rect 2044 15444 2096 15496
rect 4160 15444 4212 15496
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 6644 15444 6696 15496
rect 5724 15376 5776 15428
rect 6184 15376 6236 15428
rect 7656 15376 7708 15428
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 3388 15206 3440 15258
rect 3452 15206 3504 15258
rect 3516 15206 3568 15258
rect 3580 15206 3632 15258
rect 3644 15206 3696 15258
rect 5826 15206 5878 15258
rect 5890 15206 5942 15258
rect 5954 15206 6006 15258
rect 6018 15206 6070 15258
rect 6082 15206 6134 15258
rect 8264 15206 8316 15258
rect 8328 15206 8380 15258
rect 8392 15206 8444 15258
rect 8456 15206 8508 15258
rect 8520 15206 8572 15258
rect 10702 15206 10754 15258
rect 10766 15206 10818 15258
rect 10830 15206 10882 15258
rect 10894 15206 10946 15258
rect 10958 15206 11010 15258
rect 4160 15104 4212 15156
rect 6184 15104 6236 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 1032 14968 1084 15020
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 5540 14968 5592 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 10324 15011 10376 15020
rect 5816 14968 5868 14977
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 11060 14968 11112 15020
rect 4344 14900 4396 14952
rect 6920 14900 6972 14952
rect 8116 14900 8168 14952
rect 3884 14764 3936 14816
rect 5632 14764 5684 14816
rect 2169 14662 2221 14714
rect 2233 14662 2285 14714
rect 2297 14662 2349 14714
rect 2361 14662 2413 14714
rect 2425 14662 2477 14714
rect 4607 14662 4659 14714
rect 4671 14662 4723 14714
rect 4735 14662 4787 14714
rect 4799 14662 4851 14714
rect 4863 14662 4915 14714
rect 7045 14662 7097 14714
rect 7109 14662 7161 14714
rect 7173 14662 7225 14714
rect 7237 14662 7289 14714
rect 7301 14662 7353 14714
rect 9483 14662 9535 14714
rect 9547 14662 9599 14714
rect 9611 14662 9663 14714
rect 9675 14662 9727 14714
rect 9739 14662 9791 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 5724 14560 5776 14612
rect 9404 14560 9456 14612
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 3056 14424 3108 14476
rect 3148 14356 3200 14408
rect 3332 14356 3384 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4528 14424 4580 14476
rect 2320 14288 2372 14340
rect 3792 14288 3844 14340
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 5724 14399 5776 14408
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 6184 14424 6236 14476
rect 6736 14356 6788 14408
rect 4160 14288 4212 14340
rect 4804 14288 4856 14340
rect 7656 14492 7708 14544
rect 7748 14399 7800 14408
rect 2964 14220 3016 14272
rect 3332 14220 3384 14272
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 5816 14220 5868 14272
rect 7104 14331 7156 14340
rect 7104 14297 7113 14331
rect 7113 14297 7147 14331
rect 7147 14297 7156 14331
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 7104 14288 7156 14297
rect 8116 14288 8168 14340
rect 7196 14220 7248 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 3388 14118 3440 14170
rect 3452 14118 3504 14170
rect 3516 14118 3568 14170
rect 3580 14118 3632 14170
rect 3644 14118 3696 14170
rect 5826 14118 5878 14170
rect 5890 14118 5942 14170
rect 5954 14118 6006 14170
rect 6018 14118 6070 14170
rect 6082 14118 6134 14170
rect 8264 14118 8316 14170
rect 8328 14118 8380 14170
rect 8392 14118 8444 14170
rect 8456 14118 8508 14170
rect 8520 14118 8572 14170
rect 10702 14118 10754 14170
rect 10766 14118 10818 14170
rect 10830 14118 10882 14170
rect 10894 14118 10946 14170
rect 10958 14118 11010 14170
rect 2044 14016 2096 14068
rect 1860 13948 1912 14000
rect 4436 14016 4488 14068
rect 5540 14059 5592 14068
rect 5540 14025 5549 14059
rect 5549 14025 5583 14059
rect 5583 14025 5592 14059
rect 5540 14016 5592 14025
rect 6828 14016 6880 14068
rect 6920 14016 6972 14068
rect 7932 14016 7984 14068
rect 2044 13880 2096 13932
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 3700 13923 3752 13932
rect 2780 13812 2832 13864
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 7656 13991 7708 14000
rect 3056 13812 3108 13864
rect 3240 13744 3292 13796
rect 3976 13880 4028 13932
rect 4344 13880 4396 13932
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4804 13880 4856 13932
rect 4160 13812 4212 13864
rect 5264 13812 5316 13864
rect 5632 13923 5684 13932
rect 5632 13889 5641 13923
rect 5641 13889 5675 13923
rect 5675 13889 5684 13923
rect 5632 13880 5684 13889
rect 6644 13923 6696 13932
rect 6644 13889 6654 13923
rect 6654 13889 6688 13923
rect 6688 13889 6696 13923
rect 7656 13957 7665 13991
rect 7665 13957 7699 13991
rect 7699 13957 7708 13991
rect 7656 13948 7708 13957
rect 6644 13880 6696 13889
rect 6736 13812 6788 13864
rect 4528 13744 4580 13796
rect 6460 13744 6512 13796
rect 7104 13880 7156 13932
rect 7472 13880 7524 13932
rect 8116 13948 8168 14000
rect 7196 13812 7248 13864
rect 3056 13676 3108 13728
rect 7932 13676 7984 13728
rect 2169 13574 2221 13626
rect 2233 13574 2285 13626
rect 2297 13574 2349 13626
rect 2361 13574 2413 13626
rect 2425 13574 2477 13626
rect 4607 13574 4659 13626
rect 4671 13574 4723 13626
rect 4735 13574 4787 13626
rect 4799 13574 4851 13626
rect 4863 13574 4915 13626
rect 7045 13574 7097 13626
rect 7109 13574 7161 13626
rect 7173 13574 7225 13626
rect 7237 13574 7289 13626
rect 7301 13574 7353 13626
rect 9483 13574 9535 13626
rect 9547 13574 9599 13626
rect 9611 13574 9663 13626
rect 9675 13574 9727 13626
rect 9739 13574 9791 13626
rect 7748 13472 7800 13524
rect 1860 13268 1912 13320
rect 3148 13336 3200 13388
rect 4436 13336 4488 13388
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4160 13268 4212 13320
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 7656 13404 7708 13456
rect 5632 13336 5684 13388
rect 4988 13268 5040 13320
rect 6460 13268 6512 13320
rect 7840 13336 7892 13388
rect 8024 13311 8076 13320
rect 8024 13277 8033 13311
rect 8033 13277 8067 13311
rect 8067 13277 8076 13311
rect 8024 13268 8076 13277
rect 2780 13200 2832 13252
rect 4712 13243 4764 13252
rect 4712 13209 4721 13243
rect 4721 13209 4755 13243
rect 4755 13209 4764 13243
rect 4712 13200 4764 13209
rect 2964 13132 3016 13184
rect 4068 13132 4120 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 5080 13132 5132 13141
rect 7932 13200 7984 13252
rect 7840 13132 7892 13184
rect 8668 13132 8720 13184
rect 3388 13030 3440 13082
rect 3452 13030 3504 13082
rect 3516 13030 3568 13082
rect 3580 13030 3632 13082
rect 3644 13030 3696 13082
rect 5826 13030 5878 13082
rect 5890 13030 5942 13082
rect 5954 13030 6006 13082
rect 6018 13030 6070 13082
rect 6082 13030 6134 13082
rect 8264 13030 8316 13082
rect 8328 13030 8380 13082
rect 8392 13030 8444 13082
rect 8456 13030 8508 13082
rect 8520 13030 8572 13082
rect 10702 13030 10754 13082
rect 10766 13030 10818 13082
rect 10830 13030 10882 13082
rect 10894 13030 10946 13082
rect 10958 13030 11010 13082
rect 2780 12860 2832 12912
rect 4160 12860 4212 12912
rect 6460 12928 6512 12980
rect 3056 12792 3108 12844
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 4436 12792 4488 12844
rect 4712 12792 4764 12844
rect 5632 12860 5684 12912
rect 6644 12860 6696 12912
rect 6736 12903 6788 12912
rect 6736 12869 6745 12903
rect 6745 12869 6779 12903
rect 6779 12869 6788 12903
rect 6736 12860 6788 12869
rect 7656 12860 7708 12912
rect 7472 12835 7524 12844
rect 2964 12724 3016 12776
rect 2780 12656 2832 12708
rect 6460 12724 6512 12776
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 2596 12588 2648 12640
rect 3240 12588 3292 12640
rect 4160 12588 4212 12640
rect 5172 12588 5224 12640
rect 5356 12588 5408 12640
rect 6736 12588 6788 12640
rect 7656 12588 7708 12640
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 2169 12486 2221 12538
rect 2233 12486 2285 12538
rect 2297 12486 2349 12538
rect 2361 12486 2413 12538
rect 2425 12486 2477 12538
rect 4607 12486 4659 12538
rect 4671 12486 4723 12538
rect 4735 12486 4787 12538
rect 4799 12486 4851 12538
rect 4863 12486 4915 12538
rect 7045 12486 7097 12538
rect 7109 12486 7161 12538
rect 7173 12486 7225 12538
rect 7237 12486 7289 12538
rect 7301 12486 7353 12538
rect 9483 12486 9535 12538
rect 9547 12486 9599 12538
rect 9611 12486 9663 12538
rect 9675 12486 9727 12538
rect 9739 12486 9791 12538
rect 8852 12316 8904 12368
rect 2964 12180 3016 12232
rect 4528 12180 4580 12232
rect 4988 12180 5040 12232
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 8024 12180 8076 12232
rect 8668 12180 8720 12232
rect 9036 12112 9088 12164
rect 3056 12087 3108 12096
rect 3056 12053 3065 12087
rect 3065 12053 3099 12087
rect 3099 12053 3108 12087
rect 3056 12044 3108 12053
rect 4528 12044 4580 12096
rect 3388 11942 3440 11994
rect 3452 11942 3504 11994
rect 3516 11942 3568 11994
rect 3580 11942 3632 11994
rect 3644 11942 3696 11994
rect 5826 11942 5878 11994
rect 5890 11942 5942 11994
rect 5954 11942 6006 11994
rect 6018 11942 6070 11994
rect 6082 11942 6134 11994
rect 8264 11942 8316 11994
rect 8328 11942 8380 11994
rect 8392 11942 8444 11994
rect 8456 11942 8508 11994
rect 8520 11942 8572 11994
rect 10702 11942 10754 11994
rect 10766 11942 10818 11994
rect 10830 11942 10882 11994
rect 10894 11942 10946 11994
rect 10958 11942 11010 11994
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 6920 11840 6972 11892
rect 5172 11815 5224 11824
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 4528 11704 4580 11756
rect 5448 11704 5500 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 6828 11636 6880 11688
rect 4252 11500 4304 11552
rect 4436 11500 4488 11552
rect 7564 11500 7616 11552
rect 2169 11398 2221 11450
rect 2233 11398 2285 11450
rect 2297 11398 2349 11450
rect 2361 11398 2413 11450
rect 2425 11398 2477 11450
rect 4607 11398 4659 11450
rect 4671 11398 4723 11450
rect 4735 11398 4787 11450
rect 4799 11398 4851 11450
rect 4863 11398 4915 11450
rect 7045 11398 7097 11450
rect 7109 11398 7161 11450
rect 7173 11398 7225 11450
rect 7237 11398 7289 11450
rect 7301 11398 7353 11450
rect 9483 11398 9535 11450
rect 9547 11398 9599 11450
rect 9611 11398 9663 11450
rect 9675 11398 9727 11450
rect 9739 11398 9791 11450
rect 5356 11296 5408 11348
rect 6828 11296 6880 11348
rect 4988 11228 5040 11280
rect 5172 11228 5224 11280
rect 5080 11160 5132 11212
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 5540 11092 5592 11144
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 5724 11024 5776 11076
rect 7748 11092 7800 11144
rect 7472 10956 7524 11008
rect 3388 10854 3440 10906
rect 3452 10854 3504 10906
rect 3516 10854 3568 10906
rect 3580 10854 3632 10906
rect 3644 10854 3696 10906
rect 5826 10854 5878 10906
rect 5890 10854 5942 10906
rect 5954 10854 6006 10906
rect 6018 10854 6070 10906
rect 6082 10854 6134 10906
rect 8264 10854 8316 10906
rect 8328 10854 8380 10906
rect 8392 10854 8444 10906
rect 8456 10854 8508 10906
rect 8520 10854 8572 10906
rect 10702 10854 10754 10906
rect 10766 10854 10818 10906
rect 10830 10854 10882 10906
rect 10894 10854 10946 10906
rect 10958 10854 11010 10906
rect 4068 10752 4120 10804
rect 4528 10752 4580 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7656 10752 7708 10804
rect 4344 10684 4396 10736
rect 5172 10727 5224 10736
rect 5172 10693 5181 10727
rect 5181 10693 5215 10727
rect 5215 10693 5224 10727
rect 5172 10684 5224 10693
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 6828 10684 6880 10736
rect 7472 10659 7524 10668
rect 5080 10548 5132 10600
rect 6736 10480 6788 10532
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 7840 10616 7892 10668
rect 7564 10480 7616 10532
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 4344 10455 4396 10464
rect 4344 10421 4353 10455
rect 4353 10421 4387 10455
rect 4387 10421 4396 10455
rect 4344 10412 4396 10421
rect 5080 10412 5132 10464
rect 6644 10412 6696 10464
rect 8208 10412 8260 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 2169 10310 2221 10362
rect 2233 10310 2285 10362
rect 2297 10310 2349 10362
rect 2361 10310 2413 10362
rect 2425 10310 2477 10362
rect 4607 10310 4659 10362
rect 4671 10310 4723 10362
rect 4735 10310 4787 10362
rect 4799 10310 4851 10362
rect 4863 10310 4915 10362
rect 7045 10310 7097 10362
rect 7109 10310 7161 10362
rect 7173 10310 7225 10362
rect 7237 10310 7289 10362
rect 7301 10310 7353 10362
rect 9483 10310 9535 10362
rect 9547 10310 9599 10362
rect 9611 10310 9663 10362
rect 9675 10310 9727 10362
rect 9739 10310 9791 10362
rect 4988 10208 5040 10260
rect 4252 10072 4304 10124
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 5724 10004 5776 10056
rect 6828 10072 6880 10124
rect 6920 10072 6972 10124
rect 4896 9979 4948 9988
rect 4896 9945 4905 9979
rect 4905 9945 4939 9979
rect 4939 9945 4948 9979
rect 4896 9936 4948 9945
rect 5080 9979 5132 9988
rect 5080 9945 5105 9979
rect 5105 9945 5132 9979
rect 5080 9936 5132 9945
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6644 9979 6696 9988
rect 6644 9945 6653 9979
rect 6653 9945 6687 9979
rect 6687 9945 6696 9979
rect 6644 9936 6696 9945
rect 7656 10004 7708 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7012 9868 7064 9877
rect 8668 9868 8720 9920
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 4988 9664 5040 9716
rect 5724 9664 5776 9716
rect 8760 9664 8812 9716
rect 5080 9596 5132 9648
rect 4896 9528 4948 9580
rect 5264 9528 5316 9580
rect 8576 9596 8628 9648
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 7012 9528 7064 9580
rect 8116 9571 8168 9580
rect 5724 9435 5776 9444
rect 5724 9401 5733 9435
rect 5733 9401 5767 9435
rect 5767 9401 5776 9435
rect 5724 9392 5776 9401
rect 7472 9460 7524 9512
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 5816 9324 5868 9376
rect 8760 9324 8812 9376
rect 10048 9324 10100 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 6736 8984 6788 9036
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 5264 8916 5316 8968
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 8668 8984 8720 9036
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 5264 8780 5316 8832
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 8852 8508 8904 8560
rect 8760 8440 8812 8492
rect 9956 8304 10008 8356
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 11060 2796 11112 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 3056 2456 3108 2508
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 7932 2388 7984 2440
rect 9956 2388 10008 2440
rect 756 2252 808 2304
rect 2228 2252 2280 2304
rect 3792 2252 3844 2304
rect 5172 2252 5224 2304
rect 6644 2252 6696 2304
rect 8116 2252 8168 2304
rect 9588 2252 9640 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
<< metal2 >>
rect 754 17354 810 18000
rect 2226 17354 2282 18000
rect 3698 17354 3754 18000
rect 5170 17354 5226 18000
rect 754 17326 1072 17354
rect 754 17200 810 17326
rect 1044 15026 1072 17326
rect 2226 17326 2544 17354
rect 2226 17200 2282 17326
rect 2169 15804 2477 15813
rect 2169 15802 2175 15804
rect 2231 15802 2255 15804
rect 2311 15802 2335 15804
rect 2391 15802 2415 15804
rect 2471 15802 2477 15804
rect 2231 15750 2233 15802
rect 2413 15750 2415 15802
rect 2169 15748 2175 15750
rect 2231 15748 2255 15750
rect 2311 15748 2335 15750
rect 2391 15748 2415 15750
rect 2471 15748 2477 15750
rect 2169 15739 2477 15748
rect 2516 15570 2544 17326
rect 3698 17326 4108 17354
rect 3698 17200 3754 17326
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 4080 15450 4108 17326
rect 5170 17326 5396 17354
rect 5170 17200 5226 17326
rect 4607 15804 4915 15813
rect 4607 15802 4613 15804
rect 4669 15802 4693 15804
rect 4749 15802 4773 15804
rect 4829 15802 4853 15804
rect 4909 15802 4915 15804
rect 4669 15750 4671 15802
rect 4851 15750 4853 15802
rect 4607 15748 4613 15750
rect 4669 15748 4693 15750
rect 4749 15748 4773 15750
rect 4829 15748 4853 15750
rect 4909 15748 4915 15750
rect 4607 15739 4915 15748
rect 5368 15502 5396 17326
rect 6642 17200 6698 18000
rect 8114 17200 8170 18000
rect 9586 17354 9642 18000
rect 9416 17326 9642 17354
rect 6656 15502 6684 17200
rect 7045 15804 7353 15813
rect 7045 15802 7051 15804
rect 7107 15802 7131 15804
rect 7187 15802 7211 15804
rect 7267 15802 7291 15804
rect 7347 15802 7353 15804
rect 7107 15750 7109 15802
rect 7289 15750 7291 15802
rect 7045 15748 7051 15750
rect 7107 15748 7131 15750
rect 7187 15748 7211 15750
rect 7267 15748 7291 15750
rect 7347 15748 7353 15750
rect 7045 15739 7353 15748
rect 8128 15570 8156 17200
rect 9416 15570 9444 17326
rect 9586 17200 9642 17326
rect 11058 17200 11114 18000
rect 9483 15804 9791 15813
rect 9483 15802 9489 15804
rect 9545 15802 9569 15804
rect 9625 15802 9649 15804
rect 9705 15802 9729 15804
rect 9785 15802 9791 15804
rect 9545 15750 9547 15802
rect 9727 15750 9729 15802
rect 9483 15748 9489 15750
rect 9545 15748 9569 15750
rect 9625 15748 9649 15750
rect 9705 15748 9729 15750
rect 9785 15748 9791 15750
rect 9483 15739 9791 15748
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 4160 15496 4212 15502
rect 4080 15444 4160 15450
rect 4080 15438 4212 15444
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 1032 15020 1084 15026
rect 1032 14962 1084 14968
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14618 1624 14962
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1872 14006 1900 14894
rect 2056 14074 2084 15438
rect 4080 15422 4200 15438
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3388 15260 3696 15269
rect 3388 15258 3394 15260
rect 3450 15258 3474 15260
rect 3530 15258 3554 15260
rect 3610 15258 3634 15260
rect 3690 15258 3696 15260
rect 3450 15206 3452 15258
rect 3632 15206 3634 15258
rect 3388 15204 3394 15206
rect 3450 15204 3474 15206
rect 3530 15204 3554 15206
rect 3610 15204 3634 15206
rect 3690 15204 3696 15206
rect 3388 15195 3696 15204
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 2169 14716 2477 14725
rect 2169 14714 2175 14716
rect 2231 14714 2255 14716
rect 2311 14714 2335 14716
rect 2391 14714 2415 14716
rect 2471 14714 2477 14716
rect 2231 14662 2233 14714
rect 2413 14662 2415 14714
rect 2169 14660 2175 14662
rect 2231 14660 2255 14662
rect 2311 14660 2335 14662
rect 2391 14660 2415 14662
rect 2471 14660 2477 14662
rect 2169 14651 2477 14660
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1872 13326 1900 13942
rect 2056 13938 2084 14010
rect 2332 13938 2360 14282
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2169 13628 2477 13637
rect 2169 13626 2175 13628
rect 2231 13626 2255 13628
rect 2311 13626 2335 13628
rect 2391 13626 2415 13628
rect 2471 13626 2477 13628
rect 2231 13574 2233 13626
rect 2413 13574 2415 13626
rect 2169 13572 2175 13574
rect 2231 13572 2255 13574
rect 2311 13572 2335 13574
rect 2391 13572 2415 13574
rect 2471 13572 2477 13574
rect 2169 13563 2477 13572
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 2792 13258 2820 13806
rect 2976 13326 3004 14214
rect 3068 13870 3096 14418
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12918 2820 13194
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2792 12714 2820 12854
rect 2976 12782 3004 13126
rect 3068 12850 3096 13670
rect 3160 13394 3188 14350
rect 3344 14278 3372 14350
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3388 14172 3696 14181
rect 3388 14170 3394 14172
rect 3450 14170 3474 14172
rect 3530 14170 3554 14172
rect 3610 14170 3634 14172
rect 3690 14170 3696 14172
rect 3450 14118 3452 14170
rect 3632 14118 3634 14170
rect 3388 14116 3394 14118
rect 3450 14116 3474 14118
rect 3530 14116 3554 14118
rect 3610 14116 3634 14118
rect 3690 14116 3696 14118
rect 3388 14107 3696 14116
rect 3700 13932 3752 13938
rect 3804 13920 3832 14282
rect 3752 13892 3832 13920
rect 3700 13874 3752 13880
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2169 12540 2477 12549
rect 2169 12538 2175 12540
rect 2231 12538 2255 12540
rect 2311 12538 2335 12540
rect 2391 12538 2415 12540
rect 2471 12538 2477 12540
rect 2231 12486 2233 12538
rect 2413 12486 2415 12538
rect 2169 12484 2175 12486
rect 2231 12484 2255 12486
rect 2311 12484 2335 12486
rect 2391 12484 2415 12486
rect 2471 12484 2477 12486
rect 2169 12475 2477 12484
rect 2169 11452 2477 11461
rect 2169 11450 2175 11452
rect 2231 11450 2255 11452
rect 2311 11450 2335 11452
rect 2391 11450 2415 11452
rect 2471 11450 2477 11452
rect 2231 11398 2233 11450
rect 2413 11398 2415 11450
rect 2169 11396 2175 11398
rect 2231 11396 2255 11398
rect 2311 11396 2335 11398
rect 2391 11396 2415 11398
rect 2471 11396 2477 11398
rect 2169 11387 2477 11396
rect 2169 10364 2477 10373
rect 2169 10362 2175 10364
rect 2231 10362 2255 10364
rect 2311 10362 2335 10364
rect 2391 10362 2415 10364
rect 2471 10362 2477 10364
rect 2231 10310 2233 10362
rect 2413 10310 2415 10362
rect 2169 10308 2175 10310
rect 2231 10308 2255 10310
rect 2311 10308 2335 10310
rect 2391 10308 2415 10310
rect 2471 10308 2477 10310
rect 2169 10299 2477 10308
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2608 2446 2636 12582
rect 2976 12238 3004 12718
rect 3252 12646 3280 13738
rect 3388 13084 3696 13093
rect 3388 13082 3394 13084
rect 3450 13082 3474 13084
rect 3530 13082 3554 13084
rect 3610 13082 3634 13084
rect 3690 13082 3696 13084
rect 3450 13030 3452 13082
rect 3632 13030 3634 13082
rect 3388 13028 3394 13030
rect 3450 13028 3474 13030
rect 3530 13028 3554 13030
rect 3610 13028 3634 13030
rect 3690 13028 3696 13030
rect 3388 13019 3696 13028
rect 3896 12850 3924 14758
rect 4080 14618 4108 15302
rect 4172 15162 4200 15422
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 5736 15042 5764 15370
rect 5826 15260 6134 15269
rect 5826 15258 5832 15260
rect 5888 15258 5912 15260
rect 5968 15258 5992 15260
rect 6048 15258 6072 15260
rect 6128 15258 6134 15260
rect 5888 15206 5890 15258
rect 6070 15206 6072 15258
rect 5826 15204 5832 15206
rect 5888 15204 5912 15206
rect 5968 15204 5992 15206
rect 6048 15204 6072 15206
rect 6128 15204 6134 15206
rect 5826 15195 6134 15204
rect 6196 15162 6224 15370
rect 6656 15162 6684 15438
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 5736 15026 5856 15042
rect 5540 15020 5592 15026
rect 5736 15020 5868 15026
rect 5736 15014 5816 15020
rect 5592 14980 5672 15008
rect 5540 14962 5592 14968
rect 4344 14952 4396 14958
rect 5644 14940 5672 14980
rect 5816 14962 5868 14968
rect 5644 14912 5764 14940
rect 4344 14894 4396 14900
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13938 4016 14350
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4172 13870 4200 14282
rect 4356 14278 4384 14894
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 4607 14716 4915 14725
rect 4607 14714 4613 14716
rect 4669 14714 4693 14716
rect 4749 14714 4773 14716
rect 4829 14714 4853 14716
rect 4909 14714 4915 14716
rect 4669 14662 4671 14714
rect 4851 14662 4853 14714
rect 4607 14660 4613 14662
rect 4669 14660 4693 14662
rect 4749 14660 4773 14662
rect 4829 14660 4853 14662
rect 4909 14660 4915 14662
rect 4607 14651 4915 14660
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 13938 4384 14214
rect 4448 14074 4476 14350
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13326 4200 13806
rect 4448 13394 4476 14010
rect 4540 13938 4568 14418
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 13938 4844 14282
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14074 5580 14214
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5644 13938 5672 14758
rect 5736 14618 5764 14912
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 14414 5764 14554
rect 5724 14408 5776 14414
rect 5722 14376 5724 14385
rect 5776 14376 5778 14385
rect 5722 14311 5778 14320
rect 5828 14278 5856 14962
rect 6196 14482 6224 15098
rect 6932 14958 6960 15302
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 6748 14226 6776 14350
rect 6932 14226 6960 14894
rect 7045 14716 7353 14725
rect 7045 14714 7051 14716
rect 7107 14714 7131 14716
rect 7187 14714 7211 14716
rect 7267 14714 7291 14716
rect 7347 14714 7353 14716
rect 7107 14662 7109 14714
rect 7289 14662 7291 14714
rect 7045 14660 7051 14662
rect 7107 14660 7131 14662
rect 7187 14660 7211 14662
rect 7267 14660 7291 14662
rect 7347 14660 7353 14662
rect 7045 14651 7353 14660
rect 7668 14550 7696 15370
rect 8264 15260 8572 15269
rect 8264 15258 8270 15260
rect 8326 15258 8350 15260
rect 8406 15258 8430 15260
rect 8486 15258 8510 15260
rect 8566 15258 8572 15260
rect 8326 15206 8328 15258
rect 8508 15206 8510 15258
rect 8264 15204 8270 15206
rect 8326 15204 8350 15206
rect 8406 15204 8430 15206
rect 8486 15204 8510 15206
rect 8566 15204 8572 15206
rect 8264 15195 8572 15204
rect 8680 15162 8708 15506
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7102 14376 7158 14385
rect 7102 14311 7104 14320
rect 7156 14311 7158 14320
rect 7104 14282 7156 14288
rect 6748 14198 6960 14226
rect 5826 14172 6134 14181
rect 5826 14170 5832 14172
rect 5888 14170 5912 14172
rect 5968 14170 5992 14172
rect 6048 14170 6072 14172
rect 6128 14170 6134 14172
rect 5888 14118 5890 14170
rect 6070 14118 6072 14170
rect 5826 14116 5832 14118
rect 5888 14116 5912 14118
rect 5968 14116 5992 14118
rect 6048 14116 6072 14118
rect 6128 14116 6134 14118
rect 5826 14107 6134 14116
rect 6840 14074 6868 14198
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 2514 3096 12038
rect 3388 11996 3696 12005
rect 3388 11994 3394 11996
rect 3450 11994 3474 11996
rect 3530 11994 3554 11996
rect 3610 11994 3634 11996
rect 3690 11994 3696 11996
rect 3450 11942 3452 11994
rect 3632 11942 3634 11994
rect 3388 11940 3394 11942
rect 3450 11940 3474 11942
rect 3530 11940 3554 11942
rect 3610 11940 3634 11942
rect 3690 11940 3696 11942
rect 3388 11931 3696 11940
rect 4080 11762 4108 13126
rect 4172 12918 4200 13262
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4448 12850 4476 13330
rect 4540 13326 4568 13738
rect 4607 13628 4915 13637
rect 4607 13626 4613 13628
rect 4669 13626 4693 13628
rect 4749 13626 4773 13628
rect 4829 13626 4853 13628
rect 4909 13626 4915 13628
rect 4669 13574 4671 13626
rect 4851 13574 4853 13626
rect 4607 13572 4613 13574
rect 4669 13572 4693 13574
rect 4749 13572 4773 13574
rect 4829 13572 4853 13574
rect 4909 13572 4915 13574
rect 4607 13563 4915 13572
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 11898 4200 12582
rect 4540 12238 4568 13262
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4724 12850 4752 13194
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4607 12540 4915 12549
rect 4607 12538 4613 12540
rect 4669 12538 4693 12540
rect 4749 12538 4773 12540
rect 4829 12538 4853 12540
rect 4909 12538 4915 12540
rect 4669 12486 4671 12538
rect 4851 12486 4853 12538
rect 4607 12484 4613 12486
rect 4669 12484 4693 12486
rect 4749 12484 4773 12486
rect 4829 12484 4853 12486
rect 4909 12484 4915 12486
rect 4607 12475 4915 12484
rect 5000 12238 5028 13262
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3388 10908 3696 10917
rect 3388 10906 3394 10908
rect 3450 10906 3474 10908
rect 3530 10906 3554 10908
rect 3610 10906 3634 10908
rect 3690 10906 3696 10908
rect 3450 10854 3452 10906
rect 3632 10854 3634 10906
rect 3388 10852 3394 10854
rect 3450 10852 3474 10854
rect 3530 10852 3554 10854
rect 3610 10852 3634 10854
rect 3690 10852 3696 10854
rect 3388 10843 3696 10852
rect 4080 10810 4108 11698
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4172 10470 4200 11834
rect 4540 11762 4568 12038
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4264 10130 4292 11494
rect 4448 11098 4476 11494
rect 4356 11070 4476 11098
rect 4356 11014 4384 11070
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10742 4384 10950
rect 4540 10810 4568 11698
rect 4607 11452 4915 11461
rect 4607 11450 4613 11452
rect 4669 11450 4693 11452
rect 4749 11450 4773 11452
rect 4829 11450 4853 11452
rect 4909 11450 4915 11452
rect 4669 11398 4671 11450
rect 4851 11398 4853 11450
rect 4607 11396 4613 11398
rect 4669 11396 4693 11398
rect 4749 11396 4773 11398
rect 4829 11396 4853 11398
rect 4909 11396 4915 11398
rect 4607 11387 4915 11396
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4356 10062 4384 10406
rect 4607 10364 4915 10373
rect 4607 10362 4613 10364
rect 4669 10362 4693 10364
rect 4749 10362 4773 10364
rect 4829 10362 4853 10364
rect 4909 10362 4915 10364
rect 4669 10310 4671 10362
rect 4851 10310 4853 10362
rect 4607 10308 4613 10310
rect 4669 10308 4693 10310
rect 4749 10308 4773 10310
rect 4829 10308 4853 10310
rect 4909 10308 4915 10310
rect 4607 10299 4915 10308
rect 5000 10266 5028 11222
rect 5092 11218 5120 13126
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 11830 5212 12582
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5184 11286 5212 11766
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5092 10606 5120 11154
rect 5172 11144 5224 11150
rect 5276 11098 5304 13806
rect 5644 13394 5672 13874
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5644 12918 5672 13330
rect 6472 13326 6500 13738
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 5826 13084 6134 13093
rect 5826 13082 5832 13084
rect 5888 13082 5912 13084
rect 5968 13082 5992 13084
rect 6048 13082 6072 13084
rect 6128 13082 6134 13084
rect 5888 13030 5890 13082
rect 6070 13030 6072 13082
rect 5826 13028 5832 13030
rect 5888 13028 5912 13030
rect 5968 13028 5992 13030
rect 6048 13028 6072 13030
rect 6128 13028 6134 13030
rect 5826 13019 6134 13028
rect 6472 12986 6500 13262
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 6472 12782 6500 12922
rect 6656 12918 6684 13874
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 12918 6776 13806
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 5368 11354 5396 12582
rect 5826 11996 6134 12005
rect 5826 11994 5832 11996
rect 5888 11994 5912 11996
rect 5968 11994 5992 11996
rect 6048 11994 6072 11996
rect 6128 11994 6134 11996
rect 5888 11942 5890 11994
rect 6070 11942 6072 11994
rect 5826 11940 5832 11942
rect 5888 11940 5912 11942
rect 5968 11940 5992 11942
rect 6048 11940 6072 11942
rect 6128 11940 6134 11942
rect 5826 11931 6134 11940
rect 6748 11762 6776 12582
rect 6932 11898 6960 14010
rect 7116 13938 7144 14282
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7208 13870 7236 14214
rect 7668 14006 7696 14486
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7045 13628 7353 13637
rect 7045 13626 7051 13628
rect 7107 13626 7131 13628
rect 7187 13626 7211 13628
rect 7267 13626 7291 13628
rect 7347 13626 7353 13628
rect 7107 13574 7109 13626
rect 7289 13574 7291 13626
rect 7045 13572 7051 13574
rect 7107 13572 7131 13574
rect 7187 13572 7211 13574
rect 7267 13572 7291 13574
rect 7347 13572 7353 13574
rect 7045 13563 7353 13572
rect 7484 12850 7512 13874
rect 7668 13462 7696 13942
rect 7760 13530 7788 14350
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7668 12918 7696 13398
rect 7852 13394 7880 14214
rect 7944 14074 7972 14350
rect 8128 14346 8156 14894
rect 9416 14618 9444 15506
rect 10702 15260 11010 15269
rect 10702 15258 10708 15260
rect 10764 15258 10788 15260
rect 10844 15258 10868 15260
rect 10924 15258 10948 15260
rect 11004 15258 11010 15260
rect 10764 15206 10766 15258
rect 10946 15206 10948 15258
rect 10702 15204 10708 15206
rect 10764 15204 10788 15206
rect 10844 15204 10868 15206
rect 10924 15204 10948 15206
rect 11004 15204 11010 15206
rect 10702 15195 11010 15204
rect 11072 15026 11100 17200
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 9483 14716 9791 14725
rect 9483 14714 9489 14716
rect 9545 14714 9569 14716
rect 9625 14714 9649 14716
rect 9705 14714 9729 14716
rect 9785 14714 9791 14716
rect 9545 14662 9547 14714
rect 9727 14662 9729 14714
rect 9483 14660 9489 14662
rect 9545 14660 9569 14662
rect 9625 14660 9649 14662
rect 9705 14660 9729 14662
rect 9785 14660 9791 14662
rect 9483 14651 9791 14660
rect 10336 14618 10364 14962
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7944 13818 7972 14010
rect 8128 14006 8156 14282
rect 8264 14172 8572 14181
rect 8264 14170 8270 14172
rect 8326 14170 8350 14172
rect 8406 14170 8430 14172
rect 8486 14170 8510 14172
rect 8566 14170 8572 14172
rect 8326 14118 8328 14170
rect 8508 14118 8510 14170
rect 8264 14116 8270 14118
rect 8326 14116 8350 14118
rect 8406 14116 8430 14118
rect 8486 14116 8510 14118
rect 8566 14116 8572 14118
rect 8264 14107 8572 14116
rect 10702 14172 11010 14181
rect 10702 14170 10708 14172
rect 10764 14170 10788 14172
rect 10844 14170 10868 14172
rect 10924 14170 10948 14172
rect 11004 14170 11010 14172
rect 10764 14118 10766 14170
rect 10946 14118 10948 14170
rect 10702 14116 10708 14118
rect 10764 14116 10788 14118
rect 10844 14116 10868 14118
rect 10924 14116 10948 14118
rect 11004 14116 11010 14118
rect 10702 14107 11010 14116
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7944 13790 8064 13818
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7944 13258 7972 13670
rect 8036 13326 8064 13790
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7045 12540 7353 12549
rect 7045 12538 7051 12540
rect 7107 12538 7131 12540
rect 7187 12538 7211 12540
rect 7267 12538 7291 12540
rect 7347 12538 7353 12540
rect 7107 12486 7109 12538
rect 7289 12486 7291 12538
rect 7045 12484 7051 12486
rect 7107 12484 7131 12486
rect 7187 12484 7211 12486
rect 7267 12484 7291 12486
rect 7347 12484 7353 12486
rect 7045 12475 7353 12484
rect 7668 12238 7696 12582
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5368 11150 5396 11290
rect 5460 11234 5488 11698
rect 5460 11206 5580 11234
rect 5552 11150 5580 11206
rect 5224 11092 5304 11098
rect 5172 11086 5304 11092
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5184 11070 5304 11086
rect 5184 10742 5212 11070
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5368 10674 5396 11086
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 4264 2446 4292 9862
rect 4908 9586 4936 9930
rect 5000 9722 5028 10202
rect 5092 9994 5120 10406
rect 5736 10062 5764 11018
rect 5826 10908 6134 10917
rect 5826 10906 5832 10908
rect 5888 10906 5912 10908
rect 5968 10906 5992 10908
rect 6048 10906 6072 10908
rect 6128 10906 6134 10908
rect 5888 10854 5890 10906
rect 6070 10854 6072 10906
rect 5826 10852 5832 10854
rect 5888 10852 5912 10854
rect 5968 10852 5992 10854
rect 6048 10852 6072 10854
rect 6128 10852 6134 10854
rect 5826 10843 6134 10852
rect 6748 10538 6776 11698
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11354 6868 11630
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10742 6868 11290
rect 6932 10810 6960 11834
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7045 11452 7353 11461
rect 7045 11450 7051 11452
rect 7107 11450 7131 11452
rect 7187 11450 7211 11452
rect 7267 11450 7291 11452
rect 7347 11450 7353 11452
rect 7107 11398 7109 11450
rect 7289 11398 7291 11450
rect 7045 11396 7051 11398
rect 7107 11396 7131 11398
rect 7187 11396 7211 11398
rect 7267 11396 7291 11398
rect 7347 11396 7353 11398
rect 7045 11387 7353 11396
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 6656 9994 6684 10406
rect 6748 10010 6776 10474
rect 6840 10130 6868 10678
rect 7484 10674 7512 10950
rect 7576 10674 7604 11494
rect 7668 11234 7696 12174
rect 7668 11206 7788 11234
rect 7760 11150 7788 11206
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10538 7604 10610
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7045 10364 7353 10373
rect 7045 10362 7051 10364
rect 7107 10362 7131 10364
rect 7187 10362 7211 10364
rect 7267 10362 7291 10364
rect 7347 10362 7353 10364
rect 7107 10310 7109 10362
rect 7289 10310 7291 10362
rect 7045 10308 7051 10310
rect 7107 10308 7131 10310
rect 7187 10308 7211 10310
rect 7267 10308 7291 10310
rect 7347 10308 7353 10310
rect 7045 10299 7353 10308
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 10010 6960 10066
rect 7668 10062 7696 10746
rect 7852 10674 7880 13126
rect 7944 12850 7972 13194
rect 8128 12850 8156 13942
rect 9483 13628 9791 13637
rect 9483 13626 9489 13628
rect 9545 13626 9569 13628
rect 9625 13626 9649 13628
rect 9705 13626 9729 13628
rect 9785 13626 9791 13628
rect 9545 13574 9547 13626
rect 9727 13574 9729 13626
rect 9483 13572 9489 13574
rect 9545 13572 9569 13574
rect 9625 13572 9649 13574
rect 9705 13572 9729 13574
rect 9785 13572 9791 13574
rect 9483 13563 9791 13572
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8264 13084 8572 13093
rect 8264 13082 8270 13084
rect 8326 13082 8350 13084
rect 8406 13082 8430 13084
rect 8486 13082 8510 13084
rect 8566 13082 8572 13084
rect 8326 13030 8328 13082
rect 8508 13030 8510 13082
rect 8264 13028 8270 13030
rect 8326 13028 8350 13030
rect 8406 13028 8430 13030
rect 8486 13028 8510 13030
rect 8566 13028 8572 13030
rect 8264 13019 8572 13028
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12238 8064 12582
rect 8680 12238 8708 13126
rect 10702 13084 11010 13093
rect 10702 13082 10708 13084
rect 10764 13082 10788 13084
rect 10844 13082 10868 13084
rect 10924 13082 10948 13084
rect 11004 13082 11010 13084
rect 10764 13030 10766 13082
rect 10946 13030 10948 13082
rect 10702 13028 10708 13030
rect 10764 13028 10788 13030
rect 10844 13028 10868 13030
rect 10924 13028 10948 13030
rect 11004 13028 11010 13030
rect 10702 13019 11010 13028
rect 9483 12540 9791 12549
rect 9483 12538 9489 12540
rect 9545 12538 9569 12540
rect 9625 12538 9649 12540
rect 9705 12538 9729 12540
rect 9785 12538 9791 12540
rect 9545 12486 9547 12538
rect 9727 12486 9729 12538
rect 9483 12484 9489 12486
rect 9545 12484 9569 12486
rect 9625 12484 9649 12486
rect 9705 12484 9729 12486
rect 9785 12484 9791 12486
rect 9483 12475 9791 12484
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8264 11996 8572 12005
rect 8264 11994 8270 11996
rect 8326 11994 8350 11996
rect 8406 11994 8430 11996
rect 8486 11994 8510 11996
rect 8566 11994 8572 11996
rect 8326 11942 8328 11994
rect 8508 11942 8510 11994
rect 8264 11940 8270 11942
rect 8326 11940 8350 11942
rect 8406 11940 8430 11942
rect 8486 11940 8510 11942
rect 8566 11940 8572 11942
rect 8264 11931 8572 11940
rect 8264 10908 8572 10917
rect 8264 10906 8270 10908
rect 8326 10906 8350 10908
rect 8406 10906 8430 10908
rect 8486 10906 8510 10908
rect 8566 10906 8572 10908
rect 8326 10854 8328 10906
rect 8508 10854 8510 10906
rect 8264 10852 8270 10854
rect 8326 10852 8350 10854
rect 8406 10852 8430 10854
rect 8486 10852 8510 10854
rect 8566 10852 8572 10854
rect 8264 10843 8572 10852
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8220 10062 8248 10406
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 6644 9988 6696 9994
rect 6748 9982 6960 10010
rect 7656 10056 7708 10062
rect 8208 10056 8260 10062
rect 7656 9998 7708 10004
rect 8128 10004 8208 10010
rect 8128 9998 8260 10004
rect 8128 9982 8248 9998
rect 6644 9930 6696 9936
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 5092 9654 5120 9930
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5276 9586 5304 9862
rect 5736 9722 5764 9862
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 5000 8974 5028 9318
rect 5276 8974 5304 9522
rect 5736 9450 5764 9658
rect 7024 9586 7052 9862
rect 8128 9586 8156 9982
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 8974 5856 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7484 9042 7512 9454
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 5276 2446 5304 8774
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 6748 2446 6776 8978
rect 8588 8974 8616 9590
rect 8680 9042 8708 9862
rect 8772 9722 8800 10406
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8864 9654 8892 12310
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7944 2446 7972 8774
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8772 8498 8800 9318
rect 8864 8566 8892 9590
rect 9048 9586 9076 12106
rect 10702 11996 11010 12005
rect 10702 11994 10708 11996
rect 10764 11994 10788 11996
rect 10844 11994 10868 11996
rect 10924 11994 10948 11996
rect 11004 11994 11010 11996
rect 10764 11942 10766 11994
rect 10946 11942 10948 11994
rect 10702 11940 10708 11942
rect 10764 11940 10788 11942
rect 10844 11940 10868 11942
rect 10924 11940 10948 11942
rect 11004 11940 11010 11942
rect 10702 11931 11010 11940
rect 9483 11452 9791 11461
rect 9483 11450 9489 11452
rect 9545 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9791 11452
rect 9545 11398 9547 11450
rect 9727 11398 9729 11450
rect 9483 11396 9489 11398
rect 9545 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9791 11398
rect 9483 11387 9791 11396
rect 10702 10908 11010 10917
rect 10702 10906 10708 10908
rect 10764 10906 10788 10908
rect 10844 10906 10868 10908
rect 10924 10906 10948 10908
rect 11004 10906 11010 10908
rect 10764 10854 10766 10906
rect 10946 10854 10948 10906
rect 10702 10852 10708 10854
rect 10764 10852 10788 10854
rect 10844 10852 10868 10854
rect 10924 10852 10948 10854
rect 11004 10852 11010 10854
rect 10702 10843 11010 10852
rect 9483 10364 9791 10373
rect 9483 10362 9489 10364
rect 9545 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9791 10364
rect 9545 10310 9547 10362
rect 9727 10310 9729 10362
rect 9483 10308 9489 10310
rect 9545 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9791 10310
rect 9483 10299 9791 10308
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9968 2446 9996 8298
rect 10060 3058 10088 9318
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 756 2304 808 2310
rect 756 2246 808 2252
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 768 800 796 2246
rect 2240 800 2268 2246
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3804 1170 3832 2246
rect 3712 1142 3832 1170
rect 3712 800 3740 1142
rect 5184 800 5212 2246
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6656 800 6684 2246
rect 8128 800 8156 2246
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 9600 800 9628 2246
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 11072 800 11100 2790
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
<< via2 >>
rect 2175 15802 2231 15804
rect 2255 15802 2311 15804
rect 2335 15802 2391 15804
rect 2415 15802 2471 15804
rect 2175 15750 2221 15802
rect 2221 15750 2231 15802
rect 2255 15750 2285 15802
rect 2285 15750 2297 15802
rect 2297 15750 2311 15802
rect 2335 15750 2349 15802
rect 2349 15750 2361 15802
rect 2361 15750 2391 15802
rect 2415 15750 2425 15802
rect 2425 15750 2471 15802
rect 2175 15748 2231 15750
rect 2255 15748 2311 15750
rect 2335 15748 2391 15750
rect 2415 15748 2471 15750
rect 4613 15802 4669 15804
rect 4693 15802 4749 15804
rect 4773 15802 4829 15804
rect 4853 15802 4909 15804
rect 4613 15750 4659 15802
rect 4659 15750 4669 15802
rect 4693 15750 4723 15802
rect 4723 15750 4735 15802
rect 4735 15750 4749 15802
rect 4773 15750 4787 15802
rect 4787 15750 4799 15802
rect 4799 15750 4829 15802
rect 4853 15750 4863 15802
rect 4863 15750 4909 15802
rect 4613 15748 4669 15750
rect 4693 15748 4749 15750
rect 4773 15748 4829 15750
rect 4853 15748 4909 15750
rect 7051 15802 7107 15804
rect 7131 15802 7187 15804
rect 7211 15802 7267 15804
rect 7291 15802 7347 15804
rect 7051 15750 7097 15802
rect 7097 15750 7107 15802
rect 7131 15750 7161 15802
rect 7161 15750 7173 15802
rect 7173 15750 7187 15802
rect 7211 15750 7225 15802
rect 7225 15750 7237 15802
rect 7237 15750 7267 15802
rect 7291 15750 7301 15802
rect 7301 15750 7347 15802
rect 7051 15748 7107 15750
rect 7131 15748 7187 15750
rect 7211 15748 7267 15750
rect 7291 15748 7347 15750
rect 9489 15802 9545 15804
rect 9569 15802 9625 15804
rect 9649 15802 9705 15804
rect 9729 15802 9785 15804
rect 9489 15750 9535 15802
rect 9535 15750 9545 15802
rect 9569 15750 9599 15802
rect 9599 15750 9611 15802
rect 9611 15750 9625 15802
rect 9649 15750 9663 15802
rect 9663 15750 9675 15802
rect 9675 15750 9705 15802
rect 9729 15750 9739 15802
rect 9739 15750 9785 15802
rect 9489 15748 9545 15750
rect 9569 15748 9625 15750
rect 9649 15748 9705 15750
rect 9729 15748 9785 15750
rect 3394 15258 3450 15260
rect 3474 15258 3530 15260
rect 3554 15258 3610 15260
rect 3634 15258 3690 15260
rect 3394 15206 3440 15258
rect 3440 15206 3450 15258
rect 3474 15206 3504 15258
rect 3504 15206 3516 15258
rect 3516 15206 3530 15258
rect 3554 15206 3568 15258
rect 3568 15206 3580 15258
rect 3580 15206 3610 15258
rect 3634 15206 3644 15258
rect 3644 15206 3690 15258
rect 3394 15204 3450 15206
rect 3474 15204 3530 15206
rect 3554 15204 3610 15206
rect 3634 15204 3690 15206
rect 2175 14714 2231 14716
rect 2255 14714 2311 14716
rect 2335 14714 2391 14716
rect 2415 14714 2471 14716
rect 2175 14662 2221 14714
rect 2221 14662 2231 14714
rect 2255 14662 2285 14714
rect 2285 14662 2297 14714
rect 2297 14662 2311 14714
rect 2335 14662 2349 14714
rect 2349 14662 2361 14714
rect 2361 14662 2391 14714
rect 2415 14662 2425 14714
rect 2425 14662 2471 14714
rect 2175 14660 2231 14662
rect 2255 14660 2311 14662
rect 2335 14660 2391 14662
rect 2415 14660 2471 14662
rect 2175 13626 2231 13628
rect 2255 13626 2311 13628
rect 2335 13626 2391 13628
rect 2415 13626 2471 13628
rect 2175 13574 2221 13626
rect 2221 13574 2231 13626
rect 2255 13574 2285 13626
rect 2285 13574 2297 13626
rect 2297 13574 2311 13626
rect 2335 13574 2349 13626
rect 2349 13574 2361 13626
rect 2361 13574 2391 13626
rect 2415 13574 2425 13626
rect 2425 13574 2471 13626
rect 2175 13572 2231 13574
rect 2255 13572 2311 13574
rect 2335 13572 2391 13574
rect 2415 13572 2471 13574
rect 3394 14170 3450 14172
rect 3474 14170 3530 14172
rect 3554 14170 3610 14172
rect 3634 14170 3690 14172
rect 3394 14118 3440 14170
rect 3440 14118 3450 14170
rect 3474 14118 3504 14170
rect 3504 14118 3516 14170
rect 3516 14118 3530 14170
rect 3554 14118 3568 14170
rect 3568 14118 3580 14170
rect 3580 14118 3610 14170
rect 3634 14118 3644 14170
rect 3644 14118 3690 14170
rect 3394 14116 3450 14118
rect 3474 14116 3530 14118
rect 3554 14116 3610 14118
rect 3634 14116 3690 14118
rect 2175 12538 2231 12540
rect 2255 12538 2311 12540
rect 2335 12538 2391 12540
rect 2415 12538 2471 12540
rect 2175 12486 2221 12538
rect 2221 12486 2231 12538
rect 2255 12486 2285 12538
rect 2285 12486 2297 12538
rect 2297 12486 2311 12538
rect 2335 12486 2349 12538
rect 2349 12486 2361 12538
rect 2361 12486 2391 12538
rect 2415 12486 2425 12538
rect 2425 12486 2471 12538
rect 2175 12484 2231 12486
rect 2255 12484 2311 12486
rect 2335 12484 2391 12486
rect 2415 12484 2471 12486
rect 2175 11450 2231 11452
rect 2255 11450 2311 11452
rect 2335 11450 2391 11452
rect 2415 11450 2471 11452
rect 2175 11398 2221 11450
rect 2221 11398 2231 11450
rect 2255 11398 2285 11450
rect 2285 11398 2297 11450
rect 2297 11398 2311 11450
rect 2335 11398 2349 11450
rect 2349 11398 2361 11450
rect 2361 11398 2391 11450
rect 2415 11398 2425 11450
rect 2425 11398 2471 11450
rect 2175 11396 2231 11398
rect 2255 11396 2311 11398
rect 2335 11396 2391 11398
rect 2415 11396 2471 11398
rect 2175 10362 2231 10364
rect 2255 10362 2311 10364
rect 2335 10362 2391 10364
rect 2415 10362 2471 10364
rect 2175 10310 2221 10362
rect 2221 10310 2231 10362
rect 2255 10310 2285 10362
rect 2285 10310 2297 10362
rect 2297 10310 2311 10362
rect 2335 10310 2349 10362
rect 2349 10310 2361 10362
rect 2361 10310 2391 10362
rect 2415 10310 2425 10362
rect 2425 10310 2471 10362
rect 2175 10308 2231 10310
rect 2255 10308 2311 10310
rect 2335 10308 2391 10310
rect 2415 10308 2471 10310
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 13082 3450 13084
rect 3474 13082 3530 13084
rect 3554 13082 3610 13084
rect 3634 13082 3690 13084
rect 3394 13030 3440 13082
rect 3440 13030 3450 13082
rect 3474 13030 3504 13082
rect 3504 13030 3516 13082
rect 3516 13030 3530 13082
rect 3554 13030 3568 13082
rect 3568 13030 3580 13082
rect 3580 13030 3610 13082
rect 3634 13030 3644 13082
rect 3644 13030 3690 13082
rect 3394 13028 3450 13030
rect 3474 13028 3530 13030
rect 3554 13028 3610 13030
rect 3634 13028 3690 13030
rect 5832 15258 5888 15260
rect 5912 15258 5968 15260
rect 5992 15258 6048 15260
rect 6072 15258 6128 15260
rect 5832 15206 5878 15258
rect 5878 15206 5888 15258
rect 5912 15206 5942 15258
rect 5942 15206 5954 15258
rect 5954 15206 5968 15258
rect 5992 15206 6006 15258
rect 6006 15206 6018 15258
rect 6018 15206 6048 15258
rect 6072 15206 6082 15258
rect 6082 15206 6128 15258
rect 5832 15204 5888 15206
rect 5912 15204 5968 15206
rect 5992 15204 6048 15206
rect 6072 15204 6128 15206
rect 4613 14714 4669 14716
rect 4693 14714 4749 14716
rect 4773 14714 4829 14716
rect 4853 14714 4909 14716
rect 4613 14662 4659 14714
rect 4659 14662 4669 14714
rect 4693 14662 4723 14714
rect 4723 14662 4735 14714
rect 4735 14662 4749 14714
rect 4773 14662 4787 14714
rect 4787 14662 4799 14714
rect 4799 14662 4829 14714
rect 4853 14662 4863 14714
rect 4863 14662 4909 14714
rect 4613 14660 4669 14662
rect 4693 14660 4749 14662
rect 4773 14660 4829 14662
rect 4853 14660 4909 14662
rect 5722 14356 5724 14376
rect 5724 14356 5776 14376
rect 5776 14356 5778 14376
rect 5722 14320 5778 14356
rect 7051 14714 7107 14716
rect 7131 14714 7187 14716
rect 7211 14714 7267 14716
rect 7291 14714 7347 14716
rect 7051 14662 7097 14714
rect 7097 14662 7107 14714
rect 7131 14662 7161 14714
rect 7161 14662 7173 14714
rect 7173 14662 7187 14714
rect 7211 14662 7225 14714
rect 7225 14662 7237 14714
rect 7237 14662 7267 14714
rect 7291 14662 7301 14714
rect 7301 14662 7347 14714
rect 7051 14660 7107 14662
rect 7131 14660 7187 14662
rect 7211 14660 7267 14662
rect 7291 14660 7347 14662
rect 8270 15258 8326 15260
rect 8350 15258 8406 15260
rect 8430 15258 8486 15260
rect 8510 15258 8566 15260
rect 8270 15206 8316 15258
rect 8316 15206 8326 15258
rect 8350 15206 8380 15258
rect 8380 15206 8392 15258
rect 8392 15206 8406 15258
rect 8430 15206 8444 15258
rect 8444 15206 8456 15258
rect 8456 15206 8486 15258
rect 8510 15206 8520 15258
rect 8520 15206 8566 15258
rect 8270 15204 8326 15206
rect 8350 15204 8406 15206
rect 8430 15204 8486 15206
rect 8510 15204 8566 15206
rect 7102 14340 7158 14376
rect 7102 14320 7104 14340
rect 7104 14320 7156 14340
rect 7156 14320 7158 14340
rect 5832 14170 5888 14172
rect 5912 14170 5968 14172
rect 5992 14170 6048 14172
rect 6072 14170 6128 14172
rect 5832 14118 5878 14170
rect 5878 14118 5888 14170
rect 5912 14118 5942 14170
rect 5942 14118 5954 14170
rect 5954 14118 5968 14170
rect 5992 14118 6006 14170
rect 6006 14118 6018 14170
rect 6018 14118 6048 14170
rect 6072 14118 6082 14170
rect 6082 14118 6128 14170
rect 5832 14116 5888 14118
rect 5912 14116 5968 14118
rect 5992 14116 6048 14118
rect 6072 14116 6128 14118
rect 3394 11994 3450 11996
rect 3474 11994 3530 11996
rect 3554 11994 3610 11996
rect 3634 11994 3690 11996
rect 3394 11942 3440 11994
rect 3440 11942 3450 11994
rect 3474 11942 3504 11994
rect 3504 11942 3516 11994
rect 3516 11942 3530 11994
rect 3554 11942 3568 11994
rect 3568 11942 3580 11994
rect 3580 11942 3610 11994
rect 3634 11942 3644 11994
rect 3644 11942 3690 11994
rect 3394 11940 3450 11942
rect 3474 11940 3530 11942
rect 3554 11940 3610 11942
rect 3634 11940 3690 11942
rect 4613 13626 4669 13628
rect 4693 13626 4749 13628
rect 4773 13626 4829 13628
rect 4853 13626 4909 13628
rect 4613 13574 4659 13626
rect 4659 13574 4669 13626
rect 4693 13574 4723 13626
rect 4723 13574 4735 13626
rect 4735 13574 4749 13626
rect 4773 13574 4787 13626
rect 4787 13574 4799 13626
rect 4799 13574 4829 13626
rect 4853 13574 4863 13626
rect 4863 13574 4909 13626
rect 4613 13572 4669 13574
rect 4693 13572 4749 13574
rect 4773 13572 4829 13574
rect 4853 13572 4909 13574
rect 4613 12538 4669 12540
rect 4693 12538 4749 12540
rect 4773 12538 4829 12540
rect 4853 12538 4909 12540
rect 4613 12486 4659 12538
rect 4659 12486 4669 12538
rect 4693 12486 4723 12538
rect 4723 12486 4735 12538
rect 4735 12486 4749 12538
rect 4773 12486 4787 12538
rect 4787 12486 4799 12538
rect 4799 12486 4829 12538
rect 4853 12486 4863 12538
rect 4863 12486 4909 12538
rect 4613 12484 4669 12486
rect 4693 12484 4749 12486
rect 4773 12484 4829 12486
rect 4853 12484 4909 12486
rect 3394 10906 3450 10908
rect 3474 10906 3530 10908
rect 3554 10906 3610 10908
rect 3634 10906 3690 10908
rect 3394 10854 3440 10906
rect 3440 10854 3450 10906
rect 3474 10854 3504 10906
rect 3504 10854 3516 10906
rect 3516 10854 3530 10906
rect 3554 10854 3568 10906
rect 3568 10854 3580 10906
rect 3580 10854 3610 10906
rect 3634 10854 3644 10906
rect 3644 10854 3690 10906
rect 3394 10852 3450 10854
rect 3474 10852 3530 10854
rect 3554 10852 3610 10854
rect 3634 10852 3690 10854
rect 4613 11450 4669 11452
rect 4693 11450 4749 11452
rect 4773 11450 4829 11452
rect 4853 11450 4909 11452
rect 4613 11398 4659 11450
rect 4659 11398 4669 11450
rect 4693 11398 4723 11450
rect 4723 11398 4735 11450
rect 4735 11398 4749 11450
rect 4773 11398 4787 11450
rect 4787 11398 4799 11450
rect 4799 11398 4829 11450
rect 4853 11398 4863 11450
rect 4863 11398 4909 11450
rect 4613 11396 4669 11398
rect 4693 11396 4749 11398
rect 4773 11396 4829 11398
rect 4853 11396 4909 11398
rect 4613 10362 4669 10364
rect 4693 10362 4749 10364
rect 4773 10362 4829 10364
rect 4853 10362 4909 10364
rect 4613 10310 4659 10362
rect 4659 10310 4669 10362
rect 4693 10310 4723 10362
rect 4723 10310 4735 10362
rect 4735 10310 4749 10362
rect 4773 10310 4787 10362
rect 4787 10310 4799 10362
rect 4799 10310 4829 10362
rect 4853 10310 4863 10362
rect 4863 10310 4909 10362
rect 4613 10308 4669 10310
rect 4693 10308 4749 10310
rect 4773 10308 4829 10310
rect 4853 10308 4909 10310
rect 5832 13082 5888 13084
rect 5912 13082 5968 13084
rect 5992 13082 6048 13084
rect 6072 13082 6128 13084
rect 5832 13030 5878 13082
rect 5878 13030 5888 13082
rect 5912 13030 5942 13082
rect 5942 13030 5954 13082
rect 5954 13030 5968 13082
rect 5992 13030 6006 13082
rect 6006 13030 6018 13082
rect 6018 13030 6048 13082
rect 6072 13030 6082 13082
rect 6082 13030 6128 13082
rect 5832 13028 5888 13030
rect 5912 13028 5968 13030
rect 5992 13028 6048 13030
rect 6072 13028 6128 13030
rect 5832 11994 5888 11996
rect 5912 11994 5968 11996
rect 5992 11994 6048 11996
rect 6072 11994 6128 11996
rect 5832 11942 5878 11994
rect 5878 11942 5888 11994
rect 5912 11942 5942 11994
rect 5942 11942 5954 11994
rect 5954 11942 5968 11994
rect 5992 11942 6006 11994
rect 6006 11942 6018 11994
rect 6018 11942 6048 11994
rect 6072 11942 6082 11994
rect 6082 11942 6128 11994
rect 5832 11940 5888 11942
rect 5912 11940 5968 11942
rect 5992 11940 6048 11942
rect 6072 11940 6128 11942
rect 7051 13626 7107 13628
rect 7131 13626 7187 13628
rect 7211 13626 7267 13628
rect 7291 13626 7347 13628
rect 7051 13574 7097 13626
rect 7097 13574 7107 13626
rect 7131 13574 7161 13626
rect 7161 13574 7173 13626
rect 7173 13574 7187 13626
rect 7211 13574 7225 13626
rect 7225 13574 7237 13626
rect 7237 13574 7267 13626
rect 7291 13574 7301 13626
rect 7301 13574 7347 13626
rect 7051 13572 7107 13574
rect 7131 13572 7187 13574
rect 7211 13572 7267 13574
rect 7291 13572 7347 13574
rect 10708 15258 10764 15260
rect 10788 15258 10844 15260
rect 10868 15258 10924 15260
rect 10948 15258 11004 15260
rect 10708 15206 10754 15258
rect 10754 15206 10764 15258
rect 10788 15206 10818 15258
rect 10818 15206 10830 15258
rect 10830 15206 10844 15258
rect 10868 15206 10882 15258
rect 10882 15206 10894 15258
rect 10894 15206 10924 15258
rect 10948 15206 10958 15258
rect 10958 15206 11004 15258
rect 10708 15204 10764 15206
rect 10788 15204 10844 15206
rect 10868 15204 10924 15206
rect 10948 15204 11004 15206
rect 9489 14714 9545 14716
rect 9569 14714 9625 14716
rect 9649 14714 9705 14716
rect 9729 14714 9785 14716
rect 9489 14662 9535 14714
rect 9535 14662 9545 14714
rect 9569 14662 9599 14714
rect 9599 14662 9611 14714
rect 9611 14662 9625 14714
rect 9649 14662 9663 14714
rect 9663 14662 9675 14714
rect 9675 14662 9705 14714
rect 9729 14662 9739 14714
rect 9739 14662 9785 14714
rect 9489 14660 9545 14662
rect 9569 14660 9625 14662
rect 9649 14660 9705 14662
rect 9729 14660 9785 14662
rect 8270 14170 8326 14172
rect 8350 14170 8406 14172
rect 8430 14170 8486 14172
rect 8510 14170 8566 14172
rect 8270 14118 8316 14170
rect 8316 14118 8326 14170
rect 8350 14118 8380 14170
rect 8380 14118 8392 14170
rect 8392 14118 8406 14170
rect 8430 14118 8444 14170
rect 8444 14118 8456 14170
rect 8456 14118 8486 14170
rect 8510 14118 8520 14170
rect 8520 14118 8566 14170
rect 8270 14116 8326 14118
rect 8350 14116 8406 14118
rect 8430 14116 8486 14118
rect 8510 14116 8566 14118
rect 10708 14170 10764 14172
rect 10788 14170 10844 14172
rect 10868 14170 10924 14172
rect 10948 14170 11004 14172
rect 10708 14118 10754 14170
rect 10754 14118 10764 14170
rect 10788 14118 10818 14170
rect 10818 14118 10830 14170
rect 10830 14118 10844 14170
rect 10868 14118 10882 14170
rect 10882 14118 10894 14170
rect 10894 14118 10924 14170
rect 10948 14118 10958 14170
rect 10958 14118 11004 14170
rect 10708 14116 10764 14118
rect 10788 14116 10844 14118
rect 10868 14116 10924 14118
rect 10948 14116 11004 14118
rect 7051 12538 7107 12540
rect 7131 12538 7187 12540
rect 7211 12538 7267 12540
rect 7291 12538 7347 12540
rect 7051 12486 7097 12538
rect 7097 12486 7107 12538
rect 7131 12486 7161 12538
rect 7161 12486 7173 12538
rect 7173 12486 7187 12538
rect 7211 12486 7225 12538
rect 7225 12486 7237 12538
rect 7237 12486 7267 12538
rect 7291 12486 7301 12538
rect 7301 12486 7347 12538
rect 7051 12484 7107 12486
rect 7131 12484 7187 12486
rect 7211 12484 7267 12486
rect 7291 12484 7347 12486
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 5832 10906 5888 10908
rect 5912 10906 5968 10908
rect 5992 10906 6048 10908
rect 6072 10906 6128 10908
rect 5832 10854 5878 10906
rect 5878 10854 5888 10906
rect 5912 10854 5942 10906
rect 5942 10854 5954 10906
rect 5954 10854 5968 10906
rect 5992 10854 6006 10906
rect 6006 10854 6018 10906
rect 6018 10854 6048 10906
rect 6072 10854 6082 10906
rect 6082 10854 6128 10906
rect 5832 10852 5888 10854
rect 5912 10852 5968 10854
rect 5992 10852 6048 10854
rect 6072 10852 6128 10854
rect 7051 11450 7107 11452
rect 7131 11450 7187 11452
rect 7211 11450 7267 11452
rect 7291 11450 7347 11452
rect 7051 11398 7097 11450
rect 7097 11398 7107 11450
rect 7131 11398 7161 11450
rect 7161 11398 7173 11450
rect 7173 11398 7187 11450
rect 7211 11398 7225 11450
rect 7225 11398 7237 11450
rect 7237 11398 7267 11450
rect 7291 11398 7301 11450
rect 7301 11398 7347 11450
rect 7051 11396 7107 11398
rect 7131 11396 7187 11398
rect 7211 11396 7267 11398
rect 7291 11396 7347 11398
rect 7051 10362 7107 10364
rect 7131 10362 7187 10364
rect 7211 10362 7267 10364
rect 7291 10362 7347 10364
rect 7051 10310 7097 10362
rect 7097 10310 7107 10362
rect 7131 10310 7161 10362
rect 7161 10310 7173 10362
rect 7173 10310 7187 10362
rect 7211 10310 7225 10362
rect 7225 10310 7237 10362
rect 7237 10310 7267 10362
rect 7291 10310 7301 10362
rect 7301 10310 7347 10362
rect 7051 10308 7107 10310
rect 7131 10308 7187 10310
rect 7211 10308 7267 10310
rect 7291 10308 7347 10310
rect 9489 13626 9545 13628
rect 9569 13626 9625 13628
rect 9649 13626 9705 13628
rect 9729 13626 9785 13628
rect 9489 13574 9535 13626
rect 9535 13574 9545 13626
rect 9569 13574 9599 13626
rect 9599 13574 9611 13626
rect 9611 13574 9625 13626
rect 9649 13574 9663 13626
rect 9663 13574 9675 13626
rect 9675 13574 9705 13626
rect 9729 13574 9739 13626
rect 9739 13574 9785 13626
rect 9489 13572 9545 13574
rect 9569 13572 9625 13574
rect 9649 13572 9705 13574
rect 9729 13572 9785 13574
rect 8270 13082 8326 13084
rect 8350 13082 8406 13084
rect 8430 13082 8486 13084
rect 8510 13082 8566 13084
rect 8270 13030 8316 13082
rect 8316 13030 8326 13082
rect 8350 13030 8380 13082
rect 8380 13030 8392 13082
rect 8392 13030 8406 13082
rect 8430 13030 8444 13082
rect 8444 13030 8456 13082
rect 8456 13030 8486 13082
rect 8510 13030 8520 13082
rect 8520 13030 8566 13082
rect 8270 13028 8326 13030
rect 8350 13028 8406 13030
rect 8430 13028 8486 13030
rect 8510 13028 8566 13030
rect 10708 13082 10764 13084
rect 10788 13082 10844 13084
rect 10868 13082 10924 13084
rect 10948 13082 11004 13084
rect 10708 13030 10754 13082
rect 10754 13030 10764 13082
rect 10788 13030 10818 13082
rect 10818 13030 10830 13082
rect 10830 13030 10844 13082
rect 10868 13030 10882 13082
rect 10882 13030 10894 13082
rect 10894 13030 10924 13082
rect 10948 13030 10958 13082
rect 10958 13030 11004 13082
rect 10708 13028 10764 13030
rect 10788 13028 10844 13030
rect 10868 13028 10924 13030
rect 10948 13028 11004 13030
rect 9489 12538 9545 12540
rect 9569 12538 9625 12540
rect 9649 12538 9705 12540
rect 9729 12538 9785 12540
rect 9489 12486 9535 12538
rect 9535 12486 9545 12538
rect 9569 12486 9599 12538
rect 9599 12486 9611 12538
rect 9611 12486 9625 12538
rect 9649 12486 9663 12538
rect 9663 12486 9675 12538
rect 9675 12486 9705 12538
rect 9729 12486 9739 12538
rect 9739 12486 9785 12538
rect 9489 12484 9545 12486
rect 9569 12484 9625 12486
rect 9649 12484 9705 12486
rect 9729 12484 9785 12486
rect 8270 11994 8326 11996
rect 8350 11994 8406 11996
rect 8430 11994 8486 11996
rect 8510 11994 8566 11996
rect 8270 11942 8316 11994
rect 8316 11942 8326 11994
rect 8350 11942 8380 11994
rect 8380 11942 8392 11994
rect 8392 11942 8406 11994
rect 8430 11942 8444 11994
rect 8444 11942 8456 11994
rect 8456 11942 8486 11994
rect 8510 11942 8520 11994
rect 8520 11942 8566 11994
rect 8270 11940 8326 11942
rect 8350 11940 8406 11942
rect 8430 11940 8486 11942
rect 8510 11940 8566 11942
rect 8270 10906 8326 10908
rect 8350 10906 8406 10908
rect 8430 10906 8486 10908
rect 8510 10906 8566 10908
rect 8270 10854 8316 10906
rect 8316 10854 8326 10906
rect 8350 10854 8380 10906
rect 8380 10854 8392 10906
rect 8392 10854 8406 10906
rect 8430 10854 8444 10906
rect 8444 10854 8456 10906
rect 8456 10854 8486 10906
rect 8510 10854 8520 10906
rect 8520 10854 8566 10906
rect 8270 10852 8326 10854
rect 8350 10852 8406 10854
rect 8430 10852 8486 10854
rect 8510 10852 8566 10854
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 10708 11994 10764 11996
rect 10788 11994 10844 11996
rect 10868 11994 10924 11996
rect 10948 11994 11004 11996
rect 10708 11942 10754 11994
rect 10754 11942 10764 11994
rect 10788 11942 10818 11994
rect 10818 11942 10830 11994
rect 10830 11942 10844 11994
rect 10868 11942 10882 11994
rect 10882 11942 10894 11994
rect 10894 11942 10924 11994
rect 10948 11942 10958 11994
rect 10958 11942 11004 11994
rect 10708 11940 10764 11942
rect 10788 11940 10844 11942
rect 10868 11940 10924 11942
rect 10948 11940 11004 11942
rect 9489 11450 9545 11452
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9489 11398 9535 11450
rect 9535 11398 9545 11450
rect 9569 11398 9599 11450
rect 9599 11398 9611 11450
rect 9611 11398 9625 11450
rect 9649 11398 9663 11450
rect 9663 11398 9675 11450
rect 9675 11398 9705 11450
rect 9729 11398 9739 11450
rect 9739 11398 9785 11450
rect 9489 11396 9545 11398
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 10708 10906 10764 10908
rect 10788 10906 10844 10908
rect 10868 10906 10924 10908
rect 10948 10906 11004 10908
rect 10708 10854 10754 10906
rect 10754 10854 10764 10906
rect 10788 10854 10818 10906
rect 10818 10854 10830 10906
rect 10830 10854 10844 10906
rect 10868 10854 10882 10906
rect 10882 10854 10894 10906
rect 10894 10854 10924 10906
rect 10948 10854 10958 10906
rect 10958 10854 11004 10906
rect 10708 10852 10764 10854
rect 10788 10852 10844 10854
rect 10868 10852 10924 10854
rect 10948 10852 11004 10854
rect 9489 10362 9545 10364
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9489 10310 9535 10362
rect 9535 10310 9545 10362
rect 9569 10310 9599 10362
rect 9599 10310 9611 10362
rect 9611 10310 9625 10362
rect 9649 10310 9663 10362
rect 9663 10310 9675 10362
rect 9675 10310 9705 10362
rect 9729 10310 9739 10362
rect 9739 10310 9785 10362
rect 9489 10308 9545 10310
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
<< metal3 >>
rect 2165 15808 2481 15809
rect 2165 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2481 15808
rect 2165 15743 2481 15744
rect 4603 15808 4919 15809
rect 4603 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4919 15808
rect 4603 15743 4919 15744
rect 7041 15808 7357 15809
rect 7041 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7357 15808
rect 7041 15743 7357 15744
rect 9479 15808 9795 15809
rect 9479 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9795 15808
rect 9479 15743 9795 15744
rect 3384 15264 3700 15265
rect 3384 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3700 15264
rect 3384 15199 3700 15200
rect 5822 15264 6138 15265
rect 5822 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6138 15264
rect 5822 15199 6138 15200
rect 8260 15264 8576 15265
rect 8260 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8576 15264
rect 8260 15199 8576 15200
rect 10698 15264 11014 15265
rect 10698 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11014 15264
rect 10698 15199 11014 15200
rect 2165 14720 2481 14721
rect 2165 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2481 14720
rect 2165 14655 2481 14656
rect 4603 14720 4919 14721
rect 4603 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4919 14720
rect 4603 14655 4919 14656
rect 7041 14720 7357 14721
rect 7041 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7357 14720
rect 7041 14655 7357 14656
rect 9479 14720 9795 14721
rect 9479 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9795 14720
rect 9479 14655 9795 14656
rect 5717 14378 5783 14381
rect 7097 14378 7163 14381
rect 5717 14376 7163 14378
rect 5717 14320 5722 14376
rect 5778 14320 7102 14376
rect 7158 14320 7163 14376
rect 5717 14318 7163 14320
rect 5717 14315 5783 14318
rect 7097 14315 7163 14318
rect 3384 14176 3700 14177
rect 3384 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3700 14176
rect 3384 14111 3700 14112
rect 5822 14176 6138 14177
rect 5822 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6138 14176
rect 5822 14111 6138 14112
rect 8260 14176 8576 14177
rect 8260 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8576 14176
rect 8260 14111 8576 14112
rect 10698 14176 11014 14177
rect 10698 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11014 14176
rect 10698 14111 11014 14112
rect 2165 13632 2481 13633
rect 2165 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2481 13632
rect 2165 13567 2481 13568
rect 4603 13632 4919 13633
rect 4603 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4919 13632
rect 4603 13567 4919 13568
rect 7041 13632 7357 13633
rect 7041 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7357 13632
rect 7041 13567 7357 13568
rect 9479 13632 9795 13633
rect 9479 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9795 13632
rect 9479 13567 9795 13568
rect 3384 13088 3700 13089
rect 3384 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3700 13088
rect 3384 13023 3700 13024
rect 5822 13088 6138 13089
rect 5822 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6138 13088
rect 5822 13023 6138 13024
rect 8260 13088 8576 13089
rect 8260 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8576 13088
rect 8260 13023 8576 13024
rect 10698 13088 11014 13089
rect 10698 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11014 13088
rect 10698 13023 11014 13024
rect 2165 12544 2481 12545
rect 2165 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2481 12544
rect 2165 12479 2481 12480
rect 4603 12544 4919 12545
rect 4603 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4919 12544
rect 4603 12479 4919 12480
rect 7041 12544 7357 12545
rect 7041 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7357 12544
rect 7041 12479 7357 12480
rect 9479 12544 9795 12545
rect 9479 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9795 12544
rect 9479 12479 9795 12480
rect 3384 12000 3700 12001
rect 3384 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3700 12000
rect 3384 11935 3700 11936
rect 5822 12000 6138 12001
rect 5822 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6138 12000
rect 5822 11935 6138 11936
rect 8260 12000 8576 12001
rect 8260 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8576 12000
rect 8260 11935 8576 11936
rect 10698 12000 11014 12001
rect 10698 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11014 12000
rect 10698 11935 11014 11936
rect 2165 11456 2481 11457
rect 2165 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2481 11456
rect 2165 11391 2481 11392
rect 4603 11456 4919 11457
rect 4603 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4919 11456
rect 4603 11391 4919 11392
rect 7041 11456 7357 11457
rect 7041 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7357 11456
rect 7041 11391 7357 11392
rect 9479 11456 9795 11457
rect 9479 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9795 11456
rect 9479 11391 9795 11392
rect 3384 10912 3700 10913
rect 3384 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3700 10912
rect 3384 10847 3700 10848
rect 5822 10912 6138 10913
rect 5822 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6138 10912
rect 5822 10847 6138 10848
rect 8260 10912 8576 10913
rect 8260 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8576 10912
rect 8260 10847 8576 10848
rect 10698 10912 11014 10913
rect 10698 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11014 10912
rect 10698 10847 11014 10848
rect 2165 10368 2481 10369
rect 2165 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2481 10368
rect 2165 10303 2481 10304
rect 4603 10368 4919 10369
rect 4603 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4919 10368
rect 4603 10303 4919 10304
rect 7041 10368 7357 10369
rect 7041 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7357 10368
rect 7041 10303 7357 10304
rect 9479 10368 9795 10369
rect 9479 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9795 10368
rect 9479 10303 9795 10304
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
<< via3 >>
rect 2171 15804 2235 15808
rect 2171 15748 2175 15804
rect 2175 15748 2231 15804
rect 2231 15748 2235 15804
rect 2171 15744 2235 15748
rect 2251 15804 2315 15808
rect 2251 15748 2255 15804
rect 2255 15748 2311 15804
rect 2311 15748 2315 15804
rect 2251 15744 2315 15748
rect 2331 15804 2395 15808
rect 2331 15748 2335 15804
rect 2335 15748 2391 15804
rect 2391 15748 2395 15804
rect 2331 15744 2395 15748
rect 2411 15804 2475 15808
rect 2411 15748 2415 15804
rect 2415 15748 2471 15804
rect 2471 15748 2475 15804
rect 2411 15744 2475 15748
rect 4609 15804 4673 15808
rect 4609 15748 4613 15804
rect 4613 15748 4669 15804
rect 4669 15748 4673 15804
rect 4609 15744 4673 15748
rect 4689 15804 4753 15808
rect 4689 15748 4693 15804
rect 4693 15748 4749 15804
rect 4749 15748 4753 15804
rect 4689 15744 4753 15748
rect 4769 15804 4833 15808
rect 4769 15748 4773 15804
rect 4773 15748 4829 15804
rect 4829 15748 4833 15804
rect 4769 15744 4833 15748
rect 4849 15804 4913 15808
rect 4849 15748 4853 15804
rect 4853 15748 4909 15804
rect 4909 15748 4913 15804
rect 4849 15744 4913 15748
rect 7047 15804 7111 15808
rect 7047 15748 7051 15804
rect 7051 15748 7107 15804
rect 7107 15748 7111 15804
rect 7047 15744 7111 15748
rect 7127 15804 7191 15808
rect 7127 15748 7131 15804
rect 7131 15748 7187 15804
rect 7187 15748 7191 15804
rect 7127 15744 7191 15748
rect 7207 15804 7271 15808
rect 7207 15748 7211 15804
rect 7211 15748 7267 15804
rect 7267 15748 7271 15804
rect 7207 15744 7271 15748
rect 7287 15804 7351 15808
rect 7287 15748 7291 15804
rect 7291 15748 7347 15804
rect 7347 15748 7351 15804
rect 7287 15744 7351 15748
rect 9485 15804 9549 15808
rect 9485 15748 9489 15804
rect 9489 15748 9545 15804
rect 9545 15748 9549 15804
rect 9485 15744 9549 15748
rect 9565 15804 9629 15808
rect 9565 15748 9569 15804
rect 9569 15748 9625 15804
rect 9625 15748 9629 15804
rect 9565 15744 9629 15748
rect 9645 15804 9709 15808
rect 9645 15748 9649 15804
rect 9649 15748 9705 15804
rect 9705 15748 9709 15804
rect 9645 15744 9709 15748
rect 9725 15804 9789 15808
rect 9725 15748 9729 15804
rect 9729 15748 9785 15804
rect 9785 15748 9789 15804
rect 9725 15744 9789 15748
rect 3390 15260 3454 15264
rect 3390 15204 3394 15260
rect 3394 15204 3450 15260
rect 3450 15204 3454 15260
rect 3390 15200 3454 15204
rect 3470 15260 3534 15264
rect 3470 15204 3474 15260
rect 3474 15204 3530 15260
rect 3530 15204 3534 15260
rect 3470 15200 3534 15204
rect 3550 15260 3614 15264
rect 3550 15204 3554 15260
rect 3554 15204 3610 15260
rect 3610 15204 3614 15260
rect 3550 15200 3614 15204
rect 3630 15260 3694 15264
rect 3630 15204 3634 15260
rect 3634 15204 3690 15260
rect 3690 15204 3694 15260
rect 3630 15200 3694 15204
rect 5828 15260 5892 15264
rect 5828 15204 5832 15260
rect 5832 15204 5888 15260
rect 5888 15204 5892 15260
rect 5828 15200 5892 15204
rect 5908 15260 5972 15264
rect 5908 15204 5912 15260
rect 5912 15204 5968 15260
rect 5968 15204 5972 15260
rect 5908 15200 5972 15204
rect 5988 15260 6052 15264
rect 5988 15204 5992 15260
rect 5992 15204 6048 15260
rect 6048 15204 6052 15260
rect 5988 15200 6052 15204
rect 6068 15260 6132 15264
rect 6068 15204 6072 15260
rect 6072 15204 6128 15260
rect 6128 15204 6132 15260
rect 6068 15200 6132 15204
rect 8266 15260 8330 15264
rect 8266 15204 8270 15260
rect 8270 15204 8326 15260
rect 8326 15204 8330 15260
rect 8266 15200 8330 15204
rect 8346 15260 8410 15264
rect 8346 15204 8350 15260
rect 8350 15204 8406 15260
rect 8406 15204 8410 15260
rect 8346 15200 8410 15204
rect 8426 15260 8490 15264
rect 8426 15204 8430 15260
rect 8430 15204 8486 15260
rect 8486 15204 8490 15260
rect 8426 15200 8490 15204
rect 8506 15260 8570 15264
rect 8506 15204 8510 15260
rect 8510 15204 8566 15260
rect 8566 15204 8570 15260
rect 8506 15200 8570 15204
rect 10704 15260 10768 15264
rect 10704 15204 10708 15260
rect 10708 15204 10764 15260
rect 10764 15204 10768 15260
rect 10704 15200 10768 15204
rect 10784 15260 10848 15264
rect 10784 15204 10788 15260
rect 10788 15204 10844 15260
rect 10844 15204 10848 15260
rect 10784 15200 10848 15204
rect 10864 15260 10928 15264
rect 10864 15204 10868 15260
rect 10868 15204 10924 15260
rect 10924 15204 10928 15260
rect 10864 15200 10928 15204
rect 10944 15260 11008 15264
rect 10944 15204 10948 15260
rect 10948 15204 11004 15260
rect 11004 15204 11008 15260
rect 10944 15200 11008 15204
rect 2171 14716 2235 14720
rect 2171 14660 2175 14716
rect 2175 14660 2231 14716
rect 2231 14660 2235 14716
rect 2171 14656 2235 14660
rect 2251 14716 2315 14720
rect 2251 14660 2255 14716
rect 2255 14660 2311 14716
rect 2311 14660 2315 14716
rect 2251 14656 2315 14660
rect 2331 14716 2395 14720
rect 2331 14660 2335 14716
rect 2335 14660 2391 14716
rect 2391 14660 2395 14716
rect 2331 14656 2395 14660
rect 2411 14716 2475 14720
rect 2411 14660 2415 14716
rect 2415 14660 2471 14716
rect 2471 14660 2475 14716
rect 2411 14656 2475 14660
rect 4609 14716 4673 14720
rect 4609 14660 4613 14716
rect 4613 14660 4669 14716
rect 4669 14660 4673 14716
rect 4609 14656 4673 14660
rect 4689 14716 4753 14720
rect 4689 14660 4693 14716
rect 4693 14660 4749 14716
rect 4749 14660 4753 14716
rect 4689 14656 4753 14660
rect 4769 14716 4833 14720
rect 4769 14660 4773 14716
rect 4773 14660 4829 14716
rect 4829 14660 4833 14716
rect 4769 14656 4833 14660
rect 4849 14716 4913 14720
rect 4849 14660 4853 14716
rect 4853 14660 4909 14716
rect 4909 14660 4913 14716
rect 4849 14656 4913 14660
rect 7047 14716 7111 14720
rect 7047 14660 7051 14716
rect 7051 14660 7107 14716
rect 7107 14660 7111 14716
rect 7047 14656 7111 14660
rect 7127 14716 7191 14720
rect 7127 14660 7131 14716
rect 7131 14660 7187 14716
rect 7187 14660 7191 14716
rect 7127 14656 7191 14660
rect 7207 14716 7271 14720
rect 7207 14660 7211 14716
rect 7211 14660 7267 14716
rect 7267 14660 7271 14716
rect 7207 14656 7271 14660
rect 7287 14716 7351 14720
rect 7287 14660 7291 14716
rect 7291 14660 7347 14716
rect 7347 14660 7351 14716
rect 7287 14656 7351 14660
rect 9485 14716 9549 14720
rect 9485 14660 9489 14716
rect 9489 14660 9545 14716
rect 9545 14660 9549 14716
rect 9485 14656 9549 14660
rect 9565 14716 9629 14720
rect 9565 14660 9569 14716
rect 9569 14660 9625 14716
rect 9625 14660 9629 14716
rect 9565 14656 9629 14660
rect 9645 14716 9709 14720
rect 9645 14660 9649 14716
rect 9649 14660 9705 14716
rect 9705 14660 9709 14716
rect 9645 14656 9709 14660
rect 9725 14716 9789 14720
rect 9725 14660 9729 14716
rect 9729 14660 9785 14716
rect 9785 14660 9789 14716
rect 9725 14656 9789 14660
rect 3390 14172 3454 14176
rect 3390 14116 3394 14172
rect 3394 14116 3450 14172
rect 3450 14116 3454 14172
rect 3390 14112 3454 14116
rect 3470 14172 3534 14176
rect 3470 14116 3474 14172
rect 3474 14116 3530 14172
rect 3530 14116 3534 14172
rect 3470 14112 3534 14116
rect 3550 14172 3614 14176
rect 3550 14116 3554 14172
rect 3554 14116 3610 14172
rect 3610 14116 3614 14172
rect 3550 14112 3614 14116
rect 3630 14172 3694 14176
rect 3630 14116 3634 14172
rect 3634 14116 3690 14172
rect 3690 14116 3694 14172
rect 3630 14112 3694 14116
rect 5828 14172 5892 14176
rect 5828 14116 5832 14172
rect 5832 14116 5888 14172
rect 5888 14116 5892 14172
rect 5828 14112 5892 14116
rect 5908 14172 5972 14176
rect 5908 14116 5912 14172
rect 5912 14116 5968 14172
rect 5968 14116 5972 14172
rect 5908 14112 5972 14116
rect 5988 14172 6052 14176
rect 5988 14116 5992 14172
rect 5992 14116 6048 14172
rect 6048 14116 6052 14172
rect 5988 14112 6052 14116
rect 6068 14172 6132 14176
rect 6068 14116 6072 14172
rect 6072 14116 6128 14172
rect 6128 14116 6132 14172
rect 6068 14112 6132 14116
rect 8266 14172 8330 14176
rect 8266 14116 8270 14172
rect 8270 14116 8326 14172
rect 8326 14116 8330 14172
rect 8266 14112 8330 14116
rect 8346 14172 8410 14176
rect 8346 14116 8350 14172
rect 8350 14116 8406 14172
rect 8406 14116 8410 14172
rect 8346 14112 8410 14116
rect 8426 14172 8490 14176
rect 8426 14116 8430 14172
rect 8430 14116 8486 14172
rect 8486 14116 8490 14172
rect 8426 14112 8490 14116
rect 8506 14172 8570 14176
rect 8506 14116 8510 14172
rect 8510 14116 8566 14172
rect 8566 14116 8570 14172
rect 8506 14112 8570 14116
rect 10704 14172 10768 14176
rect 10704 14116 10708 14172
rect 10708 14116 10764 14172
rect 10764 14116 10768 14172
rect 10704 14112 10768 14116
rect 10784 14172 10848 14176
rect 10784 14116 10788 14172
rect 10788 14116 10844 14172
rect 10844 14116 10848 14172
rect 10784 14112 10848 14116
rect 10864 14172 10928 14176
rect 10864 14116 10868 14172
rect 10868 14116 10924 14172
rect 10924 14116 10928 14172
rect 10864 14112 10928 14116
rect 10944 14172 11008 14176
rect 10944 14116 10948 14172
rect 10948 14116 11004 14172
rect 11004 14116 11008 14172
rect 10944 14112 11008 14116
rect 2171 13628 2235 13632
rect 2171 13572 2175 13628
rect 2175 13572 2231 13628
rect 2231 13572 2235 13628
rect 2171 13568 2235 13572
rect 2251 13628 2315 13632
rect 2251 13572 2255 13628
rect 2255 13572 2311 13628
rect 2311 13572 2315 13628
rect 2251 13568 2315 13572
rect 2331 13628 2395 13632
rect 2331 13572 2335 13628
rect 2335 13572 2391 13628
rect 2391 13572 2395 13628
rect 2331 13568 2395 13572
rect 2411 13628 2475 13632
rect 2411 13572 2415 13628
rect 2415 13572 2471 13628
rect 2471 13572 2475 13628
rect 2411 13568 2475 13572
rect 4609 13628 4673 13632
rect 4609 13572 4613 13628
rect 4613 13572 4669 13628
rect 4669 13572 4673 13628
rect 4609 13568 4673 13572
rect 4689 13628 4753 13632
rect 4689 13572 4693 13628
rect 4693 13572 4749 13628
rect 4749 13572 4753 13628
rect 4689 13568 4753 13572
rect 4769 13628 4833 13632
rect 4769 13572 4773 13628
rect 4773 13572 4829 13628
rect 4829 13572 4833 13628
rect 4769 13568 4833 13572
rect 4849 13628 4913 13632
rect 4849 13572 4853 13628
rect 4853 13572 4909 13628
rect 4909 13572 4913 13628
rect 4849 13568 4913 13572
rect 7047 13628 7111 13632
rect 7047 13572 7051 13628
rect 7051 13572 7107 13628
rect 7107 13572 7111 13628
rect 7047 13568 7111 13572
rect 7127 13628 7191 13632
rect 7127 13572 7131 13628
rect 7131 13572 7187 13628
rect 7187 13572 7191 13628
rect 7127 13568 7191 13572
rect 7207 13628 7271 13632
rect 7207 13572 7211 13628
rect 7211 13572 7267 13628
rect 7267 13572 7271 13628
rect 7207 13568 7271 13572
rect 7287 13628 7351 13632
rect 7287 13572 7291 13628
rect 7291 13572 7347 13628
rect 7347 13572 7351 13628
rect 7287 13568 7351 13572
rect 9485 13628 9549 13632
rect 9485 13572 9489 13628
rect 9489 13572 9545 13628
rect 9545 13572 9549 13628
rect 9485 13568 9549 13572
rect 9565 13628 9629 13632
rect 9565 13572 9569 13628
rect 9569 13572 9625 13628
rect 9625 13572 9629 13628
rect 9565 13568 9629 13572
rect 9645 13628 9709 13632
rect 9645 13572 9649 13628
rect 9649 13572 9705 13628
rect 9705 13572 9709 13628
rect 9645 13568 9709 13572
rect 9725 13628 9789 13632
rect 9725 13572 9729 13628
rect 9729 13572 9785 13628
rect 9785 13572 9789 13628
rect 9725 13568 9789 13572
rect 3390 13084 3454 13088
rect 3390 13028 3394 13084
rect 3394 13028 3450 13084
rect 3450 13028 3454 13084
rect 3390 13024 3454 13028
rect 3470 13084 3534 13088
rect 3470 13028 3474 13084
rect 3474 13028 3530 13084
rect 3530 13028 3534 13084
rect 3470 13024 3534 13028
rect 3550 13084 3614 13088
rect 3550 13028 3554 13084
rect 3554 13028 3610 13084
rect 3610 13028 3614 13084
rect 3550 13024 3614 13028
rect 3630 13084 3694 13088
rect 3630 13028 3634 13084
rect 3634 13028 3690 13084
rect 3690 13028 3694 13084
rect 3630 13024 3694 13028
rect 5828 13084 5892 13088
rect 5828 13028 5832 13084
rect 5832 13028 5888 13084
rect 5888 13028 5892 13084
rect 5828 13024 5892 13028
rect 5908 13084 5972 13088
rect 5908 13028 5912 13084
rect 5912 13028 5968 13084
rect 5968 13028 5972 13084
rect 5908 13024 5972 13028
rect 5988 13084 6052 13088
rect 5988 13028 5992 13084
rect 5992 13028 6048 13084
rect 6048 13028 6052 13084
rect 5988 13024 6052 13028
rect 6068 13084 6132 13088
rect 6068 13028 6072 13084
rect 6072 13028 6128 13084
rect 6128 13028 6132 13084
rect 6068 13024 6132 13028
rect 8266 13084 8330 13088
rect 8266 13028 8270 13084
rect 8270 13028 8326 13084
rect 8326 13028 8330 13084
rect 8266 13024 8330 13028
rect 8346 13084 8410 13088
rect 8346 13028 8350 13084
rect 8350 13028 8406 13084
rect 8406 13028 8410 13084
rect 8346 13024 8410 13028
rect 8426 13084 8490 13088
rect 8426 13028 8430 13084
rect 8430 13028 8486 13084
rect 8486 13028 8490 13084
rect 8426 13024 8490 13028
rect 8506 13084 8570 13088
rect 8506 13028 8510 13084
rect 8510 13028 8566 13084
rect 8566 13028 8570 13084
rect 8506 13024 8570 13028
rect 10704 13084 10768 13088
rect 10704 13028 10708 13084
rect 10708 13028 10764 13084
rect 10764 13028 10768 13084
rect 10704 13024 10768 13028
rect 10784 13084 10848 13088
rect 10784 13028 10788 13084
rect 10788 13028 10844 13084
rect 10844 13028 10848 13084
rect 10784 13024 10848 13028
rect 10864 13084 10928 13088
rect 10864 13028 10868 13084
rect 10868 13028 10924 13084
rect 10924 13028 10928 13084
rect 10864 13024 10928 13028
rect 10944 13084 11008 13088
rect 10944 13028 10948 13084
rect 10948 13028 11004 13084
rect 11004 13028 11008 13084
rect 10944 13024 11008 13028
rect 2171 12540 2235 12544
rect 2171 12484 2175 12540
rect 2175 12484 2231 12540
rect 2231 12484 2235 12540
rect 2171 12480 2235 12484
rect 2251 12540 2315 12544
rect 2251 12484 2255 12540
rect 2255 12484 2311 12540
rect 2311 12484 2315 12540
rect 2251 12480 2315 12484
rect 2331 12540 2395 12544
rect 2331 12484 2335 12540
rect 2335 12484 2391 12540
rect 2391 12484 2395 12540
rect 2331 12480 2395 12484
rect 2411 12540 2475 12544
rect 2411 12484 2415 12540
rect 2415 12484 2471 12540
rect 2471 12484 2475 12540
rect 2411 12480 2475 12484
rect 4609 12540 4673 12544
rect 4609 12484 4613 12540
rect 4613 12484 4669 12540
rect 4669 12484 4673 12540
rect 4609 12480 4673 12484
rect 4689 12540 4753 12544
rect 4689 12484 4693 12540
rect 4693 12484 4749 12540
rect 4749 12484 4753 12540
rect 4689 12480 4753 12484
rect 4769 12540 4833 12544
rect 4769 12484 4773 12540
rect 4773 12484 4829 12540
rect 4829 12484 4833 12540
rect 4769 12480 4833 12484
rect 4849 12540 4913 12544
rect 4849 12484 4853 12540
rect 4853 12484 4909 12540
rect 4909 12484 4913 12540
rect 4849 12480 4913 12484
rect 7047 12540 7111 12544
rect 7047 12484 7051 12540
rect 7051 12484 7107 12540
rect 7107 12484 7111 12540
rect 7047 12480 7111 12484
rect 7127 12540 7191 12544
rect 7127 12484 7131 12540
rect 7131 12484 7187 12540
rect 7187 12484 7191 12540
rect 7127 12480 7191 12484
rect 7207 12540 7271 12544
rect 7207 12484 7211 12540
rect 7211 12484 7267 12540
rect 7267 12484 7271 12540
rect 7207 12480 7271 12484
rect 7287 12540 7351 12544
rect 7287 12484 7291 12540
rect 7291 12484 7347 12540
rect 7347 12484 7351 12540
rect 7287 12480 7351 12484
rect 9485 12540 9549 12544
rect 9485 12484 9489 12540
rect 9489 12484 9545 12540
rect 9545 12484 9549 12540
rect 9485 12480 9549 12484
rect 9565 12540 9629 12544
rect 9565 12484 9569 12540
rect 9569 12484 9625 12540
rect 9625 12484 9629 12540
rect 9565 12480 9629 12484
rect 9645 12540 9709 12544
rect 9645 12484 9649 12540
rect 9649 12484 9705 12540
rect 9705 12484 9709 12540
rect 9645 12480 9709 12484
rect 9725 12540 9789 12544
rect 9725 12484 9729 12540
rect 9729 12484 9785 12540
rect 9785 12484 9789 12540
rect 9725 12480 9789 12484
rect 3390 11996 3454 12000
rect 3390 11940 3394 11996
rect 3394 11940 3450 11996
rect 3450 11940 3454 11996
rect 3390 11936 3454 11940
rect 3470 11996 3534 12000
rect 3470 11940 3474 11996
rect 3474 11940 3530 11996
rect 3530 11940 3534 11996
rect 3470 11936 3534 11940
rect 3550 11996 3614 12000
rect 3550 11940 3554 11996
rect 3554 11940 3610 11996
rect 3610 11940 3614 11996
rect 3550 11936 3614 11940
rect 3630 11996 3694 12000
rect 3630 11940 3634 11996
rect 3634 11940 3690 11996
rect 3690 11940 3694 11996
rect 3630 11936 3694 11940
rect 5828 11996 5892 12000
rect 5828 11940 5832 11996
rect 5832 11940 5888 11996
rect 5888 11940 5892 11996
rect 5828 11936 5892 11940
rect 5908 11996 5972 12000
rect 5908 11940 5912 11996
rect 5912 11940 5968 11996
rect 5968 11940 5972 11996
rect 5908 11936 5972 11940
rect 5988 11996 6052 12000
rect 5988 11940 5992 11996
rect 5992 11940 6048 11996
rect 6048 11940 6052 11996
rect 5988 11936 6052 11940
rect 6068 11996 6132 12000
rect 6068 11940 6072 11996
rect 6072 11940 6128 11996
rect 6128 11940 6132 11996
rect 6068 11936 6132 11940
rect 8266 11996 8330 12000
rect 8266 11940 8270 11996
rect 8270 11940 8326 11996
rect 8326 11940 8330 11996
rect 8266 11936 8330 11940
rect 8346 11996 8410 12000
rect 8346 11940 8350 11996
rect 8350 11940 8406 11996
rect 8406 11940 8410 11996
rect 8346 11936 8410 11940
rect 8426 11996 8490 12000
rect 8426 11940 8430 11996
rect 8430 11940 8486 11996
rect 8486 11940 8490 11996
rect 8426 11936 8490 11940
rect 8506 11996 8570 12000
rect 8506 11940 8510 11996
rect 8510 11940 8566 11996
rect 8566 11940 8570 11996
rect 8506 11936 8570 11940
rect 10704 11996 10768 12000
rect 10704 11940 10708 11996
rect 10708 11940 10764 11996
rect 10764 11940 10768 11996
rect 10704 11936 10768 11940
rect 10784 11996 10848 12000
rect 10784 11940 10788 11996
rect 10788 11940 10844 11996
rect 10844 11940 10848 11996
rect 10784 11936 10848 11940
rect 10864 11996 10928 12000
rect 10864 11940 10868 11996
rect 10868 11940 10924 11996
rect 10924 11940 10928 11996
rect 10864 11936 10928 11940
rect 10944 11996 11008 12000
rect 10944 11940 10948 11996
rect 10948 11940 11004 11996
rect 11004 11940 11008 11996
rect 10944 11936 11008 11940
rect 2171 11452 2235 11456
rect 2171 11396 2175 11452
rect 2175 11396 2231 11452
rect 2231 11396 2235 11452
rect 2171 11392 2235 11396
rect 2251 11452 2315 11456
rect 2251 11396 2255 11452
rect 2255 11396 2311 11452
rect 2311 11396 2315 11452
rect 2251 11392 2315 11396
rect 2331 11452 2395 11456
rect 2331 11396 2335 11452
rect 2335 11396 2391 11452
rect 2391 11396 2395 11452
rect 2331 11392 2395 11396
rect 2411 11452 2475 11456
rect 2411 11396 2415 11452
rect 2415 11396 2471 11452
rect 2471 11396 2475 11452
rect 2411 11392 2475 11396
rect 4609 11452 4673 11456
rect 4609 11396 4613 11452
rect 4613 11396 4669 11452
rect 4669 11396 4673 11452
rect 4609 11392 4673 11396
rect 4689 11452 4753 11456
rect 4689 11396 4693 11452
rect 4693 11396 4749 11452
rect 4749 11396 4753 11452
rect 4689 11392 4753 11396
rect 4769 11452 4833 11456
rect 4769 11396 4773 11452
rect 4773 11396 4829 11452
rect 4829 11396 4833 11452
rect 4769 11392 4833 11396
rect 4849 11452 4913 11456
rect 4849 11396 4853 11452
rect 4853 11396 4909 11452
rect 4909 11396 4913 11452
rect 4849 11392 4913 11396
rect 7047 11452 7111 11456
rect 7047 11396 7051 11452
rect 7051 11396 7107 11452
rect 7107 11396 7111 11452
rect 7047 11392 7111 11396
rect 7127 11452 7191 11456
rect 7127 11396 7131 11452
rect 7131 11396 7187 11452
rect 7187 11396 7191 11452
rect 7127 11392 7191 11396
rect 7207 11452 7271 11456
rect 7207 11396 7211 11452
rect 7211 11396 7267 11452
rect 7267 11396 7271 11452
rect 7207 11392 7271 11396
rect 7287 11452 7351 11456
rect 7287 11396 7291 11452
rect 7291 11396 7347 11452
rect 7347 11396 7351 11452
rect 7287 11392 7351 11396
rect 9485 11452 9549 11456
rect 9485 11396 9489 11452
rect 9489 11396 9545 11452
rect 9545 11396 9549 11452
rect 9485 11392 9549 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 3390 10908 3454 10912
rect 3390 10852 3394 10908
rect 3394 10852 3450 10908
rect 3450 10852 3454 10908
rect 3390 10848 3454 10852
rect 3470 10908 3534 10912
rect 3470 10852 3474 10908
rect 3474 10852 3530 10908
rect 3530 10852 3534 10908
rect 3470 10848 3534 10852
rect 3550 10908 3614 10912
rect 3550 10852 3554 10908
rect 3554 10852 3610 10908
rect 3610 10852 3614 10908
rect 3550 10848 3614 10852
rect 3630 10908 3694 10912
rect 3630 10852 3634 10908
rect 3634 10852 3690 10908
rect 3690 10852 3694 10908
rect 3630 10848 3694 10852
rect 5828 10908 5892 10912
rect 5828 10852 5832 10908
rect 5832 10852 5888 10908
rect 5888 10852 5892 10908
rect 5828 10848 5892 10852
rect 5908 10908 5972 10912
rect 5908 10852 5912 10908
rect 5912 10852 5968 10908
rect 5968 10852 5972 10908
rect 5908 10848 5972 10852
rect 5988 10908 6052 10912
rect 5988 10852 5992 10908
rect 5992 10852 6048 10908
rect 6048 10852 6052 10908
rect 5988 10848 6052 10852
rect 6068 10908 6132 10912
rect 6068 10852 6072 10908
rect 6072 10852 6128 10908
rect 6128 10852 6132 10908
rect 6068 10848 6132 10852
rect 8266 10908 8330 10912
rect 8266 10852 8270 10908
rect 8270 10852 8326 10908
rect 8326 10852 8330 10908
rect 8266 10848 8330 10852
rect 8346 10908 8410 10912
rect 8346 10852 8350 10908
rect 8350 10852 8406 10908
rect 8406 10852 8410 10908
rect 8346 10848 8410 10852
rect 8426 10908 8490 10912
rect 8426 10852 8430 10908
rect 8430 10852 8486 10908
rect 8486 10852 8490 10908
rect 8426 10848 8490 10852
rect 8506 10908 8570 10912
rect 8506 10852 8510 10908
rect 8510 10852 8566 10908
rect 8566 10852 8570 10908
rect 8506 10848 8570 10852
rect 10704 10908 10768 10912
rect 10704 10852 10708 10908
rect 10708 10852 10764 10908
rect 10764 10852 10768 10908
rect 10704 10848 10768 10852
rect 10784 10908 10848 10912
rect 10784 10852 10788 10908
rect 10788 10852 10844 10908
rect 10844 10852 10848 10908
rect 10784 10848 10848 10852
rect 10864 10908 10928 10912
rect 10864 10852 10868 10908
rect 10868 10852 10924 10908
rect 10924 10852 10928 10908
rect 10864 10848 10928 10852
rect 10944 10908 11008 10912
rect 10944 10852 10948 10908
rect 10948 10852 11004 10908
rect 11004 10852 11008 10908
rect 10944 10848 11008 10852
rect 2171 10364 2235 10368
rect 2171 10308 2175 10364
rect 2175 10308 2231 10364
rect 2231 10308 2235 10364
rect 2171 10304 2235 10308
rect 2251 10364 2315 10368
rect 2251 10308 2255 10364
rect 2255 10308 2311 10364
rect 2311 10308 2315 10364
rect 2251 10304 2315 10308
rect 2331 10364 2395 10368
rect 2331 10308 2335 10364
rect 2335 10308 2391 10364
rect 2391 10308 2395 10364
rect 2331 10304 2395 10308
rect 2411 10364 2475 10368
rect 2411 10308 2415 10364
rect 2415 10308 2471 10364
rect 2471 10308 2475 10364
rect 2411 10304 2475 10308
rect 4609 10364 4673 10368
rect 4609 10308 4613 10364
rect 4613 10308 4669 10364
rect 4669 10308 4673 10364
rect 4609 10304 4673 10308
rect 4689 10364 4753 10368
rect 4689 10308 4693 10364
rect 4693 10308 4749 10364
rect 4749 10308 4753 10364
rect 4689 10304 4753 10308
rect 4769 10364 4833 10368
rect 4769 10308 4773 10364
rect 4773 10308 4829 10364
rect 4829 10308 4833 10364
rect 4769 10304 4833 10308
rect 4849 10364 4913 10368
rect 4849 10308 4853 10364
rect 4853 10308 4909 10364
rect 4909 10308 4913 10364
rect 4849 10304 4913 10308
rect 7047 10364 7111 10368
rect 7047 10308 7051 10364
rect 7051 10308 7107 10364
rect 7107 10308 7111 10364
rect 7047 10304 7111 10308
rect 7127 10364 7191 10368
rect 7127 10308 7131 10364
rect 7131 10308 7187 10364
rect 7187 10308 7191 10364
rect 7127 10304 7191 10308
rect 7207 10364 7271 10368
rect 7207 10308 7211 10364
rect 7211 10308 7267 10364
rect 7267 10308 7271 10364
rect 7207 10304 7271 10308
rect 7287 10364 7351 10368
rect 7287 10308 7291 10364
rect 7291 10308 7347 10364
rect 7347 10308 7351 10364
rect 7287 10304 7351 10308
rect 9485 10364 9549 10368
rect 9485 10308 9489 10364
rect 9489 10308 9545 10364
rect 9545 10308 9549 10364
rect 9485 10304 9549 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 15808 2483 15824
rect 2163 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2483 15808
rect 2163 14720 2483 15744
rect 2163 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2483 14720
rect 2163 13632 2483 14656
rect 2163 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2483 13632
rect 2163 12544 2483 13568
rect 2163 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2483 12544
rect 2163 11456 2483 12480
rect 2163 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2483 11456
rect 2163 10368 2483 11392
rect 2163 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2483 10368
rect 2163 9280 2483 10304
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 15264 3702 15824
rect 3382 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3702 15264
rect 3382 14176 3702 15200
rect 3382 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3702 14176
rect 3382 13088 3702 14112
rect 3382 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3702 13088
rect 3382 12000 3702 13024
rect 3382 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3702 12000
rect 3382 10912 3702 11936
rect 3382 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3702 10912
rect 3382 9824 3702 10848
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 15808 4921 15824
rect 4601 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4921 15808
rect 4601 14720 4921 15744
rect 4601 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4921 14720
rect 4601 13632 4921 14656
rect 4601 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4921 13632
rect 4601 12544 4921 13568
rect 4601 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4921 12544
rect 4601 11456 4921 12480
rect 4601 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4921 11456
rect 4601 10368 4921 11392
rect 4601 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4921 10368
rect 4601 9280 4921 10304
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 15264 6140 15824
rect 5820 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6140 15264
rect 5820 14176 6140 15200
rect 5820 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6140 14176
rect 5820 13088 6140 14112
rect 5820 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6140 13088
rect 5820 12000 6140 13024
rect 5820 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6140 12000
rect 5820 10912 6140 11936
rect 5820 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6140 10912
rect 5820 9824 6140 10848
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 15808 7359 15824
rect 7039 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7359 15808
rect 7039 14720 7359 15744
rect 7039 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7359 14720
rect 7039 13632 7359 14656
rect 7039 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7359 13632
rect 7039 12544 7359 13568
rect 7039 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7359 12544
rect 7039 11456 7359 12480
rect 7039 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7359 11456
rect 7039 10368 7359 11392
rect 7039 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7359 10368
rect 7039 9280 7359 10304
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 15264 8578 15824
rect 8258 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8578 15264
rect 8258 14176 8578 15200
rect 8258 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8578 14176
rect 8258 13088 8578 14112
rect 8258 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8578 13088
rect 8258 12000 8578 13024
rect 8258 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8578 12000
rect 8258 10912 8578 11936
rect 8258 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8578 10912
rect 8258 9824 8578 10848
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 15808 9797 15824
rect 9477 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9797 15808
rect 9477 14720 9797 15744
rect 9477 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9797 14720
rect 9477 13632 9797 14656
rect 9477 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9797 13632
rect 9477 12544 9797 13568
rect 9477 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9797 12544
rect 9477 11456 9797 12480
rect 9477 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9797 11456
rect 9477 10368 9797 11392
rect 9477 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9797 10368
rect 9477 9280 9797 10304
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 15264 11016 15824
rect 10696 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11016 15264
rect 10696 14176 11016 15200
rect 10696 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11016 14176
rect 10696 13088 11016 14112
rect 10696 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11016 13088
rect 10696 12000 11016 13024
rect 10696 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11016 12000
rect 10696 10912 11016 11936
rect 10696 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11016 10912
rect 10696 9824 11016 10848
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 1932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 4784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 9844 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 10396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35
timestamp 1666464484
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1666464484
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1666464484
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1666464484
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1666464484
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1666464484
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_84
timestamp 1666464484
transform 1 0 8832 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_96
timestamp 1666464484
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_102
timestamp 1666464484
transform 1 0 10488 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1666464484
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_56
timestamp 1666464484
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1666464484
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1666464484
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_47
timestamp 1666464484
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_65
timestamp 1666464484
transform 1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1666464484
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1666464484
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1666464484
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 1666464484
transform 1 0 4416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1666464484
transform 1 0 4784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_56
timestamp 1666464484
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1666464484
transform 1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1666464484
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1666464484
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1666464484
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1666464484
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1666464484
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_84
timestamp 1666464484
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_96
timestamp 1666464484
transform 1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1666464484
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_38
timestamp 1666464484
transform 1 0 4600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1666464484
transform 1 0 5612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1666464484
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1666464484
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 1666464484
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1666464484
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_31
timestamp 1666464484
transform 1 0 3956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 1666464484
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1666464484
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1666464484
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_65
timestamp 1666464484
transform 1 0 7084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_77
timestamp 1666464484
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1666464484
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_19
timestamp 1666464484
transform 1 0 2852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1666464484
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 1666464484
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1666464484
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1666464484
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1666464484
transform 1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1666464484
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1666464484
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1666464484
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1666464484
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_63
timestamp 1666464484
transform 1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1666464484
transform 1 0 7544 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1666464484
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1666464484
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_44
timestamp 1666464484
transform 1 0 5152 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1666464484
transform 1 0 5888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1666464484
transform 1 0 6624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1666464484
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1666464484
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1666464484
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_22
timestamp 1666464484
transform 1 0 3128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1666464484
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1666464484
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1666464484
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_67
timestamp 1666464484
transform 1 0 7268 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_78
timestamp 1666464484
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_90
timestamp 1666464484
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1666464484
transform 1 0 10488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_7
timestamp 1666464484
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_19
timestamp 1666464484
transform 1 0 2852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_40
timestamp 1666464484
transform 1 0 4784 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_55
timestamp 1666464484
transform 1 0 6164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1666464484
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1666464484
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1666464484
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1666464484
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1666464484
transform 1 0 10396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1666464484
transform 1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_40
timestamp 1666464484
transform 1 0 4784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1666464484
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1666464484
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_61
timestamp 1666464484
transform 1 0 6716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_73
timestamp 1666464484
transform 1 0 7820 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_84
timestamp 1666464484
transform 1 0 8832 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1666464484
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1666464484
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1666464484
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1666464484
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_35
timestamp 1666464484
transform 1 0 4324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_49
timestamp 1666464484
transform 1 0 5612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_55
timestamp 1666464484
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_71
timestamp 1666464484
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1666464484
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1666464484
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _054_
timestamp 1666464484
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4140 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _058_
timestamp 1666464484
transform -1 0 3128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _060_
timestamp 1666464484
transform -1 0 3496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _063_
timestamp 1666464484
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _067_
timestamp 1666464484
transform -1 0 6164 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _068_
timestamp 1666464484
transform -1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _071_
timestamp 1666464484
transform -1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _072_
timestamp 1666464484
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7268 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _074_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _075_
timestamp 1666464484
transform -1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5888 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _077_
timestamp 1666464484
transform -1 0 5612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _078_
timestamp 1666464484
transform 1 0 4508 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _079_
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _080_
timestamp 1666464484
transform -1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _082_
timestamp 1666464484
transform 1 0 6624 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _083_
timestamp 1666464484
transform 1 0 5704 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6072 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5244 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _086_
timestamp 1666464484
transform -1 0 4600 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _087_
timestamp 1666464484
transform -1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _088_
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5612 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _090_
timestamp 1666464484
transform 1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _091_
timestamp 1666464484
transform -1 0 7084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6072 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7636 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _095_
timestamp 1666464484
transform -1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _096_
timestamp 1666464484
transform 1 0 6992 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _098_
timestamp 1666464484
transform -1 0 8004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 1666464484
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _101_
timestamp 1666464484
transform -1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _102_
timestamp 1666464484
transform 1 0 7360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _103_
timestamp 1666464484
transform 1 0 8004 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _104_
timestamp 1666464484
transform 1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _105_
timestamp 1666464484
transform -1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _106_
timestamp 1666464484
transform -1 0 8648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 1666464484
transform -1 0 8372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _108_
timestamp 1666464484
transform 1 0 8188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _109_
timestamp 1666464484
transform -1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 1666464484
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _111_
timestamp 1666464484
transform -1 0 9292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1666464484
transform 1 0 2300 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1666464484
transform -1 0 8648 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform 1 0 9476 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666464484
transform -1 0 10396 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1666464484
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
<< labels >>
flabel metal2 s 754 17200 810 18000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 2226 17200 2282 18000 0 FreeSans 224 90 0 0 io_in[1]
port 1 nsew signal input
flabel metal2 s 3698 17200 3754 18000 0 FreeSans 224 90 0 0 io_in[2]
port 2 nsew signal input
flabel metal2 s 5170 17200 5226 18000 0 FreeSans 224 90 0 0 io_in[3]
port 3 nsew signal input
flabel metal2 s 6642 17200 6698 18000 0 FreeSans 224 90 0 0 io_in[4]
port 4 nsew signal input
flabel metal2 s 8114 17200 8170 18000 0 FreeSans 224 90 0 0 io_in[5]
port 5 nsew signal input
flabel metal2 s 9586 17200 9642 18000 0 FreeSans 224 90 0 0 io_in[6]
port 6 nsew signal input
flabel metal2 s 11058 17200 11114 18000 0 FreeSans 224 90 0 0 io_in[7]
port 7 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 2163 2128 2483 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 4601 2128 4921 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7039 2128 7359 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 9477 2128 9797 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 3382 2128 3702 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 5980 15776 5980 15776 0 vccd1
rlabel via1 6060 15232 6060 15232 0 vssd1
rlabel metal1 3082 12206 3082 12206 0 _000_
rlabel metal1 2944 13226 2944 13226 0 _001_
rlabel metal1 2990 12818 2990 12818 0 _002_
rlabel metal2 3910 13804 3910 13804 0 _003_
rlabel metal1 3450 12614 3450 12614 0 _004_
rlabel metal2 4186 11152 4186 11152 0 _005_
rlabel metal2 2990 13770 2990 13770 0 _006_
rlabel metal1 4462 14314 4462 14314 0 _007_
rlabel metal1 4148 10778 4148 10778 0 _008_
rlabel metal1 4462 11730 4462 11730 0 _009_
rlabel metal1 4186 10064 4186 10064 0 _010_
rlabel metal2 4370 10234 4370 10234 0 _011_
rlabel metal2 5566 14144 5566 14144 0 _012_
rlabel metal1 6578 13872 6578 13872 0 _013_
rlabel metal2 6946 11322 6946 11322 0 _014_
rlabel metal2 6762 11118 6762 11118 0 _015_
rlabel metal1 7820 11118 7820 11118 0 _016_
rlabel metal1 6210 11186 6210 11186 0 _017_
rlabel metal1 6808 11322 6808 11322 0 _018_
rlabel metal2 6670 10200 6670 10200 0 _019_
rlabel metal1 6532 10234 6532 10234 0 _020_
rlabel metal2 5658 14348 5658 14348 0 _021_
rlabel metal1 4186 11254 4186 11254 0 _022_
rlabel metal1 5198 11186 5198 11186 0 _023_
rlabel via1 5198 11101 5198 11101 0 _024_
rlabel metal1 5796 11186 5796 11186 0 _025_
rlabel metal1 5842 10030 5842 10030 0 _026_
rlabel metal1 6854 9588 6854 9588 0 _027_
rlabel metal2 5750 9656 5750 9656 0 _028_
rlabel metal2 5842 9146 5842 9146 0 _029_
rlabel metal2 4370 11033 4370 11033 0 _030_
rlabel metal1 5060 10234 5060 10234 0 _031_
rlabel via1 5114 9962 5114 9962 0 _032_
rlabel metal1 5244 8942 5244 8942 0 _033_
rlabel metal2 7498 10812 7498 10812 0 _034_
rlabel metal2 7590 11084 7590 11084 0 _035_
rlabel metal1 7222 13328 7222 13328 0 _036_
rlabel metal2 7774 13940 7774 13940 0 _037_
rlabel metal1 8096 14042 8096 14042 0 _038_
rlabel metal1 7590 13362 7590 13362 0 _039_
rlabel metal1 7820 10642 7820 10642 0 _040_
rlabel metal1 8372 9622 8372 9622 0 _041_
rlabel metal2 8234 10234 8234 10234 0 _042_
rlabel metal1 8418 8976 8418 8976 0 _043_
rlabel metal1 7590 8908 7590 8908 0 _044_
rlabel metal1 7866 9520 7866 9520 0 _045_
rlabel metal1 8556 12206 8556 12206 0 _046_
rlabel metal1 8188 12206 8188 12206 0 _047_
rlabel metal1 8832 12138 8832 12138 0 _048_
rlabel metal2 8878 10982 8878 10982 0 _049_
rlabel metal1 8556 9350 8556 9350 0 _050_
rlabel metal2 5014 9146 5014 9146 0 _051_
rlabel metal2 927 17340 927 17340 0 io_in[0]
rlabel metal2 2399 17340 2399 17340 0 io_in[1]
rlabel metal1 4232 15470 4232 15470 0 io_in[2]
rlabel metal2 5382 16405 5382 16405 0 io_in[3]
rlabel metal1 6762 15470 6762 15470 0 io_in[4]
rlabel metal1 8372 15538 8372 15538 0 io_in[5]
rlabel metal1 9476 15538 9476 15538 0 io_in[6]
rlabel metal1 10718 14994 10718 14994 0 io_in[7]
rlabel metal2 782 1520 782 1520 0 io_out[0]
rlabel metal2 2254 1520 2254 1520 0 io_out[1]
rlabel metal2 3726 959 3726 959 0 io_out[2]
rlabel metal2 5198 1520 5198 1520 0 io_out[3]
rlabel metal2 6670 1520 6670 1520 0 io_out[4]
rlabel metal2 8142 1520 8142 1520 0 io_out[5]
rlabel metal2 9614 1520 9614 1520 0 io_out[6]
rlabel metal2 11086 1792 11086 1792 0 io_out[7]
rlabel metal1 2116 13294 2116 13294 0 net1
rlabel metal1 2668 12614 2668 12614 0 net10
rlabel metal2 4278 6154 4278 6154 0 net11
rlabel metal1 5198 8806 5198 8806 0 net12
rlabel metal1 6486 9010 6486 9010 0 net13
rlabel metal1 8096 2414 8096 2414 0 net14
rlabel metal1 9844 2414 9844 2414 0 net15
rlabel metal1 9660 9350 9660 9350 0 net16
rlabel metal1 2116 13906 2116 13906 0 net2
rlabel metal1 7682 13906 7682 13906 0 net3
rlabel metal1 8050 13872 8050 13872 0 net4
rlabel metal1 2530 13328 2530 13328 0 net5
rlabel metal1 5934 15130 5934 15130 0 net6
rlabel metal1 4922 12206 4922 12206 0 net7
rlabel metal1 7958 13940 7958 13940 0 net8
rlabel metal1 2484 2482 2484 2482 0 net9
<< properties >>
string FIXED_BBOX 0 0 12000 18000
<< end >>
