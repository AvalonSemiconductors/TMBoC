magic
tech sky130B
magscale 1 2
timestamp 1683540660
<< viali >>
rect 3985 19465 4019 19499
rect 17601 19465 17635 19499
rect 18521 19465 18555 19499
rect 11069 19397 11103 19431
rect 14749 19397 14783 19431
rect 17769 19397 17803 19431
rect 17969 19397 18003 19431
rect 19625 19397 19659 19431
rect 5098 19329 5132 19363
rect 5365 19329 5399 19363
rect 8217 19329 8251 19363
rect 10885 19329 10919 19363
rect 11805 19329 11839 19363
rect 12072 19329 12106 19363
rect 14657 19329 14691 19363
rect 14841 19329 14875 19363
rect 16957 19329 16991 19363
rect 18705 19329 18739 19363
rect 8033 19261 8067 19295
rect 19441 19261 19475 19295
rect 13185 19193 13219 19227
rect 17049 19125 17083 19159
rect 17785 19125 17819 19159
rect 2973 18921 3007 18955
rect 10701 18921 10735 18955
rect 14841 18921 14875 18955
rect 17049 18921 17083 18955
rect 17693 18853 17727 18887
rect 15301 18785 15335 18819
rect 15485 18785 15519 18819
rect 17233 18785 17267 18819
rect 2513 18717 2547 18751
rect 5733 18717 5767 18751
rect 8217 18717 8251 18751
rect 9321 18717 9355 18751
rect 11805 18717 11839 18751
rect 16957 18717 16991 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18153 18717 18187 18751
rect 18337 18717 18371 18751
rect 2329 18649 2363 18683
rect 3157 18649 3191 18683
rect 3341 18649 3375 18683
rect 5978 18649 6012 18683
rect 7941 18649 7975 18683
rect 9588 18649 9622 18683
rect 12072 18649 12106 18683
rect 17233 18649 17267 18683
rect 2145 18581 2179 18615
rect 7113 18581 7147 18615
rect 13185 18581 13219 18615
rect 15209 18581 15243 18615
rect 2237 18377 2271 18411
rect 3801 18377 3835 18411
rect 9321 18377 9355 18411
rect 15761 18377 15795 18411
rect 15853 18377 15887 18411
rect 18061 18377 18095 18411
rect 4914 18309 4948 18343
rect 7113 18309 7147 18343
rect 7297 18309 7331 18343
rect 7481 18309 7515 18343
rect 8186 18309 8220 18343
rect 16037 18309 16071 18343
rect 17141 18309 17175 18343
rect 17877 18309 17911 18343
rect 2421 18241 2455 18275
rect 2605 18241 2639 18275
rect 12256 18241 12290 18275
rect 14749 18241 14783 18275
rect 15669 18241 15703 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 17693 18241 17727 18275
rect 5181 18173 5215 18207
rect 7941 18173 7975 18207
rect 11989 18173 12023 18207
rect 14933 18173 14967 18207
rect 17049 18173 17083 18207
rect 13369 18037 13403 18071
rect 14565 18037 14599 18071
rect 15485 18037 15519 18071
rect 16865 18037 16899 18071
rect 3985 17833 4019 17867
rect 7021 17833 7055 17867
rect 10977 17833 11011 17867
rect 15117 17833 15151 17867
rect 17509 17833 17543 17867
rect 15209 17765 15243 17799
rect 2145 17629 2179 17663
rect 2329 17629 2363 17663
rect 5365 17629 5399 17663
rect 8401 17629 8435 17663
rect 9597 17629 9631 17663
rect 14933 17629 14967 17663
rect 15301 17629 15335 17663
rect 17417 17629 17451 17663
rect 17601 17629 17635 17663
rect 5098 17561 5132 17595
rect 8156 17561 8190 17595
rect 9864 17561 9898 17595
rect 2513 17493 2547 17527
rect 15025 17493 15059 17527
rect 2421 17289 2455 17323
rect 15761 17289 15795 17323
rect 17325 17221 17359 17255
rect 2237 17153 2271 17187
rect 2881 17153 2915 17187
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 7674 17153 7708 17187
rect 9137 17153 9171 17187
rect 9404 17153 9438 17187
rect 12081 17153 12115 17187
rect 12348 17153 12382 17187
rect 15025 17153 15059 17187
rect 15209 17153 15243 17187
rect 15669 17153 15703 17187
rect 15853 17153 15887 17187
rect 17141 17153 17175 17187
rect 17417 17153 17451 17187
rect 2053 17085 2087 17119
rect 7941 17085 7975 17119
rect 14841 17085 14875 17119
rect 6561 17017 6595 17051
rect 10517 16949 10551 16983
rect 13461 16949 13495 16983
rect 17141 16949 17175 16983
rect 3985 16745 4019 16779
rect 15853 16745 15887 16779
rect 16681 16745 16715 16779
rect 15301 16677 15335 16711
rect 16773 16677 16807 16711
rect 10885 16609 10919 16643
rect 14933 16609 14967 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 2053 16541 2087 16575
rect 2145 16541 2179 16575
rect 5365 16541 5399 16575
rect 15117 16541 15151 16575
rect 16037 16541 16071 16575
rect 16865 16541 16899 16575
rect 17417 16541 17451 16575
rect 18705 16541 18739 16575
rect 18889 16541 18923 16575
rect 19441 16541 19475 16575
rect 19625 16541 19659 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 1869 16473 1903 16507
rect 5098 16473 5132 16507
rect 11152 16473 11186 16507
rect 16589 16473 16623 16507
rect 17785 16473 17819 16507
rect 18797 16473 18831 16507
rect 1967 16405 2001 16439
rect 12265 16405 12299 16439
rect 20085 16405 20119 16439
rect 2329 16201 2363 16235
rect 16129 16201 16163 16235
rect 17233 16201 17267 16235
rect 17509 16201 17543 16235
rect 19625 16201 19659 16235
rect 5006 16133 5040 16167
rect 9496 16133 9530 16167
rect 17141 16133 17175 16167
rect 2145 16065 2179 16099
rect 7674 16065 7708 16099
rect 7941 16065 7975 16099
rect 9229 16065 9263 16099
rect 12256 16065 12290 16099
rect 14565 16065 14599 16099
rect 14841 16065 14875 16099
rect 15025 16065 15059 16099
rect 16037 16065 16071 16099
rect 16313 16065 16347 16099
rect 17325 16065 17359 16099
rect 19441 16065 19475 16099
rect 1869 15997 1903 16031
rect 5273 15997 5307 16031
rect 11989 15997 12023 16031
rect 16957 15997 16991 16031
rect 19257 15997 19291 16031
rect 1961 15929 1995 15963
rect 14749 15929 14783 15963
rect 14933 15929 14967 15963
rect 16313 15929 16347 15963
rect 3893 15861 3927 15895
rect 6561 15861 6595 15895
rect 10609 15861 10643 15895
rect 13369 15861 13403 15895
rect 15301 15861 15335 15895
rect 2513 15657 2547 15691
rect 5733 15657 5767 15691
rect 17141 15657 17175 15691
rect 17325 15657 17359 15691
rect 19993 15657 20027 15691
rect 19441 15521 19475 15555
rect 2145 15453 2179 15487
rect 2329 15453 2363 15487
rect 18153 15453 18187 15487
rect 7021 15385 7055 15419
rect 10425 15385 10459 15419
rect 17309 15385 17343 15419
rect 17509 15385 17543 15419
rect 19809 15385 19843 15419
rect 11897 15317 11931 15351
rect 18061 15317 18095 15351
rect 19625 15317 19659 15351
rect 19717 15317 19751 15351
rect 9965 15113 9999 15147
rect 13277 15113 13311 15147
rect 19149 15113 19183 15147
rect 7012 15045 7046 15079
rect 8677 15045 8711 15079
rect 17969 15045 18003 15079
rect 19349 15045 19383 15079
rect 2237 14977 2271 15011
rect 12164 14977 12198 15011
rect 14933 14977 14967 15011
rect 15209 14977 15243 15011
rect 15945 14977 15979 15011
rect 17693 14977 17727 15011
rect 19993 14977 20027 15011
rect 1961 14909 1995 14943
rect 6745 14909 6779 14943
rect 11897 14909 11931 14943
rect 15761 14909 15795 14943
rect 20177 14909 20211 14943
rect 15025 14841 15059 14875
rect 15117 14841 15151 14875
rect 16129 14841 16163 14875
rect 2053 14773 2087 14807
rect 2421 14773 2455 14807
rect 8125 14773 8159 14807
rect 14749 14773 14783 14807
rect 18981 14773 19015 14807
rect 19165 14773 19199 14807
rect 19809 14773 19843 14807
rect 1869 14569 1903 14603
rect 6009 14569 6043 14603
rect 14933 14569 14967 14603
rect 16773 14569 16807 14603
rect 19625 14569 19659 14603
rect 15117 14501 15151 14535
rect 15393 14433 15427 14467
rect 19993 14433 20027 14467
rect 2145 14365 2179 14399
rect 5365 14365 5399 14399
rect 7389 14365 7423 14399
rect 9689 14365 9723 14399
rect 17049 14365 17083 14399
rect 17141 14365 17175 14399
rect 17233 14365 17267 14399
rect 17417 14365 17451 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 1869 14297 1903 14331
rect 5098 14297 5132 14331
rect 7122 14297 7156 14331
rect 9956 14297 9990 14331
rect 2053 14229 2087 14263
rect 3985 14229 4019 14263
rect 11069 14229 11103 14263
rect 17877 14229 17911 14263
rect 18245 14229 18279 14263
rect 19441 14229 19475 14263
rect 19625 14229 19659 14263
rect 9045 14025 9079 14059
rect 11069 14025 11103 14059
rect 13185 14025 13219 14059
rect 19717 14025 19751 14059
rect 17141 13957 17175 13991
rect 18705 13957 18739 13991
rect 2329 13889 2363 13923
rect 2513 13889 2547 13923
rect 7932 13889 7966 13923
rect 12072 13889 12106 13923
rect 17509 13889 17543 13923
rect 18521 13889 18555 13923
rect 19165 13889 19199 13923
rect 19349 13889 19383 13923
rect 19441 13889 19475 13923
rect 19533 13889 19567 13923
rect 2145 13821 2179 13855
rect 5365 13821 5399 13855
rect 5641 13821 5675 13855
rect 7665 13821 7699 13855
rect 9505 13821 9539 13855
rect 9781 13821 9815 13855
rect 11805 13821 11839 13855
rect 18337 13821 18371 13855
rect 16957 13753 16991 13787
rect 4077 13685 4111 13719
rect 17141 13685 17175 13719
rect 3985 13481 4019 13515
rect 15025 13481 15059 13515
rect 2329 13413 2363 13447
rect 1869 13345 1903 13379
rect 2789 13345 2823 13379
rect 7941 13345 7975 13379
rect 1961 13277 1995 13311
rect 2145 13277 2179 13311
rect 2973 13277 3007 13311
rect 5365 13277 5399 13311
rect 7674 13277 7708 13311
rect 11805 13277 11839 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 17141 13277 17175 13311
rect 17417 13277 17451 13311
rect 17601 13277 17635 13311
rect 19625 13277 19659 13311
rect 3157 13209 3191 13243
rect 5098 13209 5132 13243
rect 12072 13209 12106 13243
rect 6561 13141 6595 13175
rect 13185 13141 13219 13175
rect 15577 13141 15611 13175
rect 16957 13141 16991 13175
rect 19717 13141 19751 13175
rect 1967 12937 2001 12971
rect 17877 12937 17911 12971
rect 1869 12869 1903 12903
rect 2053 12869 2087 12903
rect 6828 12869 6862 12903
rect 12072 12869 12106 12903
rect 19257 12869 19291 12903
rect 19441 12869 19475 12903
rect 19901 12869 19935 12903
rect 2145 12801 2179 12835
rect 14749 12801 14783 12835
rect 17049 12801 17083 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 17969 12801 18003 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 6561 12733 6595 12767
rect 11805 12733 11839 12767
rect 14841 12733 14875 12767
rect 15117 12733 15151 12767
rect 19901 12733 19935 12767
rect 19441 12665 19475 12699
rect 7941 12597 7975 12631
rect 13185 12597 13219 12631
rect 16865 12597 16899 12631
rect 20085 12597 20119 12631
rect 11161 12393 11195 12427
rect 15301 12393 15335 12427
rect 19625 12393 19659 12427
rect 15117 12325 15151 12359
rect 19441 12325 19475 12359
rect 5641 12257 5675 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 2789 12189 2823 12223
rect 2973 12189 3007 12223
rect 5365 12189 5399 12223
rect 9781 12189 9815 12223
rect 16405 12189 16439 12223
rect 16957 12189 16991 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 18337 12189 18371 12223
rect 19993 12189 20027 12223
rect 2881 12121 2915 12155
rect 10048 12121 10082 12155
rect 14841 12121 14875 12155
rect 17233 12121 17267 12155
rect 2329 12053 2363 12087
rect 4077 12053 4111 12087
rect 16313 12053 16347 12087
rect 17509 12053 17543 12087
rect 18061 12053 18095 12087
rect 19625 12053 19659 12087
rect 2329 11849 2363 11883
rect 13277 11849 13311 11883
rect 17417 11849 17451 11883
rect 17877 11849 17911 11883
rect 19349 11849 19383 11883
rect 19717 11849 19751 11883
rect 2145 11713 2179 11747
rect 5273 11713 5307 11747
rect 5549 11713 5583 11747
rect 6929 11713 6963 11747
rect 7196 11713 7230 11747
rect 8769 11713 8803 11747
rect 12164 11713 12198 11747
rect 17049 11713 17083 11747
rect 17141 11713 17175 11747
rect 17233 11713 17267 11747
rect 18061 11713 18095 11747
rect 18245 11713 18279 11747
rect 19257 11713 19291 11747
rect 19533 11713 19567 11747
rect 1961 11645 1995 11679
rect 3893 11645 3927 11679
rect 9045 11645 9079 11679
rect 11897 11645 11931 11679
rect 15301 11645 15335 11679
rect 15393 11577 15427 11611
rect 15485 11577 15519 11611
rect 15853 11577 15887 11611
rect 8309 11509 8343 11543
rect 10149 11509 10183 11543
rect 15025 11509 15059 11543
rect 18061 11509 18095 11543
rect 15301 11305 15335 11339
rect 16865 11305 16899 11339
rect 18797 11305 18831 11339
rect 19625 11305 19659 11339
rect 4077 11237 4111 11271
rect 10517 11237 10551 11271
rect 13185 11237 13219 11271
rect 15209 11237 15243 11271
rect 17509 11169 17543 11203
rect 1869 11101 1903 11135
rect 2053 11101 2087 11135
rect 5457 11101 5491 11135
rect 6469 11101 6503 11135
rect 9137 11101 9171 11135
rect 11805 11101 11839 11135
rect 17325 11101 17359 11135
rect 18705 11101 18739 11135
rect 18889 11101 18923 11135
rect 19993 11101 20027 11135
rect 1961 11033 1995 11067
rect 5190 11033 5224 11067
rect 6736 11033 6770 11067
rect 9382 11033 9416 11067
rect 12072 11033 12106 11067
rect 14841 11033 14875 11067
rect 19625 11033 19659 11067
rect 7849 10965 7883 10999
rect 17233 10965 17267 10999
rect 19441 10965 19475 10999
rect 1777 10761 1811 10795
rect 17877 10761 17911 10795
rect 19349 10761 19383 10795
rect 3801 10693 3835 10727
rect 7849 10693 7883 10727
rect 18045 10693 18079 10727
rect 18245 10693 18279 10727
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 2237 10625 2271 10659
rect 14105 10625 14139 10659
rect 14243 10625 14277 10659
rect 14565 10625 14599 10659
rect 15301 10625 15335 10659
rect 15577 10625 15611 10659
rect 17141 10625 17175 10659
rect 17417 10625 17451 10659
rect 19257 10625 19291 10659
rect 19441 10625 19475 10659
rect 1961 10557 1995 10591
rect 5181 10557 5215 10591
rect 5457 10557 5491 10591
rect 16865 10489 16899 10523
rect 9321 10421 9355 10455
rect 14381 10421 14415 10455
rect 14473 10421 14507 10455
rect 15025 10421 15059 10455
rect 15485 10421 15519 10455
rect 17233 10421 17267 10455
rect 18061 10421 18095 10455
rect 2053 10217 2087 10251
rect 17601 10217 17635 10251
rect 19993 10217 20027 10251
rect 13277 10149 13311 10183
rect 19441 10149 19475 10183
rect 10057 10081 10091 10115
rect 11897 10081 11931 10115
rect 14841 10081 14875 10115
rect 15301 10081 15335 10115
rect 17509 10081 17543 10115
rect 1777 10013 1811 10047
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 7021 10013 7055 10047
rect 14933 10013 14967 10047
rect 17233 10013 17267 10047
rect 18705 10013 18739 10047
rect 19717 10013 19751 10047
rect 5273 9945 5307 9979
rect 10324 9945 10358 9979
rect 12164 9945 12198 9979
rect 15209 9945 15243 9979
rect 11437 9877 11471 9911
rect 14657 9877 14691 9911
rect 18797 9877 18831 9911
rect 19625 9877 19659 9911
rect 19809 9877 19843 9911
rect 19625 9673 19659 9707
rect 20085 9673 20119 9707
rect 14841 9605 14875 9639
rect 19257 9605 19291 9639
rect 19457 9605 19491 9639
rect 4885 9537 4919 9571
rect 8329 9537 8363 9571
rect 9669 9537 9703 9571
rect 11897 9537 11931 9571
rect 12164 9537 12198 9571
rect 14105 9537 14139 9571
rect 14988 9537 15022 9571
rect 17233 9537 17267 9571
rect 17601 9537 17635 9571
rect 20085 9537 20119 9571
rect 20269 9537 20303 9571
rect 4629 9469 4663 9503
rect 8585 9469 8619 9503
rect 9413 9469 9447 9503
rect 14381 9469 14415 9503
rect 15209 9469 15243 9503
rect 17325 9469 17359 9503
rect 17693 9469 17727 9503
rect 6009 9401 6043 9435
rect 14289 9401 14323 9435
rect 15117 9401 15151 9435
rect 17877 9401 17911 9435
rect 7205 9333 7239 9367
rect 10793 9333 10827 9367
rect 13277 9333 13311 9367
rect 14197 9333 14231 9367
rect 15301 9333 15335 9367
rect 19441 9333 19475 9367
rect 8493 9129 8527 9163
rect 14565 9129 14599 9163
rect 19533 9129 19567 9163
rect 2145 8993 2179 9027
rect 3985 8993 4019 9027
rect 7941 8993 7975 9027
rect 14657 8993 14691 9027
rect 2421 8925 2455 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 14841 8925 14875 8959
rect 16957 8925 16991 8959
rect 17120 8925 17154 8959
rect 17233 8925 17267 8959
rect 17325 8925 17359 8959
rect 19441 8925 19475 8959
rect 19625 8925 19659 8959
rect 4252 8857 4286 8891
rect 7674 8857 7708 8891
rect 14565 8857 14599 8891
rect 1593 8789 1627 8823
rect 5365 8789 5399 8823
rect 6561 8789 6595 8823
rect 15025 8789 15059 8823
rect 17601 8789 17635 8823
rect 2513 8585 2547 8619
rect 4629 8585 4663 8619
rect 5273 8585 5307 8619
rect 12265 8585 12299 8619
rect 16957 8585 16991 8619
rect 19533 8585 19567 8619
rect 5917 8517 5951 8551
rect 6806 8517 6840 8551
rect 18061 8517 18095 8551
rect 19701 8517 19735 8551
rect 19901 8517 19935 8551
rect 2053 8449 2087 8483
rect 2329 8449 2363 8483
rect 4445 8449 4479 8483
rect 4629 8449 4663 8483
rect 5365 8449 5399 8483
rect 6009 8449 6043 8483
rect 6561 8449 6595 8483
rect 8401 8449 8435 8483
rect 12633 8449 12667 8483
rect 14565 8449 14599 8483
rect 14841 8449 14875 8483
rect 15025 8449 15059 8483
rect 17141 8449 17175 8483
rect 17877 8449 17911 8483
rect 18153 8449 18187 8483
rect 18889 8449 18923 8483
rect 19073 8449 19107 8483
rect 12541 8381 12575 8415
rect 15209 8381 15243 8415
rect 17417 8381 17451 8415
rect 2145 8313 2179 8347
rect 7941 8313 7975 8347
rect 17325 8313 17359 8347
rect 18981 8313 19015 8347
rect 8493 8245 8527 8279
rect 12633 8245 12667 8279
rect 17877 8245 17911 8279
rect 19717 8245 19751 8279
rect 2237 8041 2271 8075
rect 4721 8041 4755 8075
rect 7021 8041 7055 8075
rect 8401 8041 8435 8075
rect 9229 8041 9263 8075
rect 10701 8041 10735 8075
rect 12449 8041 12483 8075
rect 12633 8041 12667 8075
rect 13277 8041 13311 8075
rect 14657 8041 14691 8075
rect 15117 8041 15151 8075
rect 16497 8041 16531 8075
rect 17325 8041 17359 8075
rect 18889 8041 18923 8075
rect 19809 8041 19843 8075
rect 16589 7973 16623 8007
rect 17141 7973 17175 8007
rect 18705 7973 18739 8007
rect 4077 7905 4111 7939
rect 5181 7905 5215 7939
rect 9321 7905 9355 7939
rect 13369 7905 13403 7939
rect 14933 7905 14967 7939
rect 16405 7905 16439 7939
rect 18429 7905 18463 7939
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 4445 7837 4479 7871
rect 4537 7837 4571 7871
rect 5365 7837 5399 7871
rect 5641 7837 5675 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 8033 7837 8067 7871
rect 9413 7837 9447 7871
rect 10885 7837 10919 7871
rect 10977 7837 11011 7871
rect 11161 7837 11195 7871
rect 11253 7837 11287 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 15209 7837 15243 7871
rect 16681 7837 16715 7871
rect 19441 7837 19475 7871
rect 8217 7769 8251 7803
rect 9689 7769 9723 7803
rect 12265 7769 12299 7803
rect 12481 7769 12515 7803
rect 17309 7769 17343 7803
rect 17509 7769 17543 7803
rect 19625 7769 19659 7803
rect 2053 7701 2087 7735
rect 5549 7701 5583 7735
rect 9597 7701 9631 7735
rect 4905 7497 4939 7531
rect 5733 7497 5767 7531
rect 6837 7497 6871 7531
rect 7481 7497 7515 7531
rect 10057 7497 10091 7531
rect 12173 7497 12207 7531
rect 13369 7497 13403 7531
rect 13553 7497 13587 7531
rect 17509 7497 17543 7531
rect 9873 7429 9907 7463
rect 12357 7429 12391 7463
rect 15761 7429 15795 7463
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 5181 7361 5215 7395
rect 5733 7361 5767 7395
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 8309 7361 8343 7395
rect 8493 7361 8527 7395
rect 8585 7361 8619 7395
rect 10149 7361 10183 7395
rect 10793 7361 10827 7395
rect 12081 7361 12115 7395
rect 13550 7361 13584 7395
rect 14013 7361 14047 7395
rect 15117 7361 15151 7395
rect 15669 7361 15703 7395
rect 17049 7361 17083 7395
rect 17325 7361 17359 7395
rect 6837 7293 6871 7327
rect 14841 7293 14875 7327
rect 8401 7225 8435 7259
rect 9873 7225 9907 7259
rect 12357 7225 12391 7259
rect 14933 7225 14967 7259
rect 6653 7157 6687 7191
rect 8125 7157 8159 7191
rect 10701 7157 10735 7191
rect 13921 7157 13955 7191
rect 4537 6953 4571 6987
rect 4813 6953 4847 6987
rect 6377 6953 6411 6987
rect 12449 6953 12483 6987
rect 14749 6953 14783 6987
rect 2053 6817 2087 6851
rect 5917 6817 5951 6851
rect 13001 6817 13035 6851
rect 2237 6749 2271 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 6193 6749 6227 6783
rect 10793 6749 10827 6783
rect 10885 6749 10919 6783
rect 12633 6749 12667 6783
rect 14565 6749 14599 6783
rect 15209 6749 15243 6783
rect 16773 6749 16807 6783
rect 16866 6749 16900 6783
rect 10609 6681 10643 6715
rect 12725 6681 12759 6715
rect 17141 6681 17175 6715
rect 2421 6613 2455 6647
rect 10707 6613 10741 6647
rect 12817 6613 12851 6647
rect 10425 6409 10459 6443
rect 13553 6409 13587 6443
rect 7389 6341 7423 6375
rect 13277 6341 13311 6375
rect 13829 6341 13863 6375
rect 1869 6273 1903 6307
rect 2053 6273 2087 6307
rect 4353 6273 4387 6307
rect 4537 6273 4571 6307
rect 6837 6273 6871 6307
rect 7021 6273 7055 6307
rect 7757 6273 7791 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 10333 6273 10367 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 11989 6273 12023 6307
rect 13461 6273 13495 6307
rect 13645 6273 13679 6307
rect 15393 6273 15427 6307
rect 15669 6273 15703 6307
rect 2881 6205 2915 6239
rect 6561 6205 6595 6239
rect 7941 6205 7975 6239
rect 8953 6205 8987 6239
rect 11161 6205 11195 6239
rect 12265 6205 12299 6239
rect 14381 6205 14415 6239
rect 16037 6205 16071 6239
rect 17233 6205 17267 6239
rect 17601 6205 17635 6239
rect 17693 6205 17727 6239
rect 17785 6205 17819 6239
rect 14749 6137 14783 6171
rect 15485 6137 15519 6171
rect 4445 6069 4479 6103
rect 8677 6069 8711 6103
rect 11805 6069 11839 6103
rect 12173 6069 12207 6103
rect 14841 6069 14875 6103
rect 2053 5865 2087 5899
rect 5917 5865 5951 5899
rect 10517 5865 10551 5899
rect 12541 5865 12575 5899
rect 12725 5865 12759 5899
rect 14289 5865 14323 5899
rect 14473 5865 14507 5899
rect 5181 5797 5215 5831
rect 8401 5797 8435 5831
rect 10609 5797 10643 5831
rect 13553 5797 13587 5831
rect 17141 5797 17175 5831
rect 2329 5729 2363 5763
rect 2513 5729 2547 5763
rect 4721 5729 4755 5763
rect 6469 5729 6503 5763
rect 8309 5729 8343 5763
rect 10425 5729 10459 5763
rect 14565 5729 14599 5763
rect 15577 5729 15611 5763
rect 16037 5729 16071 5763
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 3249 5661 3283 5695
rect 4629 5661 4663 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 8217 5661 8251 5695
rect 8493 5661 8527 5695
rect 10701 5661 10735 5695
rect 13369 5661 13403 5695
rect 14657 5661 14691 5695
rect 16129 5661 16163 5695
rect 17141 5661 17175 5695
rect 17693 5661 17727 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 3065 5593 3099 5627
rect 4721 5593 4755 5627
rect 6653 5593 6687 5627
rect 7021 5593 7055 5627
rect 8033 5593 8067 5627
rect 12909 5593 12943 5627
rect 3433 5525 3467 5559
rect 6745 5525 6779 5559
rect 6837 5525 6871 5559
rect 12709 5525 12743 5559
rect 15761 5525 15795 5559
rect 2145 5321 2179 5355
rect 4813 5321 4847 5355
rect 6009 5321 6043 5355
rect 10885 5321 10919 5355
rect 17509 5321 17543 5355
rect 18797 5321 18831 5355
rect 5641 5253 5675 5287
rect 5825 5253 5859 5287
rect 17601 5253 17635 5287
rect 18153 5253 18187 5287
rect 2053 5185 2087 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4997 5185 5031 5219
rect 7205 5185 7239 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 8585 5185 8619 5219
rect 9137 5185 9171 5219
rect 10149 5185 10183 5219
rect 10333 5185 10367 5219
rect 10885 5185 10919 5219
rect 11897 5185 11931 5219
rect 12081 5185 12115 5219
rect 13277 5185 13311 5219
rect 14105 5185 14139 5219
rect 14197 5185 14231 5219
rect 15025 5185 15059 5219
rect 15209 5185 15243 5219
rect 15485 5185 15519 5219
rect 17417 5185 17451 5219
rect 18300 5185 18334 5219
rect 4353 5117 4387 5151
rect 5181 5117 5215 5151
rect 8309 5117 8343 5151
rect 12357 5117 12391 5151
rect 12449 5117 12483 5151
rect 13001 5117 13035 5151
rect 13185 5117 13219 5151
rect 13369 5117 13403 5151
rect 13461 5117 13495 5151
rect 16865 5117 16899 5151
rect 17049 5117 17083 5151
rect 18521 5117 18555 5151
rect 9229 5049 9263 5083
rect 15393 5049 15427 5083
rect 18429 5049 18463 5083
rect 7757 4981 7791 5015
rect 6193 4777 6227 4811
rect 13277 4777 13311 4811
rect 15209 4777 15243 4811
rect 4353 4641 4387 4675
rect 7941 4641 7975 4675
rect 8125 4641 8159 4675
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 8309 4573 8343 4607
rect 8585 4573 8619 4607
rect 13185 4573 13219 4607
rect 13369 4573 13403 4607
rect 15209 4573 15243 4607
rect 15393 4573 15427 4607
rect 4353 4097 4387 4131
rect 5365 4097 5399 4131
rect 2145 2397 2179 2431
rect 4813 2397 4847 2431
rect 7481 2397 7515 2431
rect 9689 2397 9723 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17693 2397 17727 2431
rect 19901 2397 19935 2431
rect 1869 2329 1903 2363
rect 4537 2329 4571 2363
rect 7205 2329 7239 2363
rect 9965 2329 9999 2363
rect 12633 2329 12667 2363
rect 15301 2329 15335 2363
rect 17969 2329 18003 2363
rect 20177 2329 20211 2363
<< metal1 >>
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 14642 19700 14648 19712
rect 8076 19672 14648 19700
rect 8076 19660 8082 19672
rect 14642 19660 14648 19672
rect 14700 19700 14706 19712
rect 15654 19700 15660 19712
rect 14700 19672 15660 19700
rect 14700 19660 14706 19672
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 1104 19610 21043 19632
rect 1104 19558 5894 19610
rect 5946 19558 5958 19610
rect 6010 19558 6022 19610
rect 6074 19558 6086 19610
rect 6138 19558 6150 19610
rect 6202 19558 10839 19610
rect 10891 19558 10903 19610
rect 10955 19558 10967 19610
rect 11019 19558 11031 19610
rect 11083 19558 11095 19610
rect 11147 19558 15784 19610
rect 15836 19558 15848 19610
rect 15900 19558 15912 19610
rect 15964 19558 15976 19610
rect 16028 19558 16040 19610
rect 16092 19558 20729 19610
rect 20781 19558 20793 19610
rect 20845 19558 20857 19610
rect 20909 19558 20921 19610
rect 20973 19558 20985 19610
rect 21037 19558 21043 19610
rect 1104 19536 21043 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 2832 19468 3985 19496
rect 2832 19456 2838 19468
rect 3973 19465 3985 19468
rect 4019 19465 4031 19499
rect 3973 19459 4031 19465
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 17589 19499 17647 19505
rect 17589 19496 17601 19499
rect 13780 19468 17601 19496
rect 13780 19456 13786 19468
rect 17589 19465 17601 19468
rect 17635 19465 17647 19499
rect 18509 19499 18567 19505
rect 18509 19496 18521 19499
rect 17589 19459 17647 19465
rect 17696 19468 18521 19496
rect 11057 19431 11115 19437
rect 11057 19397 11069 19431
rect 11103 19428 11115 19431
rect 11238 19428 11244 19440
rect 11103 19400 11244 19428
rect 11103 19397 11115 19400
rect 11057 19391 11115 19397
rect 11238 19388 11244 19400
rect 11296 19388 11302 19440
rect 14737 19431 14795 19437
rect 14737 19428 14749 19431
rect 12406 19400 14749 19428
rect 4154 19320 4160 19372
rect 4212 19360 4218 19372
rect 5086 19363 5144 19369
rect 5086 19360 5098 19363
rect 4212 19332 5098 19360
rect 4212 19320 4218 19332
rect 5086 19329 5098 19332
rect 5132 19329 5144 19363
rect 5086 19323 5144 19329
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 5316 19332 5365 19360
rect 5316 19320 5322 19332
rect 5353 19329 5365 19332
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 8251 19332 10885 19360
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 10873 19329 10885 19332
rect 10919 19329 10931 19363
rect 10873 19323 10931 19329
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 11882 19360 11888 19372
rect 11839 19332 11888 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12060 19363 12118 19369
rect 12060 19329 12072 19363
rect 12106 19360 12118 19363
rect 12406 19360 12434 19400
rect 14737 19397 14749 19400
rect 14783 19397 14795 19431
rect 14737 19391 14795 19397
rect 17126 19388 17132 19440
rect 17184 19428 17190 19440
rect 17696 19428 17724 19468
rect 18509 19465 18521 19468
rect 18555 19465 18567 19499
rect 18509 19459 18567 19465
rect 17770 19437 17776 19440
rect 17184 19400 17724 19428
rect 17757 19431 17776 19437
rect 17184 19388 17190 19400
rect 17757 19397 17769 19431
rect 17757 19391 17776 19397
rect 17770 19388 17776 19391
rect 17828 19388 17834 19440
rect 17954 19388 17960 19440
rect 18012 19388 18018 19440
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 19613 19431 19671 19437
rect 19613 19428 19625 19431
rect 18288 19400 19625 19428
rect 18288 19388 18294 19400
rect 19613 19397 19625 19400
rect 19659 19397 19671 19431
rect 19613 19391 19671 19397
rect 12106 19332 12434 19360
rect 13188 19332 14596 19360
rect 12106 19329 12118 19332
rect 12060 19323 12118 19329
rect 8018 19252 8024 19304
rect 8076 19252 8082 19304
rect 13188 19233 13216 19332
rect 14568 19292 14596 19332
rect 14642 19320 14648 19372
rect 14700 19320 14706 19372
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 16942 19320 16948 19372
rect 17000 19320 17006 19372
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 15286 19292 15292 19304
rect 14568 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 18708 19292 18736 19323
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 18708 19264 19441 19292
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 13173 19227 13231 19233
rect 13173 19193 13185 19227
rect 13219 19193 13231 19227
rect 13173 19187 13231 19193
rect 17034 19116 17040 19168
rect 17092 19116 17098 19168
rect 17773 19159 17831 19165
rect 17773 19125 17785 19159
rect 17819 19156 17831 19159
rect 18046 19156 18052 19168
rect 17819 19128 18052 19156
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 1104 19066 20884 19088
rect 1104 19014 3422 19066
rect 3474 19014 3486 19066
rect 3538 19014 3550 19066
rect 3602 19014 3614 19066
rect 3666 19014 3678 19066
rect 3730 19014 8367 19066
rect 8419 19014 8431 19066
rect 8483 19014 8495 19066
rect 8547 19014 8559 19066
rect 8611 19014 8623 19066
rect 8675 19014 13312 19066
rect 13364 19014 13376 19066
rect 13428 19014 13440 19066
rect 13492 19014 13504 19066
rect 13556 19014 13568 19066
rect 13620 19014 18257 19066
rect 18309 19014 18321 19066
rect 18373 19014 18385 19066
rect 18437 19014 18449 19066
rect 18501 19014 18513 19066
rect 18565 19014 20884 19066
rect 1104 18992 20884 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 4154 18952 4160 18964
rect 3007 18924 4160 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 10735 18924 14780 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 14752 18884 14780 18924
rect 14826 18912 14832 18964
rect 14884 18912 14890 18964
rect 16114 18952 16120 18964
rect 14936 18924 16120 18952
rect 14936 18884 14964 18924
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 17034 18912 17040 18964
rect 17092 18912 17098 18964
rect 17681 18887 17739 18893
rect 17681 18884 17693 18887
rect 14752 18856 14964 18884
rect 15028 18856 17693 18884
rect 14844 18828 14872 18856
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 2464 18788 5856 18816
rect 2464 18776 2470 18788
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18748 2559 18751
rect 4062 18748 4068 18760
rect 2547 18720 4068 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 5258 18708 5264 18760
rect 5316 18748 5322 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5316 18720 5733 18748
rect 5316 18708 5322 18720
rect 5721 18717 5733 18720
rect 5767 18717 5779 18751
rect 5828 18748 5856 18788
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 8018 18748 8024 18760
rect 5828 18720 8024 18748
rect 5721 18711 5779 18717
rect 8018 18708 8024 18720
rect 8076 18748 8082 18760
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 8076 18720 8217 18748
rect 8076 18708 8082 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 9272 18720 9321 18748
rect 9272 18708 9278 18720
rect 9309 18717 9321 18720
rect 9355 18748 9367 18751
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 9355 18720 11805 18748
rect 9355 18717 9367 18720
rect 9309 18711 9367 18717
rect 11793 18717 11805 18720
rect 11839 18748 11851 18751
rect 11882 18748 11888 18760
rect 11839 18720 11888 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 15028 18748 15056 18856
rect 17681 18853 17693 18856
rect 17727 18853 17739 18887
rect 17681 18847 17739 18853
rect 15286 18776 15292 18828
rect 15344 18776 15350 18828
rect 15470 18776 15476 18828
rect 15528 18776 15534 18828
rect 17126 18816 17132 18828
rect 16960 18788 17132 18816
rect 16960 18757 16988 18788
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17770 18816 17776 18828
rect 17276 18788 17776 18816
rect 17276 18776 17282 18788
rect 17770 18776 17776 18788
rect 17828 18816 17834 18828
rect 17828 18788 18092 18816
rect 17828 18776 17834 18788
rect 11992 18720 15056 18748
rect 16945 18751 17003 18757
rect 2317 18683 2375 18689
rect 2317 18649 2329 18683
rect 2363 18680 2375 18683
rect 3142 18680 3148 18692
rect 2363 18652 3148 18680
rect 2363 18649 2375 18652
rect 2317 18643 2375 18649
rect 3142 18640 3148 18652
rect 3200 18640 3206 18692
rect 3329 18683 3387 18689
rect 3329 18649 3341 18683
rect 3375 18680 3387 18683
rect 3786 18680 3792 18692
rect 3375 18652 3792 18680
rect 3375 18649 3387 18652
rect 3329 18643 3387 18649
rect 3786 18640 3792 18652
rect 3844 18640 3850 18692
rect 5966 18683 6024 18689
rect 5966 18680 5978 18683
rect 4172 18652 5978 18680
rect 2130 18572 2136 18624
rect 2188 18572 2194 18624
rect 2222 18572 2228 18624
rect 2280 18612 2286 18624
rect 4172 18612 4200 18652
rect 5966 18649 5978 18652
rect 6012 18649 6024 18683
rect 5966 18643 6024 18649
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 7929 18683 7987 18689
rect 7929 18680 7941 18683
rect 7340 18652 7941 18680
rect 7340 18640 7346 18652
rect 7929 18649 7941 18652
rect 7975 18649 7987 18683
rect 7929 18643 7987 18649
rect 9576 18683 9634 18689
rect 9576 18649 9588 18683
rect 9622 18680 9634 18683
rect 11992 18680 12020 18720
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 18064 18757 18092 18788
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17092 18720 17969 18748
rect 17092 18708 17098 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 9622 18652 12020 18680
rect 12060 18683 12118 18689
rect 9622 18649 9634 18652
rect 9576 18643 9634 18649
rect 12060 18649 12072 18683
rect 12106 18680 12118 18683
rect 13722 18680 13728 18692
rect 12106 18652 13728 18680
rect 12106 18649 12118 18652
rect 12060 18643 12118 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 14918 18640 14924 18692
rect 14976 18680 14982 18692
rect 17221 18683 17279 18689
rect 14976 18652 17172 18680
rect 14976 18640 14982 18652
rect 2280 18584 4200 18612
rect 2280 18572 2286 18584
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18612 13231 18615
rect 15010 18612 15016 18624
rect 13219 18584 15016 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15194 18572 15200 18624
rect 15252 18572 15258 18624
rect 17144 18612 17172 18652
rect 17221 18649 17233 18683
rect 17267 18680 17279 18683
rect 18156 18680 18184 18711
rect 17267 18652 18184 18680
rect 17267 18649 17279 18652
rect 17221 18643 17279 18649
rect 17954 18612 17960 18624
rect 17144 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18612 18018 18624
rect 18340 18612 18368 18711
rect 19242 18612 19248 18624
rect 18012 18584 19248 18612
rect 18012 18572 18018 18584
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 1104 18522 21043 18544
rect 1104 18470 5894 18522
rect 5946 18470 5958 18522
rect 6010 18470 6022 18522
rect 6074 18470 6086 18522
rect 6138 18470 6150 18522
rect 6202 18470 10839 18522
rect 10891 18470 10903 18522
rect 10955 18470 10967 18522
rect 11019 18470 11031 18522
rect 11083 18470 11095 18522
rect 11147 18470 15784 18522
rect 15836 18470 15848 18522
rect 15900 18470 15912 18522
rect 15964 18470 15976 18522
rect 16028 18470 16040 18522
rect 16092 18470 20729 18522
rect 20781 18470 20793 18522
rect 20845 18470 20857 18522
rect 20909 18470 20921 18522
rect 20973 18470 20985 18522
rect 21037 18470 21043 18522
rect 1104 18448 21043 18470
rect 2222 18368 2228 18420
rect 2280 18368 2286 18420
rect 3786 18368 3792 18420
rect 3844 18368 3850 18420
rect 9309 18411 9367 18417
rect 9309 18377 9321 18411
rect 9355 18377 9367 18411
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 9309 18371 9367 18377
rect 15580 18380 15761 18408
rect 2130 18300 2136 18352
rect 2188 18340 2194 18352
rect 4902 18343 4960 18349
rect 4902 18340 4914 18343
rect 2188 18312 4914 18340
rect 2188 18300 2194 18312
rect 4902 18309 4914 18312
rect 4948 18309 4960 18343
rect 4902 18303 4960 18309
rect 7098 18300 7104 18352
rect 7156 18300 7162 18352
rect 7282 18300 7288 18352
rect 7340 18300 7346 18352
rect 7469 18343 7527 18349
rect 7469 18309 7481 18343
rect 7515 18340 7527 18343
rect 8174 18343 8232 18349
rect 8174 18340 8186 18343
rect 7515 18312 8186 18340
rect 7515 18309 7527 18312
rect 7469 18303 7527 18309
rect 8174 18309 8186 18312
rect 8220 18309 8232 18343
rect 9324 18340 9352 18371
rect 9324 18312 12434 18340
rect 8174 18303 8232 18309
rect 2406 18232 2412 18284
rect 2464 18232 2470 18284
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3878 18272 3884 18284
rect 2639 18244 3884 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 7300 18272 7328 18300
rect 12250 18281 12256 18284
rect 3988 18244 7328 18272
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3988 18204 4016 18244
rect 12244 18235 12256 18281
rect 12250 18232 12256 18235
rect 12308 18232 12314 18284
rect 12406 18272 12434 18312
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 15580 18340 15608 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 15749 18371 15807 18377
rect 15838 18368 15844 18420
rect 15896 18368 15902 18420
rect 18046 18368 18052 18420
rect 18104 18368 18110 18420
rect 15436 18312 15608 18340
rect 16025 18343 16083 18349
rect 15436 18300 15442 18312
rect 16025 18309 16037 18343
rect 16071 18340 16083 18343
rect 16114 18340 16120 18352
rect 16071 18312 16120 18340
rect 16071 18309 16083 18312
rect 16025 18303 16083 18309
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 17092 18312 17141 18340
rect 17092 18300 17098 18312
rect 17129 18309 17141 18312
rect 17175 18340 17187 18343
rect 17865 18343 17923 18349
rect 17865 18340 17877 18343
rect 17175 18312 17877 18340
rect 17175 18309 17187 18312
rect 17129 18303 17187 18309
rect 17865 18309 17877 18312
rect 17911 18309 17923 18343
rect 17865 18303 17923 18309
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 12406 18244 14749 18272
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 14737 18235 14795 18241
rect 15580 18244 15669 18272
rect 3200 18176 4016 18204
rect 5169 18207 5227 18213
rect 3200 18164 3206 18176
rect 5169 18173 5181 18207
rect 5215 18204 5227 18207
rect 5258 18204 5264 18216
rect 5215 18176 5264 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 7926 18164 7932 18216
rect 7984 18164 7990 18216
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 11940 18176 11989 18204
rect 11940 18164 11946 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 13630 18164 13636 18216
rect 13688 18204 13694 18216
rect 14918 18204 14924 18216
rect 13688 18176 14924 18204
rect 13688 18164 13694 18176
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 15580 18136 15608 18244
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16960 18244 17233 18272
rect 16114 18204 16120 18216
rect 15948 18176 16120 18204
rect 15948 18136 15976 18176
rect 16114 18164 16120 18176
rect 16172 18204 16178 18216
rect 16960 18204 16988 18244
rect 17221 18241 17233 18244
rect 17267 18272 17279 18275
rect 17586 18272 17592 18284
rect 17267 18244 17592 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17586 18232 17592 18244
rect 17644 18272 17650 18284
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 17644 18244 17693 18272
rect 17644 18232 17650 18244
rect 17681 18241 17693 18244
rect 17727 18241 17739 18275
rect 17681 18235 17739 18241
rect 16172 18176 16988 18204
rect 17037 18207 17095 18213
rect 16172 18164 16178 18176
rect 17037 18173 17049 18207
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 15580 18108 15976 18136
rect 16206 18096 16212 18148
rect 16264 18136 16270 18148
rect 16942 18136 16948 18148
rect 16264 18108 16948 18136
rect 16264 18096 16270 18108
rect 16942 18096 16948 18108
rect 17000 18136 17006 18148
rect 17052 18136 17080 18167
rect 17000 18108 17080 18136
rect 17000 18096 17006 18108
rect 13357 18071 13415 18077
rect 13357 18037 13369 18071
rect 13403 18068 13415 18071
rect 14366 18068 14372 18080
rect 13403 18040 14372 18068
rect 13403 18037 13415 18040
rect 13357 18031 13415 18037
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14550 18028 14556 18080
rect 14608 18028 14614 18080
rect 15470 18028 15476 18080
rect 15528 18028 15534 18080
rect 15562 18028 15568 18080
rect 15620 18068 15626 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 15620 18040 16865 18068
rect 15620 18028 15626 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 1104 17978 20884 18000
rect 1104 17926 3422 17978
rect 3474 17926 3486 17978
rect 3538 17926 3550 17978
rect 3602 17926 3614 17978
rect 3666 17926 3678 17978
rect 3730 17926 8367 17978
rect 8419 17926 8431 17978
rect 8483 17926 8495 17978
rect 8547 17926 8559 17978
rect 8611 17926 8623 17978
rect 8675 17926 13312 17978
rect 13364 17926 13376 17978
rect 13428 17926 13440 17978
rect 13492 17926 13504 17978
rect 13556 17926 13568 17978
rect 13620 17926 18257 17978
rect 18309 17926 18321 17978
rect 18373 17926 18385 17978
rect 18437 17926 18449 17978
rect 18501 17926 18513 17978
rect 18565 17926 20884 17978
rect 1104 17904 20884 17926
rect 3878 17824 3884 17876
rect 3936 17864 3942 17876
rect 3973 17867 4031 17873
rect 3973 17864 3985 17867
rect 3936 17836 3985 17864
rect 3936 17824 3942 17836
rect 3973 17833 3985 17836
rect 4019 17833 4031 17867
rect 3973 17827 4031 17833
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 7009 17867 7067 17873
rect 7009 17864 7021 17867
rect 4120 17836 7021 17864
rect 4120 17824 4126 17836
rect 7009 17833 7021 17836
rect 7055 17833 7067 17867
rect 7009 17827 7067 17833
rect 10962 17824 10968 17876
rect 11020 17824 11026 17876
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 15562 17864 15568 17876
rect 15151 17836 15568 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 15197 17799 15255 17805
rect 15197 17765 15209 17799
rect 15243 17796 15255 17799
rect 15746 17796 15752 17808
rect 15243 17768 15752 17796
rect 15243 17765 15255 17768
rect 15197 17759 15255 17765
rect 15580 17740 15608 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 15470 17728 15476 17740
rect 14936 17700 15476 17728
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 2133 17663 2191 17669
rect 2133 17660 2145 17663
rect 2096 17632 2145 17660
rect 2096 17620 2102 17632
rect 2133 17629 2145 17632
rect 2179 17629 2191 17663
rect 2133 17623 2191 17629
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2774 17660 2780 17672
rect 2363 17632 2780 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 5258 17620 5264 17672
rect 5316 17660 5322 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 5316 17632 5365 17660
rect 5316 17620 5322 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 8389 17663 8447 17669
rect 8389 17660 8401 17663
rect 5353 17623 5411 17629
rect 7944 17632 8401 17660
rect 7944 17604 7972 17632
rect 8389 17629 8401 17632
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9585 17663 9643 17669
rect 9585 17660 9597 17663
rect 9272 17632 9597 17660
rect 9272 17620 9278 17632
rect 9585 17629 9597 17632
rect 9631 17629 9643 17663
rect 14550 17660 14556 17672
rect 9585 17623 9643 17629
rect 9784 17632 14556 17660
rect 2406 17552 2412 17604
rect 2464 17592 2470 17604
rect 5086 17595 5144 17601
rect 5086 17592 5098 17595
rect 2464 17564 5098 17592
rect 2464 17552 2470 17564
rect 5086 17561 5098 17564
rect 5132 17561 5144 17595
rect 5086 17555 5144 17561
rect 7926 17552 7932 17604
rect 7984 17552 7990 17604
rect 8144 17595 8202 17601
rect 8144 17561 8156 17595
rect 8190 17592 8202 17595
rect 9784 17592 9812 17632
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 14936 17669 14964 17700
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15562 17688 15568 17740
rect 15620 17688 15626 17740
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 17126 17660 17132 17672
rect 15335 17632 17132 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 8190 17564 9812 17592
rect 9852 17595 9910 17601
rect 8190 17561 8202 17564
rect 8144 17555 8202 17561
rect 9852 17561 9864 17595
rect 9898 17592 9910 17595
rect 9898 17564 12434 17592
rect 9898 17561 9910 17564
rect 9852 17555 9910 17561
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 4982 17524 4988 17536
rect 2547 17496 4988 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 12406 17524 12434 17564
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 17034 17592 17040 17604
rect 15528 17564 17040 17592
rect 15528 17552 15534 17564
rect 17034 17552 17040 17564
rect 17092 17592 17098 17604
rect 17420 17592 17448 17623
rect 17586 17620 17592 17672
rect 17644 17620 17650 17672
rect 17092 17564 17448 17592
rect 17092 17552 17098 17564
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 12406 17496 15025 17524
rect 15013 17493 15025 17496
rect 15059 17493 15071 17527
rect 15013 17487 15071 17493
rect 1104 17434 21043 17456
rect 1104 17382 5894 17434
rect 5946 17382 5958 17434
rect 6010 17382 6022 17434
rect 6074 17382 6086 17434
rect 6138 17382 6150 17434
rect 6202 17382 10839 17434
rect 10891 17382 10903 17434
rect 10955 17382 10967 17434
rect 11019 17382 11031 17434
rect 11083 17382 11095 17434
rect 11147 17382 15784 17434
rect 15836 17382 15848 17434
rect 15900 17382 15912 17434
rect 15964 17382 15976 17434
rect 16028 17382 16040 17434
rect 16092 17382 20729 17434
rect 20781 17382 20793 17434
rect 20845 17382 20857 17434
rect 20909 17382 20921 17434
rect 20973 17382 20985 17434
rect 21037 17382 21043 17434
rect 1104 17360 21043 17382
rect 2406 17280 2412 17332
rect 2464 17280 2470 17332
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 15252 17292 15761 17320
rect 15252 17280 15258 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 2038 17212 2044 17264
rect 2096 17252 2102 17264
rect 2096 17224 2912 17252
rect 2096 17212 2102 17224
rect 2884 17193 2912 17224
rect 3970 17212 3976 17264
rect 4028 17252 4034 17264
rect 8754 17252 8760 17264
rect 4028 17224 8760 17252
rect 4028 17212 4034 17224
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 17313 17255 17371 17261
rect 15344 17224 15700 17252
rect 15344 17212 15350 17224
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 2038 17076 2044 17128
rect 2096 17076 2102 17128
rect 2240 17048 2268 17147
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17184 3295 17187
rect 7662 17187 7720 17193
rect 7662 17184 7674 17187
rect 3283 17156 7674 17184
rect 3283 17153 3295 17156
rect 3237 17147 3295 17153
rect 7662 17153 7674 17156
rect 7708 17153 7720 17187
rect 7662 17147 7720 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9214 17184 9220 17196
rect 9171 17156 9220 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9398 17193 9404 17196
rect 9392 17184 9404 17193
rect 9359 17156 9404 17184
rect 9392 17147 9404 17156
rect 9398 17144 9404 17147
rect 9456 17144 9462 17196
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11940 17156 12081 17184
rect 11940 17144 11946 17156
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12336 17187 12394 17193
rect 12336 17153 12348 17187
rect 12382 17184 12394 17187
rect 12382 17156 14964 17184
rect 12382 17153 12394 17156
rect 12336 17147 12394 17153
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17085 14887 17119
rect 14936 17116 14964 17156
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 15470 17184 15476 17196
rect 15243 17156 15476 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 15672 17193 15700 17224
rect 17313 17221 17325 17255
rect 17359 17252 17371 17255
rect 17494 17252 17500 17264
rect 17359 17224 17500 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 16390 17184 16396 17196
rect 15887 17156 16396 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 16632 17156 17141 17184
rect 16632 17144 16638 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17402 17144 17408 17196
rect 17460 17144 17466 17196
rect 16666 17116 16672 17128
rect 14936 17088 16672 17116
rect 14829 17079 14887 17085
rect 6549 17051 6607 17057
rect 6549 17048 6561 17051
rect 2240 17020 6561 17048
rect 6549 17017 6561 17020
rect 6595 17017 6607 17051
rect 14844 17048 14872 17079
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 15194 17048 15200 17060
rect 14844 17020 15200 17048
rect 6549 17011 6607 17017
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 12342 16980 12348 16992
rect 10551 16952 12348 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 13449 16983 13507 16989
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 15010 16980 15016 16992
rect 13495 16952 15016 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 16758 16940 16764 16992
rect 16816 16980 16822 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 16816 16952 17141 16980
rect 16816 16940 16822 16952
rect 17129 16949 17141 16952
rect 17175 16949 17187 16983
rect 17129 16943 17187 16949
rect 1104 16890 20884 16912
rect 1104 16838 3422 16890
rect 3474 16838 3486 16890
rect 3538 16838 3550 16890
rect 3602 16838 3614 16890
rect 3666 16838 3678 16890
rect 3730 16838 8367 16890
rect 8419 16838 8431 16890
rect 8483 16838 8495 16890
rect 8547 16838 8559 16890
rect 8611 16838 8623 16890
rect 8675 16838 13312 16890
rect 13364 16838 13376 16890
rect 13428 16838 13440 16890
rect 13492 16838 13504 16890
rect 13556 16838 13568 16890
rect 13620 16838 18257 16890
rect 18309 16838 18321 16890
rect 18373 16838 18385 16890
rect 18437 16838 18449 16890
rect 18501 16838 18513 16890
rect 18565 16838 20884 16890
rect 1104 16816 20884 16838
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3973 16779 4031 16785
rect 3973 16776 3985 16779
rect 3108 16748 3985 16776
rect 3108 16736 3114 16748
rect 3973 16745 3985 16748
rect 4019 16745 4031 16779
rect 3973 16739 4031 16745
rect 9398 16736 9404 16788
rect 9456 16776 9462 16788
rect 15841 16779 15899 16785
rect 15841 16776 15853 16779
rect 9456 16748 15853 16776
rect 9456 16736 9462 16748
rect 15841 16745 15853 16748
rect 15887 16745 15899 16779
rect 15841 16739 15899 16745
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 15194 16708 15200 16720
rect 14936 16680 15200 16708
rect 14936 16649 14964 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 15289 16711 15347 16717
rect 15289 16677 15301 16711
rect 15335 16708 15347 16711
rect 16574 16708 16580 16720
rect 15335 16680 16580 16708
rect 15335 16677 15347 16680
rect 15289 16671 15347 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 16758 16668 16764 16720
rect 16816 16668 16822 16720
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 14921 16643 14979 16649
rect 10919 16612 11008 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 1762 16532 1768 16584
rect 1820 16572 1826 16584
rect 2041 16575 2099 16581
rect 2041 16572 2053 16575
rect 1820 16544 2053 16572
rect 1820 16532 1826 16544
rect 2041 16541 2053 16544
rect 2087 16541 2099 16575
rect 2041 16535 2099 16541
rect 2130 16532 2136 16584
rect 2188 16532 2194 16584
rect 5258 16532 5264 16584
rect 5316 16572 5322 16584
rect 5353 16575 5411 16581
rect 5353 16572 5365 16575
rect 5316 16544 5365 16572
rect 5316 16532 5322 16544
rect 5353 16541 5365 16544
rect 5399 16541 5411 16575
rect 10980 16572 11008 16612
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15010 16600 15016 16652
rect 15068 16640 15074 16652
rect 15068 16612 15148 16640
rect 15068 16600 15074 16612
rect 11882 16572 11888 16584
rect 10980 16544 11888 16572
rect 5353 16535 5411 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 15120 16581 15148 16612
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15620 16612 15761 16640
rect 15620 16600 15626 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16298 16640 16304 16652
rect 15979 16612 16304 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 15105 16575 15163 16581
rect 15105 16541 15117 16575
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 1854 16464 1860 16516
rect 1912 16504 1918 16516
rect 2222 16504 2228 16516
rect 1912 16476 2228 16504
rect 1912 16464 1918 16476
rect 2222 16464 2228 16476
rect 2280 16464 2286 16516
rect 2314 16464 2320 16516
rect 2372 16504 2378 16516
rect 5086 16507 5144 16513
rect 5086 16504 5098 16507
rect 2372 16476 5098 16504
rect 2372 16464 2378 16476
rect 5086 16473 5098 16476
rect 5132 16473 5144 16507
rect 5086 16467 5144 16473
rect 11140 16507 11198 16513
rect 11140 16473 11152 16507
rect 11186 16504 11198 16507
rect 13170 16504 13176 16516
rect 11186 16476 13176 16504
rect 11186 16473 11198 16476
rect 11140 16467 11198 16473
rect 13170 16464 13176 16476
rect 13228 16464 13234 16516
rect 1946 16396 1952 16448
rect 2004 16445 2010 16448
rect 2004 16399 2013 16445
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 12710 16436 12716 16448
rect 12299 16408 12716 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 2004 16396 2010 16399
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 15764 16436 15792 16603
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17494 16600 17500 16652
rect 17552 16640 17558 16652
rect 17552 16612 18920 16640
rect 17552 16600 17558 16612
rect 18892 16584 18920 16612
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19300 16612 19472 16640
rect 19300 16600 19306 16612
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16572 16083 16575
rect 16114 16572 16120 16584
rect 16071 16544 16120 16572
rect 16071 16541 16083 16544
rect 16025 16535 16083 16541
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 16850 16532 16856 16584
rect 16908 16532 16914 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17052 16544 17417 16572
rect 16577 16507 16635 16513
rect 16577 16473 16589 16507
rect 16623 16504 16635 16507
rect 16666 16504 16672 16516
rect 16623 16476 16672 16504
rect 16623 16473 16635 16476
rect 16577 16467 16635 16473
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 17052 16436 17080 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 17770 16464 17776 16516
rect 17828 16464 17834 16516
rect 15764 16408 17080 16436
rect 18708 16436 18736 16535
rect 18874 16532 18880 16584
rect 18932 16532 18938 16584
rect 19444 16581 19472 16612
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 18785 16507 18843 16513
rect 18785 16473 18797 16507
rect 18831 16504 18843 16507
rect 19628 16504 19656 16535
rect 19702 16532 19708 16584
rect 19760 16532 19766 16584
rect 19794 16532 19800 16584
rect 19852 16532 19858 16584
rect 18831 16476 19656 16504
rect 18831 16473 18843 16476
rect 18785 16467 18843 16473
rect 19702 16436 19708 16448
rect 18708 16408 19708 16436
rect 19702 16396 19708 16408
rect 19760 16396 19766 16448
rect 20070 16396 20076 16448
rect 20128 16396 20134 16448
rect 1104 16346 21043 16368
rect 1104 16294 5894 16346
rect 5946 16294 5958 16346
rect 6010 16294 6022 16346
rect 6074 16294 6086 16346
rect 6138 16294 6150 16346
rect 6202 16294 10839 16346
rect 10891 16294 10903 16346
rect 10955 16294 10967 16346
rect 11019 16294 11031 16346
rect 11083 16294 11095 16346
rect 11147 16294 15784 16346
rect 15836 16294 15848 16346
rect 15900 16294 15912 16346
rect 15964 16294 15976 16346
rect 16028 16294 16040 16346
rect 16092 16294 20729 16346
rect 20781 16294 20793 16346
rect 20845 16294 20857 16346
rect 20909 16294 20921 16346
rect 20973 16294 20985 16346
rect 21037 16294 21043 16346
rect 1104 16272 21043 16294
rect 2314 16192 2320 16244
rect 2372 16192 2378 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16390 16232 16396 16244
rect 16163 16204 16396 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 16632 16204 17233 16232
rect 16632 16192 16638 16204
rect 17221 16201 17233 16204
rect 17267 16232 17279 16235
rect 17310 16232 17316 16244
rect 17267 16204 17316 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 19613 16235 19671 16241
rect 19613 16201 19625 16235
rect 19659 16232 19671 16235
rect 19794 16232 19800 16244
rect 19659 16204 19800 16232
rect 19659 16201 19671 16204
rect 19613 16195 19671 16201
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 2038 16124 2044 16176
rect 2096 16164 2102 16176
rect 2222 16164 2228 16176
rect 2096 16136 2228 16164
rect 2096 16124 2102 16136
rect 2222 16124 2228 16136
rect 2280 16124 2286 16176
rect 4982 16124 4988 16176
rect 5040 16173 5046 16176
rect 5040 16164 5052 16173
rect 9484 16167 9542 16173
rect 5040 16136 5085 16164
rect 5040 16127 5052 16136
rect 9484 16133 9496 16167
rect 9530 16164 9542 16167
rect 9582 16164 9588 16176
rect 9530 16136 9588 16164
rect 9530 16133 9542 16136
rect 9484 16127 9542 16133
rect 5040 16124 5046 16127
rect 9582 16124 9588 16136
rect 9640 16124 9646 16176
rect 12342 16124 12348 16176
rect 12400 16164 12406 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 12400 16136 17141 16164
rect 12400 16124 12406 16136
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 2004 16068 2145 16096
rect 2004 16056 2010 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2498 16056 2504 16108
rect 2556 16096 2562 16108
rect 7662 16099 7720 16105
rect 7662 16096 7674 16099
rect 2556 16068 7674 16096
rect 2556 16056 2562 16068
rect 7662 16065 7674 16068
rect 7708 16065 7720 16099
rect 7662 16059 7720 16065
rect 7926 16056 7932 16108
rect 7984 16056 7990 16108
rect 9214 16056 9220 16108
rect 9272 16056 9278 16108
rect 12244 16099 12302 16105
rect 12244 16065 12256 16099
rect 12290 16096 12302 16099
rect 13722 16096 13728 16108
rect 12290 16068 13728 16096
rect 12290 16065 12302 16068
rect 12244 16059 12302 16065
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 14550 16056 14556 16108
rect 14608 16056 14614 16108
rect 14844 16105 14872 16136
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15654 16096 15660 16108
rect 15059 16068 15660 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 16040 16105 16068 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16850 16096 16856 16108
rect 16347 16068 16856 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 17402 16096 17408 16108
rect 17359 16068 17408 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 18874 16056 18880 16108
rect 18932 16096 18938 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 18932 16068 19441 16096
rect 18932 16056 18938 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 1857 16031 1915 16037
rect 1857 16028 1869 16031
rect 1820 16000 1869 16028
rect 1820 15988 1826 16000
rect 1857 15997 1869 16000
rect 1903 16028 1915 16031
rect 2038 16028 2044 16040
rect 1903 16000 2044 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 5258 15988 5264 16040
rect 5316 15988 5322 16040
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11940 16000 11989 16028
rect 11940 15988 11946 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 11977 15991 12035 15997
rect 14752 16000 16957 16028
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2130 15960 2136 15972
rect 1995 15932 2136 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2130 15920 2136 15932
rect 2188 15960 2194 15972
rect 14752 15969 14780 16000
rect 16945 15997 16957 16000
rect 16991 16028 17003 16031
rect 17494 16028 17500 16040
rect 16991 16000 17500 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 19245 16031 19303 16037
rect 19245 15997 19257 16031
rect 19291 16028 19303 16031
rect 19886 16028 19892 16040
rect 19291 16000 19892 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 14737 15963 14795 15969
rect 14737 15960 14749 15963
rect 2188 15932 4016 15960
rect 2188 15920 2194 15932
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 2372 15864 3893 15892
rect 2372 15852 2378 15864
rect 3881 15861 3893 15864
rect 3927 15861 3939 15895
rect 3988 15892 4016 15932
rect 13280 15932 14749 15960
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 3988 15864 6561 15892
rect 3881 15855 3939 15861
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 6730 15852 6736 15904
rect 6788 15892 6794 15904
rect 7926 15892 7932 15904
rect 6788 15864 7932 15892
rect 6788 15852 6794 15864
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 10597 15895 10655 15901
rect 10597 15861 10609 15895
rect 10643 15892 10655 15895
rect 13280 15892 13308 15932
rect 14737 15929 14749 15932
rect 14783 15929 14795 15963
rect 14737 15923 14795 15929
rect 14826 15920 14832 15972
rect 14884 15960 14890 15972
rect 14921 15963 14979 15969
rect 14921 15960 14933 15963
rect 14884 15932 14933 15960
rect 14884 15920 14890 15932
rect 14921 15929 14933 15932
rect 14967 15929 14979 15963
rect 14921 15923 14979 15929
rect 16298 15920 16304 15972
rect 16356 15920 16362 15972
rect 16390 15920 16396 15972
rect 16448 15960 16454 15972
rect 19260 15960 19288 15991
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 16448 15932 19288 15960
rect 16448 15920 16454 15932
rect 10643 15864 13308 15892
rect 13357 15895 13415 15901
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 13357 15861 13369 15895
rect 13403 15892 13415 15895
rect 14458 15892 14464 15904
rect 13403 15864 14464 15892
rect 13403 15861 13415 15864
rect 13357 15855 13415 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15289 15895 15347 15901
rect 15289 15861 15301 15895
rect 15335 15892 15347 15895
rect 15378 15892 15384 15904
rect 15335 15864 15384 15892
rect 15335 15861 15347 15864
rect 15289 15855 15347 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 1104 15802 20884 15824
rect 1104 15750 3422 15802
rect 3474 15750 3486 15802
rect 3538 15750 3550 15802
rect 3602 15750 3614 15802
rect 3666 15750 3678 15802
rect 3730 15750 8367 15802
rect 8419 15750 8431 15802
rect 8483 15750 8495 15802
rect 8547 15750 8559 15802
rect 8611 15750 8623 15802
rect 8675 15750 13312 15802
rect 13364 15750 13376 15802
rect 13428 15750 13440 15802
rect 13492 15750 13504 15802
rect 13556 15750 13568 15802
rect 13620 15750 18257 15802
rect 18309 15750 18321 15802
rect 18373 15750 18385 15802
rect 18437 15750 18449 15802
rect 18501 15750 18513 15802
rect 18565 15750 20884 15802
rect 1104 15728 20884 15750
rect 2498 15648 2504 15700
rect 2556 15648 2562 15700
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 5316 15660 5733 15688
rect 5316 15648 5322 15660
rect 5721 15657 5733 15660
rect 5767 15688 5779 15691
rect 6730 15688 6736 15700
rect 5767 15660 6736 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 16908 15660 17141 15688
rect 16908 15648 16914 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 17310 15648 17316 15700
rect 17368 15648 17374 15700
rect 19702 15648 19708 15700
rect 19760 15688 19766 15700
rect 19981 15691 20039 15697
rect 19981 15688 19993 15691
rect 19760 15660 19993 15688
rect 19760 15648 19766 15660
rect 19981 15657 19993 15660
rect 20027 15657 20039 15691
rect 19981 15651 20039 15657
rect 16666 15580 16672 15632
rect 16724 15620 16730 15632
rect 17770 15620 17776 15632
rect 16724 15592 17776 15620
rect 16724 15580 16730 15592
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 17310 15552 17316 15564
rect 14516 15524 17316 15552
rect 14516 15512 14522 15524
rect 17310 15512 17316 15524
rect 17368 15552 17374 15564
rect 19334 15552 19340 15564
rect 17368 15524 19340 15552
rect 17368 15512 17374 15524
rect 19334 15512 19340 15524
rect 19392 15552 19398 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19392 15524 19441 15552
rect 19392 15512 19398 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 2130 15444 2136 15496
rect 2188 15444 2194 15496
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 5810 15484 5816 15496
rect 2363 15456 5816 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 17402 15444 17408 15496
rect 17460 15484 17466 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 17460 15456 18153 15484
rect 17460 15444 17466 15456
rect 18141 15453 18153 15456
rect 18187 15484 18199 15487
rect 19720 15484 19748 15648
rect 18187 15456 19748 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 7006 15376 7012 15428
rect 7064 15416 7070 15428
rect 9950 15416 9956 15428
rect 7064 15388 9956 15416
rect 7064 15376 7070 15388
rect 9950 15376 9956 15388
rect 10008 15416 10014 15428
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 10008 15388 10425 15416
rect 10008 15376 10014 15388
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10413 15379 10471 15385
rect 17297 15419 17355 15425
rect 17297 15385 17309 15419
rect 17343 15416 17355 15419
rect 17420 15416 17448 15444
rect 17343 15388 17448 15416
rect 17343 15385 17355 15388
rect 17297 15379 17355 15385
rect 17494 15376 17500 15428
rect 17552 15376 17558 15428
rect 19518 15376 19524 15428
rect 19576 15416 19582 15428
rect 19797 15419 19855 15425
rect 19797 15416 19809 15419
rect 19576 15388 19809 15416
rect 19576 15376 19582 15388
rect 19797 15385 19809 15388
rect 19843 15385 19855 15419
rect 19797 15379 19855 15385
rect 11882 15308 11888 15360
rect 11940 15308 11946 15360
rect 18046 15308 18052 15360
rect 18104 15308 18110 15360
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 18196 15320 19625 15348
rect 18196 15308 18202 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 19702 15308 19708 15360
rect 19760 15308 19766 15360
rect 1104 15258 21043 15280
rect 1104 15206 5894 15258
rect 5946 15206 5958 15258
rect 6010 15206 6022 15258
rect 6074 15206 6086 15258
rect 6138 15206 6150 15258
rect 6202 15206 10839 15258
rect 10891 15206 10903 15258
rect 10955 15206 10967 15258
rect 11019 15206 11031 15258
rect 11083 15206 11095 15258
rect 11147 15206 15784 15258
rect 15836 15206 15848 15258
rect 15900 15206 15912 15258
rect 15964 15206 15976 15258
rect 16028 15206 16040 15258
rect 16092 15206 20729 15258
rect 20781 15206 20793 15258
rect 20845 15206 20857 15258
rect 20909 15206 20921 15258
rect 20973 15206 20985 15258
rect 21037 15206 21043 15258
rect 1104 15184 21043 15206
rect 9950 15104 9956 15156
rect 10008 15104 10014 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 14550 15144 14556 15156
rect 13311 15116 14556 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15654 15104 15660 15156
rect 15712 15144 15718 15156
rect 19137 15147 19195 15153
rect 15712 15116 18000 15144
rect 15712 15104 15718 15116
rect 7000 15079 7058 15085
rect 7000 15045 7012 15079
rect 7046 15076 7058 15079
rect 7098 15076 7104 15088
rect 7046 15048 7104 15076
rect 7046 15045 7058 15048
rect 7000 15039 7058 15045
rect 7098 15036 7104 15048
rect 7156 15036 7162 15088
rect 8665 15079 8723 15085
rect 8665 15045 8677 15079
rect 8711 15076 8723 15079
rect 8754 15076 8760 15088
rect 8711 15048 8760 15076
rect 8711 15045 8723 15048
rect 8665 15039 8723 15045
rect 8754 15036 8760 15048
rect 8812 15036 8818 15088
rect 14568 15076 14596 15104
rect 17972 15088 18000 15116
rect 19137 15113 19149 15147
rect 19183 15144 19195 15147
rect 19518 15144 19524 15156
rect 19183 15116 19524 15144
rect 19183 15113 19195 15116
rect 19137 15107 19195 15113
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 14568 15048 15976 15076
rect 2222 14968 2228 15020
rect 2280 14968 2286 15020
rect 12152 15011 12210 15017
rect 12152 14977 12164 15011
rect 12198 15008 12210 15011
rect 14921 15011 14979 15017
rect 12198 14980 14872 15008
rect 12198 14977 12210 14980
rect 12152 14971 12210 14977
rect 1946 14900 1952 14952
rect 2004 14900 2010 14952
rect 6730 14900 6736 14952
rect 6788 14900 6794 14952
rect 11882 14900 11888 14952
rect 11940 14900 11946 14952
rect 14844 14940 14872 14980
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15010 15008 15016 15020
rect 14967 14980 15016 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15948 15017 15976 15048
rect 17954 15036 17960 15088
rect 18012 15036 18018 15088
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 15933 15011 15991 15017
rect 15252 14980 15792 15008
rect 15252 14968 15258 14980
rect 15654 14940 15660 14952
rect 14844 14912 15660 14940
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 15764 14949 15792 14980
rect 15933 14977 15945 15011
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 17678 14968 17684 15020
rect 17736 14968 17742 15020
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19576 14980 19993 15008
rect 19576 14968 19582 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 16390 14940 16396 14952
rect 15795 14912 16396 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 19702 14940 19708 14952
rect 19168 14912 19708 14940
rect 14918 14832 14924 14884
rect 14976 14872 14982 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 14976 14844 15025 14872
rect 14976 14832 14982 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14841 15163 14875
rect 15105 14835 15163 14841
rect 16117 14875 16175 14881
rect 16117 14841 16129 14875
rect 16163 14872 16175 14875
rect 18138 14872 18144 14884
rect 16163 14844 18144 14872
rect 16163 14841 16175 14844
rect 16117 14835 16175 14841
rect 2038 14764 2044 14816
rect 2096 14764 2102 14816
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 6914 14804 6920 14816
rect 2455 14776 6920 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 13998 14804 14004 14816
rect 8159 14776 14004 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14734 14764 14740 14816
rect 14792 14764 14798 14816
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 15120 14804 15148 14835
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 19168 14816 19196 14912
rect 19702 14900 19708 14912
rect 19760 14940 19766 14952
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 19760 14912 20177 14940
rect 19760 14900 19766 14912
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 14884 14776 15148 14804
rect 14884 14764 14890 14776
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 18969 14807 19027 14813
rect 18969 14804 18981 14807
rect 17184 14776 18981 14804
rect 17184 14764 17190 14776
rect 18969 14773 18981 14776
rect 19015 14773 19027 14807
rect 18969 14767 19027 14773
rect 19150 14764 19156 14816
rect 19208 14764 19214 14816
rect 19794 14764 19800 14816
rect 19852 14764 19858 14816
rect 1104 14714 20884 14736
rect 1104 14662 3422 14714
rect 3474 14662 3486 14714
rect 3538 14662 3550 14714
rect 3602 14662 3614 14714
rect 3666 14662 3678 14714
rect 3730 14662 8367 14714
rect 8419 14662 8431 14714
rect 8483 14662 8495 14714
rect 8547 14662 8559 14714
rect 8611 14662 8623 14714
rect 8675 14662 13312 14714
rect 13364 14662 13376 14714
rect 13428 14662 13440 14714
rect 13492 14662 13504 14714
rect 13556 14662 13568 14714
rect 13620 14662 18257 14714
rect 18309 14662 18321 14714
rect 18373 14662 18385 14714
rect 18437 14662 18449 14714
rect 18501 14662 18513 14714
rect 18565 14662 20884 14714
rect 1104 14640 20884 14662
rect 1857 14603 1915 14609
rect 1857 14569 1869 14603
rect 1903 14600 1915 14603
rect 2222 14600 2228 14612
rect 1903 14572 2228 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5868 14572 6009 14600
rect 5868 14560 5874 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 14921 14603 14979 14609
rect 14921 14600 14933 14603
rect 14884 14572 14933 14600
rect 14884 14560 14890 14572
rect 14921 14569 14933 14572
rect 14967 14569 14979 14603
rect 14921 14563 14979 14569
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 15712 14572 16773 14600
rect 15712 14560 15718 14572
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 18046 14600 18052 14612
rect 16761 14563 16819 14569
rect 17328 14572 18052 14600
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 15105 14535 15163 14541
rect 15105 14532 15117 14535
rect 13136 14504 15117 14532
rect 13136 14492 13142 14504
rect 15105 14501 15117 14504
rect 15151 14532 15163 14535
rect 15151 14504 15700 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15672 14476 15700 14504
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 10744 14436 12434 14464
rect 10744 14424 10750 14436
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 2096 14368 2145 14396
rect 2096 14356 2102 14368
rect 2133 14365 2145 14368
rect 2179 14396 2191 14399
rect 5353 14399 5411 14405
rect 2179 14368 4016 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 1854 14288 1860 14340
rect 1912 14288 1918 14340
rect 2038 14220 2044 14272
rect 2096 14220 2102 14272
rect 3988 14269 4016 14368
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5534 14396 5540 14408
rect 5399 14368 5540 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 6788 14368 7389 14396
rect 6788 14356 6794 14368
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 7377 14359 7435 14365
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 11882 14396 11888 14408
rect 9723 14368 11888 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12406 14396 12434 14436
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 15381 14467 15439 14473
rect 15381 14464 15393 14467
rect 14424 14436 15393 14464
rect 14424 14424 14430 14436
rect 15381 14433 15393 14436
rect 15427 14464 15439 14467
rect 15470 14464 15476 14476
rect 15427 14436 15476 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 16942 14396 16948 14408
rect 12406 14368 16948 14396
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 5086 14331 5144 14337
rect 5086 14328 5098 14331
rect 4212 14300 5098 14328
rect 4212 14288 4218 14300
rect 5086 14297 5098 14300
rect 5132 14297 5144 14331
rect 5086 14291 5144 14297
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 7110 14331 7168 14337
rect 7110 14328 7122 14331
rect 6972 14300 7122 14328
rect 6972 14288 6978 14300
rect 7110 14297 7122 14300
rect 7156 14297 7168 14331
rect 7110 14291 7168 14297
rect 9944 14331 10002 14337
rect 9944 14297 9956 14331
rect 9990 14328 10002 14331
rect 12250 14328 12256 14340
rect 9990 14300 12256 14328
rect 9990 14297 10002 14300
rect 9944 14291 10002 14297
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 17052 14328 17080 14359
rect 17126 14356 17132 14408
rect 17184 14356 17190 14408
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 17328 14396 17356 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 19628 14532 19656 14560
rect 17420 14504 19656 14532
rect 17420 14408 17448 14504
rect 19794 14464 19800 14476
rect 18064 14436 19800 14464
rect 17267 14368 17356 14396
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 17402 14356 17408 14408
rect 17460 14356 17466 14408
rect 18064 14405 18092 14436
rect 19794 14424 19800 14436
rect 19852 14464 19858 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19852 14436 19993 14464
rect 19852 14424 19858 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 19334 14396 19340 14408
rect 18371 14368 19340 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 18138 14328 18144 14340
rect 17052 14300 18144 14328
rect 18138 14288 18144 14300
rect 18196 14288 18202 14340
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 14550 14260 14556 14272
rect 11103 14232 14556 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17865 14263 17923 14269
rect 17865 14260 17877 14263
rect 17184 14232 17877 14260
rect 17184 14220 17190 14232
rect 17865 14229 17877 14232
rect 17911 14229 17923 14263
rect 17865 14223 17923 14229
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18233 14263 18291 14269
rect 18233 14260 18245 14263
rect 18012 14232 18245 14260
rect 18012 14220 18018 14232
rect 18233 14229 18245 14232
rect 18279 14260 18291 14263
rect 19334 14260 19340 14272
rect 18279 14232 19340 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19426 14220 19432 14272
rect 19484 14220 19490 14272
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 19702 14260 19708 14272
rect 19659 14232 19708 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 1104 14170 21043 14192
rect 1104 14118 5894 14170
rect 5946 14118 5958 14170
rect 6010 14118 6022 14170
rect 6074 14118 6086 14170
rect 6138 14118 6150 14170
rect 6202 14118 10839 14170
rect 10891 14118 10903 14170
rect 10955 14118 10967 14170
rect 11019 14118 11031 14170
rect 11083 14118 11095 14170
rect 11147 14118 15784 14170
rect 15836 14118 15848 14170
rect 15900 14118 15912 14170
rect 15964 14118 15976 14170
rect 16028 14118 16040 14170
rect 16092 14118 20729 14170
rect 20781 14118 20793 14170
rect 20845 14118 20857 14170
rect 20909 14118 20921 14170
rect 20973 14118 20985 14170
rect 21037 14118 21043 14170
rect 1104 14096 21043 14118
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 10686 14056 10692 14068
rect 9079 14028 10692 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 13078 14056 13084 14068
rect 11103 14028 13084 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 14826 14056 14832 14068
rect 13219 14028 14832 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 19426 14056 19432 14068
rect 15948 14028 19432 14056
rect 15948 13988 15976 14028
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19518 14016 19524 14068
rect 19576 14016 19582 14068
rect 19702 14016 19708 14068
rect 19760 14016 19766 14068
rect 11992 13960 12434 13988
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 5718 13920 5724 13932
rect 2547 13892 5724 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2130 13812 2136 13864
rect 2188 13812 2194 13864
rect 2332 13852 2360 13883
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 7920 13923 7978 13929
rect 7920 13889 7932 13923
rect 7966 13920 7978 13923
rect 11992 13920 12020 13960
rect 12066 13929 12072 13932
rect 7966 13892 12020 13920
rect 7966 13889 7978 13892
rect 7920 13883 7978 13889
rect 12060 13883 12072 13929
rect 12066 13880 12072 13883
rect 12124 13880 12130 13932
rect 12406 13920 12434 13960
rect 13188 13960 15976 13988
rect 17129 13991 17187 13997
rect 12406 13892 12848 13920
rect 3970 13852 3976 13864
rect 2332 13824 3976 13852
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 4120 13824 5365 13852
rect 4120 13812 4126 13824
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5500 13824 5641 13852
rect 5500 13812 5506 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 7653 13855 7711 13861
rect 7653 13852 7665 13855
rect 5675 13824 7665 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 7653 13821 7665 13824
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 2148 13784 2176 13812
rect 2682 13784 2688 13796
rect 2148 13756 2688 13784
rect 2682 13744 2688 13756
rect 2740 13744 2746 13796
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 4065 13719 4123 13725
rect 4065 13716 4077 13719
rect 3292 13688 4077 13716
rect 3292 13676 3298 13688
rect 4065 13685 4077 13688
rect 4111 13685 4123 13719
rect 7668 13716 7696 13815
rect 9306 13812 9312 13864
rect 9364 13852 9370 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9364 13824 9505 13852
rect 9364 13812 9370 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10410 13852 10416 13864
rect 9815 13824 10416 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 12820 13852 12848 13892
rect 13188 13852 13216 13960
rect 17129 13957 17141 13991
rect 17175 13988 17187 13991
rect 17402 13988 17408 14000
rect 17175 13960 17408 13988
rect 17175 13957 17187 13960
rect 17129 13951 17187 13957
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 18693 13991 18751 13997
rect 18693 13957 18705 13991
rect 18739 13988 18751 13991
rect 19536 13988 19564 14016
rect 18739 13960 19564 13988
rect 18739 13957 18751 13960
rect 18693 13951 18751 13957
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17000 13892 17080 13920
rect 17000 13880 17006 13892
rect 12820 13824 13216 13852
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 17052 13852 17080 13892
rect 17218 13880 17224 13932
rect 17276 13920 17282 13932
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 17276 13892 17509 13920
rect 17276 13880 17282 13892
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 17497 13883 17555 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 18598 13920 18604 13932
rect 18555 13892 18604 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 13780 13824 16988 13852
rect 17052 13824 18337 13852
rect 13780 13812 13786 13824
rect 16960 13793 16988 13824
rect 18325 13821 18337 13824
rect 18371 13852 18383 13855
rect 18616 13852 18644 13880
rect 19352 13852 19380 13883
rect 19426 13880 19432 13932
rect 19484 13880 19490 13932
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19536 13852 19564 13883
rect 18371 13824 18552 13852
rect 18616 13824 19380 13852
rect 19444 13824 19564 13852
rect 18371 13821 18383 13824
rect 18325 13815 18383 13821
rect 16945 13787 17003 13793
rect 16945 13753 16957 13787
rect 16991 13753 17003 13787
rect 18524 13784 18552 13824
rect 19444 13784 19472 13824
rect 18524 13756 19472 13784
rect 16945 13747 17003 13753
rect 19518 13744 19524 13796
rect 19576 13784 19582 13796
rect 19886 13784 19892 13796
rect 19576 13756 19892 13784
rect 19576 13744 19582 13756
rect 19886 13744 19892 13756
rect 19944 13744 19950 13796
rect 7926 13716 7932 13728
rect 7668 13688 7932 13716
rect 4065 13679 4123 13685
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 17126 13676 17132 13728
rect 17184 13676 17190 13728
rect 1104 13626 20884 13648
rect 1104 13574 3422 13626
rect 3474 13574 3486 13626
rect 3538 13574 3550 13626
rect 3602 13574 3614 13626
rect 3666 13574 3678 13626
rect 3730 13574 8367 13626
rect 8419 13574 8431 13626
rect 8483 13574 8495 13626
rect 8547 13574 8559 13626
rect 8611 13574 8623 13626
rect 8675 13574 13312 13626
rect 13364 13574 13376 13626
rect 13428 13574 13440 13626
rect 13492 13574 13504 13626
rect 13556 13574 13568 13626
rect 13620 13574 18257 13626
rect 18309 13574 18321 13626
rect 18373 13574 18385 13626
rect 18437 13574 18449 13626
rect 18501 13574 18513 13626
rect 18565 13574 20884 13626
rect 1104 13552 20884 13574
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 15013 13515 15071 13521
rect 15013 13481 15025 13515
rect 15059 13512 15071 13515
rect 15286 13512 15292 13524
rect 15059 13484 15292 13512
rect 15059 13481 15071 13484
rect 15013 13475 15071 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 4154 13444 4160 13456
rect 2363 13416 4160 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 4154 13404 4160 13416
rect 4212 13404 4218 13456
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 2038 13376 2044 13388
rect 1903 13348 2044 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 2038 13336 2044 13348
rect 2096 13376 2102 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2096 13348 2789 13376
rect 2096 13336 2102 13348
rect 2777 13345 2789 13348
rect 2823 13376 2835 13379
rect 3234 13376 3240 13388
rect 2823 13348 3240 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 7926 13336 7932 13388
rect 7984 13336 7990 13388
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17000 13348 17540 13376
rect 17000 13336 17006 13348
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 1964 13172 1992 13271
rect 2130 13268 2136 13320
rect 2188 13268 2194 13320
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2740 13280 2973 13308
rect 2740 13268 2746 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 7662 13311 7720 13317
rect 7662 13308 7674 13311
rect 5776 13280 7674 13308
rect 5776 13268 5782 13280
rect 7662 13277 7674 13280
rect 7708 13277 7720 13311
rect 7662 13271 7720 13277
rect 11790 13268 11796 13320
rect 11848 13268 11854 13320
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 14829 13311 14887 13317
rect 14829 13308 14841 13311
rect 14700 13280 14841 13308
rect 14700 13268 14706 13280
rect 14829 13277 14841 13280
rect 14875 13277 14887 13311
rect 14829 13271 14887 13277
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17129 13311 17187 13317
rect 17129 13308 17141 13311
rect 17092 13280 17141 13308
rect 17092 13268 17098 13280
rect 17129 13277 17141 13280
rect 17175 13308 17187 13311
rect 17218 13308 17224 13320
rect 17175 13280 17224 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17402 13268 17408 13320
rect 17460 13268 17466 13320
rect 17512 13308 17540 13348
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17512 13280 17601 13308
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19392 13280 19625 13308
rect 19392 13268 19398 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 3145 13243 3203 13249
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 5086 13243 5144 13249
rect 5086 13240 5098 13243
rect 3191 13212 5098 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 5086 13209 5098 13212
rect 5132 13209 5144 13243
rect 5086 13203 5144 13209
rect 12060 13243 12118 13249
rect 12060 13209 12072 13243
rect 12106 13240 12118 13243
rect 19426 13240 19432 13252
rect 12106 13212 19432 13240
rect 12106 13209 12118 13212
rect 12060 13203 12118 13209
rect 19426 13200 19432 13212
rect 19484 13200 19490 13252
rect 2222 13172 2228 13184
rect 1964 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13172 2286 13184
rect 6549 13175 6607 13181
rect 6549 13172 6561 13175
rect 2280 13144 6561 13172
rect 2280 13132 2286 13144
rect 6549 13141 6561 13144
rect 6595 13141 6607 13175
rect 6549 13135 6607 13141
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 15010 13172 15016 13184
rect 13219 13144 15016 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15562 13132 15568 13184
rect 15620 13132 15626 13184
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13172 17003 13175
rect 17126 13172 17132 13184
rect 16991 13144 17132 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19705 13175 19763 13181
rect 19705 13172 19717 13175
rect 19576 13144 19717 13172
rect 19576 13132 19582 13144
rect 19705 13141 19717 13144
rect 19751 13141 19763 13175
rect 19705 13135 19763 13141
rect 1104 13082 21043 13104
rect 1104 13030 5894 13082
rect 5946 13030 5958 13082
rect 6010 13030 6022 13082
rect 6074 13030 6086 13082
rect 6138 13030 6150 13082
rect 6202 13030 10839 13082
rect 10891 13030 10903 13082
rect 10955 13030 10967 13082
rect 11019 13030 11031 13082
rect 11083 13030 11095 13082
rect 11147 13030 15784 13082
rect 15836 13030 15848 13082
rect 15900 13030 15912 13082
rect 15964 13030 15976 13082
rect 16028 13030 16040 13082
rect 16092 13030 20729 13082
rect 20781 13030 20793 13082
rect 20845 13030 20857 13082
rect 20909 13030 20921 13082
rect 20973 13030 20985 13082
rect 21037 13030 21043 13082
rect 1104 13008 21043 13030
rect 1955 12971 2013 12977
rect 1955 12937 1967 12971
rect 2001 12968 2013 12971
rect 2130 12968 2136 12980
rect 2001 12940 2136 12968
rect 2001 12937 2013 12940
rect 1955 12931 2013 12937
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15344 12940 17632 12968
rect 15344 12928 15350 12940
rect 1854 12860 1860 12912
rect 1912 12860 1918 12912
rect 2038 12860 2044 12912
rect 2096 12860 2102 12912
rect 6816 12903 6874 12909
rect 6816 12869 6828 12903
rect 6862 12900 6874 12903
rect 6914 12900 6920 12912
rect 6862 12872 6920 12900
rect 6862 12869 6874 12872
rect 6816 12863 6874 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 12060 12903 12118 12909
rect 12060 12869 12072 12903
rect 12106 12900 12118 12903
rect 16758 12900 16764 12912
rect 12106 12872 16764 12900
rect 12106 12869 12118 12872
rect 12060 12863 12118 12869
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 17402 12900 17408 12912
rect 17144 12872 17408 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2222 12832 2228 12844
rect 2179 12804 2228 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14700 12804 14749 12832
rect 14700 12792 14706 12804
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17144 12841 17172 12872
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 17604 12900 17632 12940
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 17865 12971 17923 12977
rect 17865 12968 17877 12971
rect 17736 12940 17877 12968
rect 17736 12928 17742 12940
rect 17865 12937 17877 12940
rect 17911 12937 17923 12971
rect 17865 12931 17923 12937
rect 18598 12900 18604 12912
rect 17604 12872 18604 12900
rect 18598 12860 18604 12872
rect 18656 12900 18662 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18656 12872 19257 12900
rect 18656 12860 18662 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 19245 12863 19303 12869
rect 19429 12903 19487 12909
rect 19429 12869 19441 12903
rect 19475 12900 19487 12903
rect 19889 12903 19947 12909
rect 19889 12900 19901 12903
rect 19475 12872 19901 12900
rect 19475 12869 19487 12872
rect 19429 12863 19487 12869
rect 19889 12869 19901 12872
rect 19935 12869 19947 12903
rect 19889 12863 19947 12869
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 17000 12804 17049 12832
rect 17000 12792 17006 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 14826 12724 14832 12776
rect 14884 12724 14890 12776
rect 15102 12724 15108 12776
rect 15160 12724 15166 12776
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 17144 12764 17172 12795
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17954 12832 17960 12844
rect 17276 12804 17960 12832
rect 17276 12792 17282 12804
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 19260 12832 19288 12863
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19260 12804 20177 12832
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 16172 12736 17172 12764
rect 16172 12724 16178 12736
rect 7929 12631 7987 12637
rect 7929 12597 7941 12631
rect 7975 12628 7987 12631
rect 8018 12628 8024 12640
rect 7975 12600 8024 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 13173 12631 13231 12637
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 14090 12628 14096 12640
rect 13219 12600 14096 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 14090 12588 14096 12600
rect 14148 12628 14154 12640
rect 15102 12628 15108 12640
rect 14148 12600 15108 12628
rect 14148 12588 14154 12600
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 16942 12628 16948 12640
rect 16899 12600 16948 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 19168 12628 19196 12792
rect 19610 12724 19616 12776
rect 19668 12764 19674 12776
rect 19889 12767 19947 12773
rect 19889 12764 19901 12767
rect 19668 12736 19901 12764
rect 19668 12724 19674 12736
rect 19889 12733 19901 12736
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 19426 12656 19432 12708
rect 19484 12656 19490 12708
rect 19978 12628 19984 12640
rect 19168 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12628 20042 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 20036 12600 20085 12628
rect 20036 12588 20042 12600
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 20073 12591 20131 12597
rect 1104 12538 20884 12560
rect 1104 12486 3422 12538
rect 3474 12486 3486 12538
rect 3538 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 8367 12538
rect 8419 12486 8431 12538
rect 8483 12486 8495 12538
rect 8547 12486 8559 12538
rect 8611 12486 8623 12538
rect 8675 12486 13312 12538
rect 13364 12486 13376 12538
rect 13428 12486 13440 12538
rect 13492 12486 13504 12538
rect 13556 12486 13568 12538
rect 13620 12486 18257 12538
rect 18309 12486 18321 12538
rect 18373 12486 18385 12538
rect 18437 12486 18449 12538
rect 18501 12486 18513 12538
rect 18565 12486 20884 12538
rect 1104 12464 20884 12486
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 14642 12424 14648 12436
rect 11195 12396 14648 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15252 12396 15301 12424
rect 15252 12384 15258 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 19610 12384 19616 12436
rect 19668 12384 19674 12436
rect 2222 12356 2228 12368
rect 1964 12328 2228 12356
rect 1964 12229 1992 12328
rect 2222 12316 2228 12328
rect 2280 12356 2286 12368
rect 3142 12356 3148 12368
rect 2280 12328 3148 12356
rect 2280 12316 2286 12328
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2314 12220 2320 12232
rect 2179 12192 2320 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2976 12229 3004 12328
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 15102 12316 15108 12368
rect 15160 12316 15166 12368
rect 19429 12359 19487 12365
rect 19429 12356 19441 12359
rect 15948 12328 19441 12356
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5500 12260 5641 12288
rect 5500 12248 5506 12260
rect 5629 12257 5641 12260
rect 5675 12288 5687 12291
rect 6546 12288 6552 12300
rect 5675 12260 6552 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 2961 12183 3019 12189
rect 4172 12192 5365 12220
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 2792 12152 2820 12183
rect 2096 12124 2820 12152
rect 2869 12155 2927 12161
rect 2096 12112 2102 12124
rect 2314 12044 2320 12096
rect 2372 12044 2378 12096
rect 2746 12084 2774 12124
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 4172 12152 4200 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9364 12192 9781 12220
rect 9364 12180 9370 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 15948 12220 15976 12328
rect 19429 12325 19441 12328
rect 19475 12325 19487 12359
rect 19429 12319 19487 12325
rect 17954 12288 17960 12300
rect 16408 12260 17960 12288
rect 16408 12229 16436 12260
rect 17954 12248 17960 12260
rect 18012 12288 18018 12300
rect 18012 12260 18368 12288
rect 18012 12248 18018 12260
rect 12400 12192 15976 12220
rect 16393 12223 16451 12229
rect 12400 12180 12406 12192
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16942 12180 16948 12232
rect 17000 12180 17006 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 17402 12220 17408 12232
rect 17359 12192 17408 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 18340 12229 18368 12260
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 2915 12124 4200 12152
rect 10036 12155 10094 12161
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 10036 12121 10048 12155
rect 10082 12152 10094 12155
rect 10502 12152 10508 12164
rect 10082 12124 10508 12152
rect 10082 12121 10094 12124
rect 10036 12115 10094 12121
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14608 12124 14841 12152
rect 14608 12112 14614 12124
rect 14829 12121 14841 12124
rect 14875 12152 14887 12155
rect 14918 12152 14924 12164
rect 14875 12124 14924 12152
rect 14875 12121 14887 12124
rect 14829 12115 14887 12121
rect 14918 12112 14924 12124
rect 14976 12112 14982 12164
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 17862 12152 17868 12164
rect 17267 12124 17868 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 2746 12056 4077 12084
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 16301 12087 16359 12093
rect 16301 12053 16313 12087
rect 16347 12084 16359 12087
rect 17034 12084 17040 12096
rect 16347 12056 17040 12084
rect 16347 12053 16359 12056
rect 16301 12047 16359 12053
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17494 12044 17500 12096
rect 17552 12044 17558 12096
rect 18046 12044 18052 12096
rect 18104 12044 18110 12096
rect 19613 12087 19671 12093
rect 19613 12053 19625 12087
rect 19659 12084 19671 12087
rect 19702 12084 19708 12096
rect 19659 12056 19708 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 1104 11994 21043 12016
rect 1104 11942 5894 11994
rect 5946 11942 5958 11994
rect 6010 11942 6022 11994
rect 6074 11942 6086 11994
rect 6138 11942 6150 11994
rect 6202 11942 10839 11994
rect 10891 11942 10903 11994
rect 10955 11942 10967 11994
rect 11019 11942 11031 11994
rect 11083 11942 11095 11994
rect 11147 11942 15784 11994
rect 15836 11942 15848 11994
rect 15900 11942 15912 11994
rect 15964 11942 15976 11994
rect 16028 11942 16040 11994
rect 16092 11942 20729 11994
rect 20781 11942 20793 11994
rect 20845 11942 20857 11994
rect 20909 11942 20921 11994
rect 20973 11942 20985 11994
rect 21037 11942 21043 11994
rect 1104 11920 21043 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 4062 11880 4068 11892
rect 2363 11852 4068 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 2682 11812 2688 11824
rect 2148 11784 2688 11812
rect 2148 11753 2176 11784
rect 2682 11772 2688 11784
rect 2740 11772 2746 11824
rect 13280 11812 13308 11843
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 17862 11840 17868 11892
rect 17920 11840 17926 11892
rect 19337 11883 19395 11889
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19518 11880 19524 11892
rect 19383 11852 19524 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 19702 11840 19708 11892
rect 19760 11840 19766 11892
rect 14274 11812 14280 11824
rect 13280 11784 14280 11812
rect 14274 11772 14280 11784
rect 14332 11812 14338 11824
rect 14332 11784 18276 11812
rect 14332 11772 14338 11784
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 2372 11716 5273 11744
rect 2372 11704 2378 11716
rect 5261 11713 5273 11716
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5500 11716 5549 11744
rect 5500 11704 5506 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 7190 11753 7196 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6604 11716 6929 11744
rect 6604 11704 6610 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 7184 11707 7196 11753
rect 7190 11704 7196 11707
rect 7248 11704 7254 11756
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 9306 11744 9312 11756
rect 8803 11716 9312 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 12152 11747 12210 11753
rect 12152 11713 12164 11747
rect 12198 11744 12210 11747
rect 12710 11744 12716 11756
rect 12198 11716 12716 11744
rect 12198 11713 12210 11716
rect 12152 11707 12210 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 16666 11744 16672 11756
rect 14700 11716 16672 11744
rect 14700 11704 14706 11716
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 17034 11704 17040 11756
rect 17092 11704 17098 11756
rect 17144 11753 17172 11784
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17218 11704 17224 11756
rect 17276 11704 17282 11756
rect 18046 11704 18052 11756
rect 18104 11704 18110 11756
rect 18248 11753 18276 11784
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 19521 11747 19579 11753
rect 19521 11744 19533 11747
rect 19392 11716 19533 11744
rect 19392 11704 19398 11716
rect 19521 11713 19533 11716
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2866 11676 2872 11688
rect 1995 11648 2872 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 2924 11648 3893 11676
rect 2924 11636 2930 11648
rect 3881 11645 3893 11648
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 9030 11636 9036 11688
rect 9088 11636 9094 11688
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11848 11648 11897 11676
rect 11848 11636 11854 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 17494 11676 17500 11688
rect 15335 11648 17500 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 15378 11568 15384 11620
rect 15436 11568 15442 11620
rect 15473 11611 15531 11617
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 15562 11608 15568 11620
rect 15519 11580 15568 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 15841 11611 15899 11617
rect 15841 11577 15853 11611
rect 15887 11608 15899 11611
rect 16850 11608 16856 11620
rect 15887 11580 16856 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 8297 11543 8355 11549
rect 8297 11509 8309 11543
rect 8343 11540 8355 11543
rect 9122 11540 9128 11552
rect 8343 11512 9128 11540
rect 8343 11509 8355 11512
rect 8297 11503 8355 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 15013 11543 15071 11549
rect 15013 11540 15025 11543
rect 14700 11512 15025 11540
rect 14700 11500 14706 11512
rect 15013 11509 15025 11512
rect 15059 11509 15071 11543
rect 15013 11503 15071 11509
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17276 11512 18061 11540
rect 17276 11500 17282 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 1104 11450 20884 11472
rect 1104 11398 3422 11450
rect 3474 11398 3486 11450
rect 3538 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 8367 11450
rect 8419 11398 8431 11450
rect 8483 11398 8495 11450
rect 8547 11398 8559 11450
rect 8611 11398 8623 11450
rect 8675 11398 13312 11450
rect 13364 11398 13376 11450
rect 13428 11398 13440 11450
rect 13492 11398 13504 11450
rect 13556 11398 13568 11450
rect 13620 11398 18257 11450
rect 18309 11398 18321 11450
rect 18373 11398 18385 11450
rect 18437 11398 18449 11450
rect 18501 11398 18513 11450
rect 18565 11398 20884 11450
rect 1104 11376 20884 11398
rect 15286 11296 15292 11348
rect 15344 11296 15350 11348
rect 16850 11296 16856 11348
rect 16908 11296 16914 11348
rect 18785 11339 18843 11345
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 18831 11308 19625 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 2130 11228 2136 11280
rect 2188 11268 2194 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 2188 11240 4077 11268
rect 2188 11228 2194 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4065 11231 4123 11237
rect 10318 11228 10324 11280
rect 10376 11268 10382 11280
rect 10505 11271 10563 11277
rect 10505 11268 10517 11271
rect 10376 11240 10517 11268
rect 10376 11228 10382 11240
rect 10505 11237 10517 11240
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 13173 11271 13231 11277
rect 13173 11237 13185 11271
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 13188 11200 13216 11231
rect 15010 11228 15016 11280
rect 15068 11268 15074 11280
rect 15197 11271 15255 11277
rect 15197 11268 15209 11271
rect 15068 11240 15209 11268
rect 15068 11228 15074 11240
rect 15197 11237 15209 11240
rect 15243 11237 15255 11271
rect 15197 11231 15255 11237
rect 17218 11200 17224 11212
rect 13188 11172 17224 11200
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 17552 11172 18920 11200
rect 17552 11160 17558 11172
rect 1854 11092 1860 11144
rect 1912 11092 1918 11144
rect 2038 11092 2044 11144
rect 2096 11092 2102 11144
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 5500 11104 6469 11132
rect 5500 11092 5506 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9214 11132 9220 11144
rect 9171 11104 9220 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9214 11092 9220 11104
rect 9272 11132 9278 11144
rect 11790 11132 11796 11144
rect 9272 11104 11796 11132
rect 9272 11092 9278 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 17313 11135 17371 11141
rect 14056 11104 17264 11132
rect 14056 11092 14062 11104
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 5178 11067 5236 11073
rect 5178 11064 5190 11067
rect 1995 11036 5190 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 5178 11033 5190 11036
rect 5224 11033 5236 11067
rect 5178 11027 5236 11033
rect 6724 11067 6782 11073
rect 6724 11033 6736 11067
rect 6770 11064 6782 11067
rect 6822 11064 6828 11076
rect 6770 11036 6828 11064
rect 6770 11033 6782 11036
rect 6724 11027 6782 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 12066 11073 12072 11076
rect 9370 11067 9428 11073
rect 9370 11064 9382 11067
rect 8996 11036 9382 11064
rect 8996 11024 9002 11036
rect 9370 11033 9382 11036
rect 9416 11033 9428 11067
rect 9370 11027 9428 11033
rect 12060 11027 12072 11073
rect 12066 11024 12072 11027
rect 12124 11024 12130 11076
rect 14829 11067 14887 11073
rect 14829 11033 14841 11067
rect 14875 11064 14887 11067
rect 15194 11064 15200 11076
rect 14875 11036 15200 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 7834 10956 7840 11008
rect 7892 10956 7898 11008
rect 17236 11005 17264 11104
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17402 11132 17408 11144
rect 17359 11104 17408 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 18892 11141 18920 11172
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 19392 11104 19993 11132
rect 19392 11092 19398 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 19610 11024 19616 11076
rect 19668 11024 19674 11076
rect 17221 10999 17279 11005
rect 17221 10965 17233 10999
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 19426 10956 19432 11008
rect 19484 10956 19490 11008
rect 1104 10906 21043 10928
rect 1104 10854 5894 10906
rect 5946 10854 5958 10906
rect 6010 10854 6022 10906
rect 6074 10854 6086 10906
rect 6138 10854 6150 10906
rect 6202 10854 10839 10906
rect 10891 10854 10903 10906
rect 10955 10854 10967 10906
rect 11019 10854 11031 10906
rect 11083 10854 11095 10906
rect 11147 10854 15784 10906
rect 15836 10854 15848 10906
rect 15900 10854 15912 10906
rect 15964 10854 15976 10906
rect 16028 10854 16040 10906
rect 16092 10854 20729 10906
rect 20781 10854 20793 10906
rect 20845 10854 20857 10906
rect 20909 10854 20921 10906
rect 20973 10854 20985 10906
rect 21037 10854 21043 10906
rect 1104 10832 21043 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 1854 10792 1860 10804
rect 1811 10764 1860 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 15194 10792 15200 10804
rect 14108 10764 15200 10792
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 2056 10696 3801 10724
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2056 10665 2084 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 7006 10684 7012 10736
rect 7064 10724 7070 10736
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 7064 10696 7849 10724
rect 7064 10684 7070 10696
rect 7837 10693 7849 10696
rect 7883 10693 7895 10727
rect 7837 10687 7895 10693
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1912 10628 2053 10656
rect 1912 10616 1918 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2130 10616 2136 10668
rect 2188 10616 2194 10668
rect 2222 10616 2228 10668
rect 2280 10616 2286 10668
rect 14108 10665 14136 10764
rect 15194 10752 15200 10764
rect 15252 10792 15258 10804
rect 15252 10764 15332 10792
rect 15252 10752 15258 10764
rect 15010 10724 15016 10736
rect 14476 10696 15016 10724
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14231 10659 14289 10665
rect 14231 10625 14243 10659
rect 14277 10656 14289 10659
rect 14476 10656 14504 10696
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15304 10724 15332 10764
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 17865 10795 17923 10801
rect 17865 10792 17877 10795
rect 16816 10764 17877 10792
rect 16816 10752 16822 10764
rect 17865 10761 17877 10764
rect 17911 10761 17923 10795
rect 17865 10755 17923 10761
rect 17972 10764 18276 10792
rect 17034 10724 17040 10736
rect 15304 10696 17040 10724
rect 15304 10665 15332 10696
rect 17034 10684 17040 10696
rect 17092 10724 17098 10736
rect 17092 10696 17172 10724
rect 17092 10684 17098 10696
rect 14277 10628 14504 10656
rect 14553 10659 14611 10665
rect 14277 10625 14289 10628
rect 14231 10619 14289 10625
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 14553 10619 14611 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 4212 10560 5181 10588
rect 4212 10548 4218 10560
rect 5169 10557 5181 10560
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5442 10588 5448 10600
rect 5316 10560 5448 10588
rect 5316 10548 5322 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 14568 10588 14596 10619
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 17144 10665 17172 10696
rect 17770 10684 17776 10736
rect 17828 10724 17834 10736
rect 17972 10724 18000 10764
rect 18046 10733 18052 10736
rect 17828 10696 18000 10724
rect 18033 10727 18052 10733
rect 17828 10684 17834 10696
rect 18033 10693 18045 10727
rect 18033 10687 18052 10693
rect 18046 10684 18052 10687
rect 18104 10684 18110 10736
rect 18248 10733 18276 10764
rect 19334 10752 19340 10804
rect 19392 10752 19398 10804
rect 18233 10727 18291 10733
rect 18233 10693 18245 10727
rect 18279 10693 18291 10727
rect 18233 10687 18291 10693
rect 18690 10684 18696 10736
rect 18748 10724 18754 10736
rect 18748 10696 19472 10724
rect 18748 10684 18754 10696
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 15528 10628 15577 10656
rect 15528 10616 15534 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17368 10628 17417 10656
rect 17368 10616 17374 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 19444 10665 19472 10696
rect 19245 10659 19303 10665
rect 19245 10656 19257 10659
rect 17552 10628 19257 10656
rect 17552 10616 17558 10628
rect 19245 10625 19257 10628
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 19429 10659 19487 10665
rect 19429 10625 19441 10659
rect 19475 10656 19487 10659
rect 20070 10656 20076 10668
rect 19475 10628 20076 10656
rect 19475 10625 19487 10628
rect 19429 10619 19487 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 14568 10560 14688 10588
rect 14660 10520 14688 10560
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15160 10560 16988 10588
rect 15160 10548 15166 10560
rect 16853 10523 16911 10529
rect 16853 10520 16865 10523
rect 14660 10492 16865 10520
rect 16853 10489 16865 10492
rect 16899 10489 16911 10523
rect 16960 10520 16988 10560
rect 17328 10520 17356 10616
rect 17770 10548 17776 10600
rect 17828 10588 17834 10600
rect 19610 10588 19616 10600
rect 17828 10560 19616 10588
rect 17828 10548 17834 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 16960 10492 17356 10520
rect 16853 10483 16911 10489
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14240 10424 14381 10452
rect 14240 10412 14246 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14369 10415 14427 10421
rect 14458 10412 14464 10464
rect 14516 10412 14522 10464
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14608 10424 15025 10452
rect 14608 10412 14614 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10452 15531 10455
rect 15654 10452 15660 10464
rect 15519 10424 15660 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 17218 10412 17224 10464
rect 17276 10412 17282 10464
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10452 18107 10455
rect 18690 10452 18696 10464
rect 18095 10424 18696 10452
rect 18095 10421 18107 10424
rect 18049 10415 18107 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 1104 10362 20884 10384
rect 1104 10310 3422 10362
rect 3474 10310 3486 10362
rect 3538 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 8367 10362
rect 8419 10310 8431 10362
rect 8483 10310 8495 10362
rect 8547 10310 8559 10362
rect 8611 10310 8623 10362
rect 8675 10310 13312 10362
rect 13364 10310 13376 10362
rect 13428 10310 13440 10362
rect 13492 10310 13504 10362
rect 13556 10310 13568 10362
rect 13620 10310 18257 10362
rect 18309 10310 18321 10362
rect 18373 10310 18385 10362
rect 18437 10310 18449 10362
rect 18501 10310 18513 10362
rect 18565 10310 20884 10362
rect 1104 10288 20884 10310
rect 2038 10208 2044 10260
rect 2096 10208 2102 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 15194 10248 15200 10260
rect 14240 10220 15200 10248
rect 14240 10208 14246 10220
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 17552 10220 17601 10248
rect 17552 10208 17558 10220
rect 17589 10217 17601 10220
rect 17635 10217 17647 10251
rect 17589 10211 17647 10217
rect 13265 10183 13323 10189
rect 13265 10149 13277 10183
rect 13311 10180 13323 10183
rect 13311 10152 17540 10180
rect 13311 10149 13323 10152
rect 13265 10143 13323 10149
rect 1946 10112 1952 10124
rect 1780 10084 1952 10112
rect 1780 10053 1808 10084
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9364 10084 10057 10112
rect 9364 10072 9370 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11848 10084 11897 10112
rect 11848 10072 11854 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15102 10112 15108 10124
rect 14875 10084 15108 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15286 10072 15292 10124
rect 15344 10072 15350 10124
rect 17512 10121 17540 10152
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10081 17555 10115
rect 17497 10075 17555 10081
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 2130 10044 2136 10056
rect 2087 10016 2136 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 15028 10016 15976 10044
rect 5258 9936 5264 9988
rect 5316 9936 5322 9988
rect 10312 9979 10370 9985
rect 10312 9945 10324 9979
rect 10358 9976 10370 9979
rect 10594 9976 10600 9988
rect 10358 9948 10600 9976
rect 10358 9945 10370 9948
rect 10312 9939 10370 9945
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 12152 9979 12210 9985
rect 12152 9945 12164 9979
rect 12198 9976 12210 9979
rect 15028 9976 15056 10016
rect 12198 9948 15056 9976
rect 12198 9945 12210 9948
rect 12152 9939 12210 9945
rect 15194 9936 15200 9988
rect 15252 9936 15258 9988
rect 15948 9976 15976 10016
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 17092 10016 17233 10044
rect 17092 10004 17098 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17604 10044 17632 10211
rect 19978 10208 19984 10260
rect 20036 10208 20042 10260
rect 19242 10140 19248 10192
rect 19300 10180 19306 10192
rect 19429 10183 19487 10189
rect 19429 10180 19441 10183
rect 19300 10152 19441 10180
rect 19300 10140 19306 10152
rect 19429 10149 19441 10152
rect 19475 10149 19487 10183
rect 19429 10143 19487 10149
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 17604 10016 18705 10044
rect 17221 10007 17279 10013
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 19610 10004 19616 10056
rect 19668 10044 19674 10056
rect 19705 10047 19763 10053
rect 19705 10044 19717 10047
rect 19668 10016 19717 10044
rect 19668 10004 19674 10016
rect 19705 10013 19717 10016
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19334 9976 19340 9988
rect 15948 9948 19340 9976
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 11422 9868 11428 9920
rect 11480 9868 11486 9920
rect 14645 9911 14703 9917
rect 14645 9877 14657 9911
rect 14691 9908 14703 9911
rect 15102 9908 15108 9920
rect 14691 9880 15108 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 18785 9911 18843 9917
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 18831 9880 19625 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 19794 9868 19800 9920
rect 19852 9868 19858 9920
rect 1104 9818 21043 9840
rect 1104 9766 5894 9818
rect 5946 9766 5958 9818
rect 6010 9766 6022 9818
rect 6074 9766 6086 9818
rect 6138 9766 6150 9818
rect 6202 9766 10839 9818
rect 10891 9766 10903 9818
rect 10955 9766 10967 9818
rect 11019 9766 11031 9818
rect 11083 9766 11095 9818
rect 11147 9766 15784 9818
rect 15836 9766 15848 9818
rect 15900 9766 15912 9818
rect 15964 9766 15976 9818
rect 16028 9766 16040 9818
rect 16092 9766 20729 9818
rect 20781 9766 20793 9818
rect 20845 9766 20857 9818
rect 20909 9766 20921 9818
rect 20973 9766 20985 9818
rect 21037 9766 21043 9818
rect 1104 9744 21043 9766
rect 5258 9704 5264 9716
rect 4632 9676 5264 9704
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4632 9509 4660 9676
rect 5258 9664 5264 9676
rect 5316 9704 5322 9716
rect 6546 9704 6552 9716
rect 5316 9676 6552 9704
rect 5316 9664 5322 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 19613 9707 19671 9713
rect 14660 9676 14964 9704
rect 14660 9636 14688 9676
rect 14108 9608 14688 9636
rect 14108 9580 14136 9608
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14792 9608 14841 9636
rect 14792 9596 14798 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 14936 9636 14964 9676
rect 19613 9673 19625 9707
rect 19659 9704 19671 9707
rect 19794 9704 19800 9716
rect 19659 9676 19800 9704
rect 19659 9673 19671 9676
rect 19613 9667 19671 9673
rect 19794 9664 19800 9676
rect 19852 9664 19858 9716
rect 20070 9664 20076 9716
rect 20128 9664 20134 9716
rect 14936 9608 16252 9636
rect 14829 9599 14887 9605
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 4873 9571 4931 9577
rect 4873 9568 4885 9571
rect 4764 9540 4885 9568
rect 4764 9528 4770 9540
rect 4873 9537 4885 9540
rect 4919 9537 4931 9571
rect 4873 9531 4931 9537
rect 8317 9571 8375 9577
rect 8317 9537 8329 9571
rect 8363 9568 8375 9571
rect 8846 9568 8852 9580
rect 8363 9540 8852 9568
rect 8363 9537 8375 9540
rect 8317 9531 8375 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 9214 9528 9220 9580
rect 9272 9568 9278 9580
rect 9657 9571 9715 9577
rect 9657 9568 9669 9571
rect 9272 9540 9669 9568
rect 9272 9528 9278 9540
rect 9657 9537 9669 9540
rect 9703 9537 9715 9571
rect 9657 9531 9715 9537
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 12158 9577 12164 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11848 9540 11897 9568
rect 11848 9528 11854 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12152 9531 12164 9577
rect 12158 9528 12164 9531
rect 12216 9528 12222 9580
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 14976 9571 15034 9577
rect 14976 9568 14988 9571
rect 14516 9540 14988 9568
rect 14516 9528 14522 9540
rect 14976 9537 14988 9540
rect 15022 9537 15034 9571
rect 16224 9568 16252 9608
rect 17126 9596 17132 9648
rect 17184 9636 17190 9648
rect 19150 9636 19156 9648
rect 17184 9608 19156 9636
rect 17184 9596 17190 9608
rect 19150 9596 19156 9608
rect 19208 9636 19214 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 19208 9608 19257 9636
rect 19208 9596 19214 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19445 9639 19503 9645
rect 19445 9636 19457 9639
rect 19245 9599 19303 9605
rect 19352 9608 19457 9636
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 16224 9540 17233 9568
rect 14976 9531 15034 9537
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4028 9472 4629 9500
rect 4028 9460 4034 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 8754 9500 8760 9512
rect 8619 9472 8760 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 8754 9460 8760 9472
rect 8812 9500 8818 9512
rect 9306 9500 9312 9512
rect 8812 9472 9312 9500
rect 8812 9460 8818 9472
rect 9306 9460 9312 9472
rect 9364 9500 9370 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9364 9472 9413 9500
rect 9364 9460 9370 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14550 9500 14556 9512
rect 14415 9472 14556 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 15197 9503 15255 9509
rect 15197 9500 15209 9503
rect 14752 9472 15209 9500
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 14277 9435 14335 9441
rect 6043 9404 7696 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 7466 9364 7472 9376
rect 7239 9336 7472 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 7668 9364 7696 9404
rect 14277 9401 14289 9435
rect 14323 9432 14335 9435
rect 14752 9432 14780 9472
rect 15197 9469 15209 9472
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 14323 9404 14780 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 15102 9392 15108 9444
rect 15160 9392 15166 9444
rect 9766 9364 9772 9376
rect 7668 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 10744 9336 10793 9364
rect 10744 9324 10750 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13814 9364 13820 9376
rect 13311 9336 13820 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 15286 9364 15292 9376
rect 14516 9336 15292 9364
rect 14516 9324 14522 9336
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 16776 9364 16804 9540
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 17552 9540 17601 9568
rect 17552 9528 17558 9540
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17313 9503 17371 9509
rect 16908 9492 17172 9500
rect 17313 9492 17325 9503
rect 16908 9472 17325 9492
rect 16908 9460 16914 9472
rect 17144 9469 17325 9472
rect 17359 9469 17371 9503
rect 17144 9464 17371 9469
rect 17313 9463 17371 9464
rect 17328 9432 17356 9463
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19352 9500 19380 9608
rect 19445 9605 19457 9608
rect 19491 9605 19503 9639
rect 19812 9636 19840 9664
rect 19812 9608 20300 9636
rect 19445 9599 19503 9605
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 20272 9577 20300 9608
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19668 9540 20085 9568
rect 19668 9528 19674 9540
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 19300 9472 19380 9500
rect 19300 9460 19306 9472
rect 17586 9432 17592 9444
rect 17328 9404 17592 9432
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 17865 9435 17923 9441
rect 17865 9401 17877 9435
rect 17911 9432 17923 9435
rect 18046 9432 18052 9444
rect 17911 9404 18052 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 16776 9336 19441 9364
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 1104 9274 20884 9296
rect 1104 9222 3422 9274
rect 3474 9222 3486 9274
rect 3538 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 8367 9274
rect 8419 9222 8431 9274
rect 8483 9222 8495 9274
rect 8547 9222 8559 9274
rect 8611 9222 8623 9274
rect 8675 9222 13312 9274
rect 13364 9222 13376 9274
rect 13428 9222 13440 9274
rect 13492 9222 13504 9274
rect 13556 9222 13568 9274
rect 13620 9222 18257 9274
rect 18309 9222 18321 9274
rect 18373 9222 18385 9274
rect 18437 9222 18449 9274
rect 18501 9222 18513 9274
rect 18565 9222 20884 9274
rect 1104 9200 20884 9222
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8938 9160 8944 9172
rect 8527 9132 8944 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 14553 9163 14611 9169
rect 14553 9160 14565 9163
rect 14332 9132 14565 9160
rect 14332 9120 14338 9132
rect 14553 9129 14565 9132
rect 14599 9129 14611 9163
rect 14553 9123 14611 9129
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17494 9160 17500 9172
rect 17092 9132 17500 9160
rect 17092 9120 17098 9132
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 19521 9163 19579 9169
rect 19521 9160 19533 9163
rect 17736 9132 19533 9160
rect 17736 9120 17742 9132
rect 19521 9129 19533 9132
rect 19567 9129 19579 9163
rect 19521 9123 19579 9129
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 17586 9092 17592 9104
rect 10560 9064 17592 9092
rect 10560 9052 10566 9064
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 2130 8984 2136 9036
rect 2188 8984 2194 9036
rect 3970 8984 3976 9036
rect 4028 8984 4034 9036
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 9024 7987 9027
rect 8754 9024 8760 9036
rect 7975 8996 8760 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14608 8996 14657 9024
rect 14608 8984 14614 8996
rect 14645 8993 14657 8996
rect 14691 9024 14703 9027
rect 15010 9024 15016 9036
rect 14691 8996 15016 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 17696 9024 17724 9120
rect 17052 8996 17724 9024
rect 2406 8916 2412 8968
rect 2464 8916 2470 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 6788 8928 8401 8956
rect 6788 8916 6794 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8938 8956 8944 8968
rect 8619 8928 8944 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9548 8928 14688 8956
rect 9548 8916 9554 8928
rect 14660 8900 14688 8928
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 16942 8916 16948 8968
rect 17000 8916 17006 8968
rect 17052 8956 17080 8996
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19300 8996 19656 9024
rect 19300 8984 19306 8996
rect 17108 8959 17166 8965
rect 17108 8956 17120 8959
rect 17052 8928 17120 8956
rect 17108 8925 17120 8928
rect 17154 8925 17166 8959
rect 17108 8919 17166 8925
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8958 17371 8959
rect 17494 8958 17500 8968
rect 17359 8930 17500 8958
rect 17359 8925 17371 8930
rect 17313 8919 17371 8925
rect 4240 8891 4298 8897
rect 4240 8857 4252 8891
rect 4286 8888 4298 8891
rect 4522 8888 4528 8900
rect 4286 8860 4528 8888
rect 4286 8857 4298 8860
rect 4240 8851 4298 8857
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 7662 8891 7720 8897
rect 7662 8888 7674 8891
rect 5776 8860 7674 8888
rect 5776 8848 5782 8860
rect 7662 8857 7674 8860
rect 7708 8857 7720 8891
rect 7662 8851 7720 8857
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 14056 8860 14565 8888
rect 14056 8848 14062 8860
rect 14553 8857 14565 8860
rect 14599 8857 14611 8891
rect 14553 8851 14611 8857
rect 14642 8848 14648 8900
rect 14700 8888 14706 8900
rect 14700 8860 15148 8888
rect 14700 8848 14706 8860
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1854 8820 1860 8832
rect 1627 8792 1860 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 5353 8823 5411 8829
rect 5353 8820 5365 8823
rect 4856 8792 5365 8820
rect 4856 8780 4862 8792
rect 5353 8789 5365 8792
rect 5399 8789 5411 8823
rect 5353 8783 5411 8789
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6420 8792 6561 8820
rect 6420 8780 6426 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 15010 8780 15016 8832
rect 15068 8780 15074 8832
rect 15120 8820 15148 8860
rect 15286 8848 15292 8900
rect 15344 8888 15350 8900
rect 16574 8888 16580 8900
rect 15344 8860 16580 8888
rect 15344 8848 15350 8860
rect 16574 8848 16580 8860
rect 16632 8888 16638 8900
rect 17236 8888 17264 8919
rect 16632 8860 17264 8888
rect 16632 8848 16638 8860
rect 17328 8820 17356 8919
rect 17494 8916 17500 8930
rect 17552 8916 17558 8968
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 19628 8965 19656 8996
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19208 8928 19441 8956
rect 19208 8916 19214 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 15120 8792 17356 8820
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17862 8820 17868 8832
rect 17635 8792 17868 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 1104 8730 21043 8752
rect 1104 8678 5894 8730
rect 5946 8678 5958 8730
rect 6010 8678 6022 8730
rect 6074 8678 6086 8730
rect 6138 8678 6150 8730
rect 6202 8678 10839 8730
rect 10891 8678 10903 8730
rect 10955 8678 10967 8730
rect 11019 8678 11031 8730
rect 11083 8678 11095 8730
rect 11147 8678 15784 8730
rect 15836 8678 15848 8730
rect 15900 8678 15912 8730
rect 15964 8678 15976 8730
rect 16028 8678 16040 8730
rect 16092 8678 20729 8730
rect 20781 8678 20793 8730
rect 20845 8678 20857 8730
rect 20909 8678 20921 8730
rect 20973 8678 20985 8730
rect 21037 8678 21043 8730
rect 1104 8656 21043 8678
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 4154 8616 4160 8628
rect 2547 8588 4160 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4706 8616 4712 8628
rect 4663 8588 4712 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 7190 8616 7196 8628
rect 5307 8588 7196 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 12216 8588 12265 8616
rect 12216 8576 12222 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 17644 8588 19533 8616
rect 17644 8576 17650 8588
rect 19521 8585 19533 8588
rect 19567 8585 19579 8619
rect 19521 8579 19579 8585
rect 19628 8588 19932 8616
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5905 8551 5963 8557
rect 5905 8548 5917 8551
rect 5592 8520 5917 8548
rect 5592 8508 5598 8520
rect 5905 8517 5917 8520
rect 5951 8548 5963 8551
rect 6794 8551 6852 8557
rect 6794 8548 6806 8551
rect 5951 8520 6806 8548
rect 5951 8517 5963 8520
rect 5905 8511 5963 8517
rect 6794 8517 6806 8520
rect 6840 8517 6852 8551
rect 6794 8511 6852 8517
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 14458 8548 14464 8560
rect 9640 8520 14464 8548
rect 9640 8508 9646 8520
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 14918 8548 14924 8560
rect 14568 8520 14924 8548
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 2004 8452 2053 8480
rect 2004 8440 2010 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4522 8480 4528 8492
rect 4479 8452 4528 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5626 8480 5632 8492
rect 5399 8452 5632 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 7944 8452 8401 8480
rect 2038 8304 2044 8356
rect 2096 8344 2102 8356
rect 7944 8353 7972 8452
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 14568 8489 14596 8520
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 16724 8520 18061 8548
rect 16724 8508 16730 8520
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 12406 8384 12541 8412
rect 2133 8347 2191 8353
rect 2133 8344 2145 8347
rect 2096 8316 2145 8344
rect 2096 8304 2102 8316
rect 2133 8313 2145 8316
rect 2179 8313 2191 8347
rect 2133 8307 2191 8313
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8313 7987 8347
rect 7929 8307 7987 8313
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8276 8539 8279
rect 8754 8276 8760 8288
rect 8527 8248 8760 8276
rect 8527 8245 8539 8248
rect 8481 8239 8539 8245
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 12406 8276 12434 8384
rect 12529 8381 12541 8384
rect 12575 8412 12587 8415
rect 13722 8412 13728 8424
rect 12575 8384 13728 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 11020 8248 12434 8276
rect 11020 8236 11026 8248
rect 12618 8236 12624 8288
rect 12676 8236 12682 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 14568 8276 14596 8443
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14829 8483 14887 8489
rect 14829 8480 14841 8483
rect 14700 8452 14841 8480
rect 14700 8440 14706 8452
rect 14829 8449 14841 8452
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 16908 8452 17141 8480
rect 16908 8440 16914 8452
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 14792 8384 15209 8412
rect 14792 8372 14798 8384
rect 15197 8381 15209 8384
rect 15243 8412 15255 8415
rect 17034 8412 17040 8424
rect 15243 8384 17040 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 17236 8412 17264 8520
rect 18049 8517 18061 8520
rect 18095 8517 18107 8551
rect 19242 8548 19248 8560
rect 18049 8511 18107 8517
rect 18892 8520 19248 8548
rect 18892 8492 18920 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 19628 8548 19656 8588
rect 19392 8520 19656 8548
rect 19689 8551 19747 8557
rect 19392 8508 19398 8520
rect 19689 8517 19701 8551
rect 19735 8548 19747 8551
rect 19794 8548 19800 8560
rect 19735 8520 19800 8548
rect 19735 8517 19747 8520
rect 19689 8511 19747 8517
rect 19794 8508 19800 8520
rect 19852 8508 19858 8560
rect 19904 8557 19932 8588
rect 19889 8551 19947 8557
rect 19889 8517 19901 8551
rect 19935 8517 19947 8551
rect 19889 8511 19947 8517
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17862 8480 17868 8492
rect 17368 8452 17868 8480
rect 17368 8440 17374 8452
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 17236 8384 17417 8412
rect 17405 8381 17417 8384
rect 17451 8412 17463 8415
rect 17586 8412 17592 8424
rect 17451 8384 17592 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18156 8412 18184 8443
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19107 8452 19656 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19628 8424 19656 8452
rect 17736 8384 18184 8412
rect 17736 8372 17742 8384
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 17184 8316 17325 8344
rect 17184 8304 17190 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 18969 8347 19027 8353
rect 18969 8313 18981 8347
rect 19015 8344 19027 8347
rect 19015 8316 19748 8344
rect 19015 8313 19027 8316
rect 18969 8307 19027 8313
rect 12860 8248 14596 8276
rect 17865 8279 17923 8285
rect 12860 8236 12866 8248
rect 17865 8245 17877 8279
rect 17911 8276 17923 8279
rect 17954 8276 17960 8288
rect 17911 8248 17960 8276
rect 17911 8245 17923 8248
rect 17865 8239 17923 8245
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 19720 8285 19748 8316
rect 19705 8279 19763 8285
rect 19705 8245 19717 8279
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 1104 8186 20884 8208
rect 1104 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 8367 8186
rect 8419 8134 8431 8186
rect 8483 8134 8495 8186
rect 8547 8134 8559 8186
rect 8611 8134 8623 8186
rect 8675 8134 13312 8186
rect 13364 8134 13376 8186
rect 13428 8134 13440 8186
rect 13492 8134 13504 8186
rect 13556 8134 13568 8186
rect 13620 8134 18257 8186
rect 18309 8134 18321 8186
rect 18373 8134 18385 8186
rect 18437 8134 18449 8186
rect 18501 8134 18513 8186
rect 18565 8134 20884 8186
rect 1104 8112 20884 8134
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2314 8072 2320 8084
rect 2271 8044 2320 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 5718 8072 5724 8084
rect 4755 8044 5724 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7009 8075 7067 8081
rect 7009 8072 7021 8075
rect 6972 8044 7021 8072
rect 6972 8032 6978 8044
rect 7009 8041 7021 8044
rect 7055 8041 7067 8075
rect 7009 8035 7067 8041
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8846 8072 8852 8084
rect 8435 8044 8852 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 9088 8044 9229 8072
rect 9088 8032 9094 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10652 8044 10701 8072
rect 10652 8032 10658 8044
rect 10689 8041 10701 8044
rect 10735 8041 10747 8075
rect 12437 8075 12495 8081
rect 10689 8035 10747 8041
rect 10796 8044 11284 8072
rect 8478 7964 8484 8016
rect 8536 8004 8542 8016
rect 10796 8004 10824 8044
rect 8536 7976 10824 8004
rect 8536 7964 8542 7976
rect 10962 7964 10968 8016
rect 11020 7964 11026 8016
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4614 7936 4620 7948
rect 4111 7908 4620 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4614 7896 4620 7908
rect 4672 7936 4678 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4672 7908 5181 7936
rect 4672 7896 4678 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7936 9367 7939
rect 10226 7936 10232 7948
rect 9355 7908 10232 7936
rect 9355 7905 9367 7908
rect 9309 7899 9367 7905
rect 10226 7896 10232 7908
rect 10284 7936 10290 7948
rect 10980 7936 11008 7964
rect 11256 7936 11284 8044
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12483 8044 12517 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 12452 8004 12480 8035
rect 12618 8032 12624 8084
rect 12676 8032 12682 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13228 8044 13277 8072
rect 13228 8032 13234 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 14642 8032 14648 8084
rect 14700 8032 14706 8084
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 15378 8072 15384 8084
rect 15151 8044 15384 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 15378 8032 15384 8044
rect 15436 8072 15442 8084
rect 16114 8072 16120 8084
rect 15436 8044 16120 8072
rect 15436 8032 15442 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16485 8075 16543 8081
rect 16485 8041 16497 8075
rect 16531 8041 16543 8075
rect 16485 8035 16543 8041
rect 12802 8004 12808 8016
rect 12400 7976 12808 8004
rect 12400 7964 12406 7976
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 16500 8004 16528 8035
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17092 8044 17325 8072
rect 17092 8032 17098 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 18874 8032 18880 8084
rect 18932 8032 18938 8084
rect 19794 8032 19800 8084
rect 19852 8032 19858 8084
rect 13004 7976 16528 8004
rect 16577 8007 16635 8013
rect 12618 7936 12624 7948
rect 10284 7908 11192 7936
rect 10284 7896 10290 7908
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 2038 7868 2044 7880
rect 1995 7840 2044 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4706 7868 4712 7880
rect 4571 7840 4712 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 2240 7800 2268 7828
rect 1820 7772 2268 7800
rect 4448 7800 4476 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7868 5411 7871
rect 5534 7868 5540 7880
rect 5399 7840 5540 7868
rect 5399 7837 5411 7840
rect 5353 7831 5411 7837
rect 5368 7800 5396 7831
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6052 7840 6377 7868
rect 6052 7828 6058 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 4448 7772 5396 7800
rect 6380 7800 6408 7831
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6512 7840 6561 7868
rect 6512 7828 6518 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6696 7840 6837 7868
rect 6696 7828 6702 7840
rect 6825 7837 6837 7840
rect 6871 7868 6883 7871
rect 8021 7871 8079 7877
rect 6871 7840 7512 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7374 7800 7380 7812
rect 6380 7772 7380 7800
rect 1820 7760 1826 7772
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 7484 7800 7512 7840
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8294 7868 8300 7880
rect 8067 7840 8300 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8294 7828 8300 7840
rect 8352 7868 8358 7880
rect 8938 7868 8944 7880
rect 8352 7840 8944 7868
rect 8352 7828 8358 7840
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9858 7868 9864 7880
rect 9447 7840 9864 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10652 7840 10885 7868
rect 10652 7828 10658 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11054 7868 11060 7880
rect 11011 7840 11060 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11164 7877 11192 7908
rect 11256 7908 12624 7936
rect 11256 7877 11284 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 13004 7868 13032 7976
rect 16577 7973 16589 8007
rect 16623 8004 16635 8007
rect 17129 8007 17187 8013
rect 17129 8004 17141 8007
rect 16623 7976 17141 8004
rect 16623 7973 16635 7976
rect 16577 7967 16635 7973
rect 17129 7973 17141 7976
rect 17175 7973 17187 8007
rect 17129 7967 17187 7973
rect 17586 7964 17592 8016
rect 17644 8004 17650 8016
rect 18693 8007 18751 8013
rect 18693 8004 18705 8007
rect 17644 7976 18705 8004
rect 17644 7964 17650 7976
rect 18693 7973 18705 7976
rect 18739 7973 18751 8007
rect 18693 7967 18751 7973
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13320 7908 13369 7936
rect 13320 7896 13326 7908
rect 13357 7905 13369 7908
rect 13403 7936 13415 7939
rect 13630 7936 13636 7948
rect 13403 7908 13636 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 15654 7936 15660 7948
rect 14967 7908 15660 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 12124 7840 13032 7868
rect 13081 7871 13139 7877
rect 12124 7828 12130 7840
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 8205 7803 8263 7809
rect 8205 7800 8217 7803
rect 7484 7772 8217 7800
rect 8205 7769 8217 7772
rect 8251 7800 8263 7803
rect 9214 7800 9220 7812
rect 8251 7772 9220 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 9674 7760 9680 7812
rect 9732 7760 9738 7812
rect 12250 7800 12256 7812
rect 10152 7772 12256 7800
rect 10152 7744 10180 7772
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 12434 7760 12440 7812
rect 12492 7809 12498 7812
rect 12492 7803 12527 7809
rect 12515 7800 12527 7803
rect 13096 7800 13124 7831
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 14936 7868 14964 7899
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 16393 7939 16451 7945
rect 16393 7905 16405 7939
rect 16439 7936 16451 7939
rect 16482 7936 16488 7948
rect 16439 7908 16488 7936
rect 16439 7905 16451 7908
rect 16393 7899 16451 7905
rect 13596 7840 14964 7868
rect 15197 7871 15255 7877
rect 13596 7828 13602 7840
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15286 7868 15292 7880
rect 15243 7840 15292 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 12515 7772 13124 7800
rect 12515 7769 12527 7772
rect 12492 7763 12527 7769
rect 12492 7760 12498 7763
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 16408 7800 16436 7899
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18417 7939 18475 7945
rect 18417 7936 18429 7939
rect 18196 7908 18429 7936
rect 18196 7896 18202 7908
rect 18417 7905 18429 7908
rect 18463 7905 18475 7939
rect 18417 7899 18475 7905
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17954 7868 17960 7880
rect 16715 7840 17960 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 18932 7840 19441 7868
rect 18932 7828 18938 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 17310 7809 17316 7812
rect 13780 7772 16436 7800
rect 17297 7803 17316 7809
rect 13780 7760 13786 7772
rect 17297 7769 17309 7803
rect 17297 7763 17316 7769
rect 17310 7760 17316 7763
rect 17368 7760 17374 7812
rect 17497 7803 17555 7809
rect 17497 7769 17509 7803
rect 17543 7800 17555 7803
rect 17586 7800 17592 7812
rect 17543 7772 17592 7800
rect 17543 7769 17555 7772
rect 17497 7763 17555 7769
rect 17586 7760 17592 7772
rect 17644 7760 17650 7812
rect 19610 7760 19616 7812
rect 19668 7760 19674 7812
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 2004 7704 2053 7732
rect 2004 7692 2010 7704
rect 2041 7701 2053 7704
rect 2087 7732 2099 7735
rect 2130 7732 2136 7744
rect 2087 7704 2136 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2130 7692 2136 7704
rect 2188 7732 2194 7744
rect 3142 7732 3148 7744
rect 2188 7704 3148 7732
rect 2188 7692 2194 7704
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 5537 7735 5595 7741
rect 5537 7732 5549 7735
rect 4764 7704 5549 7732
rect 4764 7692 4770 7704
rect 5537 7701 5549 7704
rect 5583 7732 5595 7735
rect 6638 7732 6644 7744
rect 5583 7704 6644 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 9585 7735 9643 7741
rect 9585 7701 9597 7735
rect 9631 7732 9643 7735
rect 10134 7732 10140 7744
rect 9631 7704 10140 7732
rect 9631 7701 9643 7704
rect 9585 7695 9643 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 17678 7732 17684 7744
rect 12676 7704 17684 7732
rect 12676 7692 12682 7704
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 1104 7642 21043 7664
rect 1104 7590 5894 7642
rect 5946 7590 5958 7642
rect 6010 7590 6022 7642
rect 6074 7590 6086 7642
rect 6138 7590 6150 7642
rect 6202 7590 10839 7642
rect 10891 7590 10903 7642
rect 10955 7590 10967 7642
rect 11019 7590 11031 7642
rect 11083 7590 11095 7642
rect 11147 7590 15784 7642
rect 15836 7590 15848 7642
rect 15900 7590 15912 7642
rect 15964 7590 15976 7642
rect 16028 7590 16040 7642
rect 16092 7590 20729 7642
rect 20781 7590 20793 7642
rect 20845 7590 20857 7642
rect 20909 7590 20921 7642
rect 20973 7590 20985 7642
rect 21037 7590 21043 7642
rect 1104 7568 21043 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 2832 7500 4905 7528
rect 2832 7488 2838 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 2958 7420 2964 7472
rect 3016 7420 3022 7472
rect 4908 7460 4936 7491
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5684 7500 5733 7528
rect 5684 7488 5690 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 8294 7528 8300 7540
rect 7515 7500 8300 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10594 7528 10600 7540
rect 10091 7500 10600 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 12250 7528 12256 7540
rect 12207 7500 12256 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 13228 7500 13369 7528
rect 13228 7488 13234 7500
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13357 7491 13415 7497
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13722 7528 13728 7540
rect 13587 7500 13728 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 15378 7528 15384 7540
rect 13832 7500 15384 7528
rect 9490 7460 9496 7472
rect 4908 7432 5764 7460
rect 5736 7404 5764 7432
rect 8312 7432 9496 7460
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5258 7392 5264 7404
rect 5215 7364 5264 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6454 7392 6460 7404
rect 5951 7364 6460 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6638 7392 6644 7404
rect 6595 7364 6644 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6564 7324 6592 7355
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7248 7364 7297 7392
rect 7248 7352 7254 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 8312 7401 8340 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 9861 7463 9919 7469
rect 9861 7460 9873 7463
rect 9732 7432 9873 7460
rect 9732 7420 9738 7432
rect 9861 7429 9873 7432
rect 9907 7460 9919 7463
rect 9907 7432 12112 7460
rect 9907 7429 9919 7432
rect 9861 7423 9919 7429
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7432 7364 7481 7392
rect 7432 7352 7438 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8754 7392 8760 7404
rect 8619 7364 8760 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 12084 7401 12112 7432
rect 10781 7395 10839 7401
rect 10781 7392 10793 7395
rect 10744 7364 10793 7392
rect 10744 7352 10750 7364
rect 10781 7361 10793 7364
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12268 7392 12296 7488
rect 12342 7420 12348 7472
rect 12400 7420 12406 7472
rect 13832 7460 13860 7500
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 17770 7528 17776 7540
rect 17543 7500 17776 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 17770 7488 17776 7500
rect 17828 7528 17834 7540
rect 19334 7528 19340 7540
rect 17828 7500 19340 7528
rect 17828 7488 17834 7500
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 15194 7460 15200 7472
rect 13372 7432 13860 7460
rect 14016 7432 15200 7460
rect 13372 7392 13400 7432
rect 13538 7392 13544 7404
rect 12268 7364 13400 7392
rect 13464 7364 13544 7392
rect 12069 7355 12127 7361
rect 6144 7296 6592 7324
rect 6144 7284 6150 7296
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 8496 7324 8524 7352
rect 9030 7324 9036 7336
rect 8496 7296 9036 7324
rect 6825 7287 6883 7293
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 12084 7324 12112 7355
rect 12250 7324 12256 7336
rect 12084 7296 12256 7324
rect 12250 7284 12256 7296
rect 12308 7324 12314 7336
rect 12434 7324 12440 7336
rect 12308 7296 12440 7324
rect 12308 7284 12314 7296
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13464 7324 13492 7364
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 14016 7401 14044 7432
rect 15194 7420 15200 7432
rect 15252 7460 15258 7472
rect 15749 7463 15807 7469
rect 15749 7460 15761 7463
rect 15252 7432 15761 7460
rect 15252 7420 15258 7432
rect 15749 7429 15761 7432
rect 15795 7429 15807 7463
rect 15749 7423 15807 7429
rect 16482 7420 16488 7472
rect 16540 7460 16546 7472
rect 16540 7432 17356 7460
rect 16540 7420 16546 7432
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15344 7364 15669 7392
rect 15344 7352 15350 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 17328 7401 17356 7432
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16172 7364 17049 7392
rect 16172 7352 16178 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 12860 7296 13492 7324
rect 12860 7284 12866 7296
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13872 7296 14841 7324
rect 13872 7284 13878 7296
rect 14829 7293 14841 7296
rect 14875 7324 14887 7327
rect 15010 7324 15016 7336
rect 14875 7296 15016 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7256 8447 7259
rect 9582 7256 9588 7268
rect 8435 7228 9588 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 9858 7216 9864 7268
rect 9916 7216 9922 7268
rect 12345 7259 12403 7265
rect 12345 7225 12357 7259
rect 12391 7256 12403 7259
rect 12526 7256 12532 7268
rect 12391 7228 12532 7256
rect 12391 7225 12403 7228
rect 12345 7219 12403 7225
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 14918 7216 14924 7268
rect 14976 7216 14982 7268
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6512 7160 6653 7188
rect 6512 7148 6518 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 8110 7148 8116 7200
rect 8168 7148 8174 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 9732 7160 10701 7188
rect 9732 7148 9738 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 15102 7188 15108 7200
rect 13955 7160 15108 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 1104 7098 20884 7120
rect 1104 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 8367 7098
rect 8419 7046 8431 7098
rect 8483 7046 8495 7098
rect 8547 7046 8559 7098
rect 8611 7046 8623 7098
rect 8675 7046 13312 7098
rect 13364 7046 13376 7098
rect 13428 7046 13440 7098
rect 13492 7046 13504 7098
rect 13556 7046 13568 7098
rect 13620 7046 18257 7098
rect 18309 7046 18321 7098
rect 18373 7046 18385 7098
rect 18437 7046 18449 7098
rect 18501 7046 18513 7098
rect 18565 7046 20884 7098
rect 1104 7024 20884 7046
rect 4522 6944 4528 6996
rect 4580 6944 4586 6996
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 6365 6987 6423 6993
rect 6365 6984 6377 6987
rect 4847 6956 6377 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 6365 6953 6377 6956
rect 6411 6984 6423 6987
rect 6730 6984 6736 6996
rect 6411 6956 6736 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12308 6956 12449 6984
rect 12308 6944 12314 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14240 6956 14749 6984
rect 14240 6944 14246 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 14737 6947 14795 6953
rect 16850 6916 16856 6928
rect 12452 6888 12940 6916
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2866 6848 2872 6860
rect 2087 6820 2872 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4706 6848 4712 6860
rect 4356 6820 4712 6848
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 4356 6789 4384 6820
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6848 5963 6851
rect 7374 6848 7380 6860
rect 5951 6820 7380 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 10594 6808 10600 6860
rect 10652 6848 10658 6860
rect 12452 6848 12480 6888
rect 12802 6848 12808 6860
rect 10652 6820 12480 6848
rect 12544 6820 12808 6848
rect 10652 6808 10658 6820
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 2188 6752 2237 6780
rect 2188 6740 2194 6752
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4540 6712 4568 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5776 6752 6009 6780
rect 5776 6740 5782 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6454 6780 6460 6792
rect 6227 6752 6460 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6196 6712 6224 6743
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 10796 6789 10824 6820
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11238 6780 11244 6792
rect 10919 6752 11244 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11238 6740 11244 6752
rect 11296 6780 11302 6792
rect 12544 6780 12572 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12912 6848 12940 6888
rect 14936 6888 16856 6916
rect 12989 6851 13047 6857
rect 12989 6848 13001 6851
rect 12912 6820 13001 6848
rect 12989 6817 13001 6820
rect 13035 6848 13047 6851
rect 14936 6848 14964 6888
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 13035 6820 14964 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 17218 6848 17224 6860
rect 15068 6820 17224 6848
rect 15068 6808 15074 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 11296 6752 12572 6780
rect 12621 6783 12679 6789
rect 11296 6740 11302 6752
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 13722 6780 13728 6792
rect 12667 6752 13728 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 4540 6684 6224 6712
rect 10597 6715 10655 6721
rect 10597 6681 10609 6715
rect 10643 6712 10655 6715
rect 12636 6712 12664 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 15160 6752 15209 6780
rect 15160 6740 15166 6752
rect 15197 6749 15209 6752
rect 15243 6780 15255 6783
rect 16758 6780 16764 6792
rect 15243 6752 16764 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 16908 6752 16953 6780
rect 16908 6740 16914 6752
rect 10643 6684 12664 6712
rect 12713 6715 12771 6721
rect 10643 6681 10655 6684
rect 10597 6675 10655 6681
rect 12713 6681 12725 6715
rect 12759 6712 12771 6715
rect 12894 6712 12900 6724
rect 12759 6684 12900 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 17129 6715 17187 6721
rect 17129 6712 17141 6715
rect 13504 6684 17141 6712
rect 13504 6672 13510 6684
rect 17129 6681 17141 6684
rect 17175 6712 17187 6715
rect 17402 6712 17408 6724
rect 17175 6684 17408 6712
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2498 6644 2504 6656
rect 2455 6616 2504 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 10686 6604 10692 6656
rect 10744 6653 10750 6656
rect 10744 6607 10753 6653
rect 10744 6604 10750 6607
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 12912 6644 12940 6672
rect 15286 6644 15292 6656
rect 12912 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 21043 6576
rect 1104 6502 5894 6554
rect 5946 6502 5958 6554
rect 6010 6502 6022 6554
rect 6074 6502 6086 6554
rect 6138 6502 6150 6554
rect 6202 6502 10839 6554
rect 10891 6502 10903 6554
rect 10955 6502 10967 6554
rect 11019 6502 11031 6554
rect 11083 6502 11095 6554
rect 11147 6502 15784 6554
rect 15836 6502 15848 6554
rect 15900 6502 15912 6554
rect 15964 6502 15976 6554
rect 16028 6502 16040 6554
rect 16092 6502 20729 6554
rect 20781 6502 20793 6554
rect 20845 6502 20857 6554
rect 20909 6502 20921 6554
rect 20973 6502 20985 6554
rect 21037 6502 21043 6554
rect 1104 6480 21043 6502
rect 9582 6440 9588 6452
rect 8772 6412 9588 6440
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 1854 6264 1860 6316
rect 1912 6264 1918 6316
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 4338 6264 4344 6316
rect 4396 6264 4402 6316
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 6914 6304 6920 6316
rect 6871 6276 6920 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8110 6304 8116 6316
rect 7791 6276 8116 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6236 2927 6239
rect 4614 6236 4620 6248
rect 2915 6208 4620 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 5960 6208 6561 6236
rect 5960 6196 5966 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 7024 6236 7052 6267
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 6788 6208 7052 6236
rect 6788 6196 6794 6208
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7248 6208 7941 6236
rect 7248 6196 7254 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 8772 6236 8800 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 13446 6440 13452 6452
rect 11992 6412 13452 6440
rect 9490 6372 9496 6384
rect 8864 6344 9496 6372
rect 8864 6313 8892 6344
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9674 6304 9680 6316
rect 9355 6276 9680 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8772 6208 8953 6236
rect 7929 6199 7987 6205
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 5718 6128 5724 6180
rect 5776 6168 5782 6180
rect 9140 6168 9168 6267
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10284 6276 10333 6304
rect 10284 6264 10290 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10686 6304 10692 6316
rect 10643 6276 10692 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11238 6304 11244 6316
rect 10919 6276 11244 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11992 6313 12020 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13541 6443 13599 6449
rect 13541 6409 13553 6443
rect 13587 6440 13599 6443
rect 13630 6440 13636 6452
rect 13587 6412 13636 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 16850 6440 16856 6452
rect 14056 6412 16856 6440
rect 14056 6400 14062 6412
rect 16850 6400 16856 6412
rect 16908 6440 16914 6452
rect 17770 6440 17776 6452
rect 16908 6412 17776 6440
rect 16908 6400 16914 6412
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 13265 6375 13323 6381
rect 13265 6372 13277 6375
rect 12406 6344 13277 6372
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 12406 6304 12434 6344
rect 13265 6341 13277 6344
rect 13311 6372 13323 6375
rect 13722 6372 13728 6384
rect 13311 6344 13728 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 14274 6372 14280 6384
rect 13863 6344 14280 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 14274 6332 14280 6344
rect 14332 6372 14338 6384
rect 14458 6372 14464 6384
rect 14332 6344 14464 6372
rect 14332 6332 14338 6344
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 14550 6332 14556 6384
rect 14608 6372 14614 6384
rect 14608 6344 15700 6372
rect 14608 6332 14614 6344
rect 11977 6267 12035 6273
rect 12084 6276 12434 6304
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 12084 6236 12112 6276
rect 13078 6264 13084 6316
rect 13136 6304 13142 6316
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 13136 6276 13461 6304
rect 13136 6264 13142 6276
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 13998 6304 14004 6316
rect 13679 6276 14004 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 15672 6313 15700 6344
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 18138 6372 18144 6384
rect 16816 6344 18144 6372
rect 16816 6332 16822 6344
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 11204 6208 12112 6236
rect 11204 6196 11210 6208
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 14366 6196 14372 6248
rect 14424 6196 14430 6248
rect 14826 6236 14832 6248
rect 14752 6208 14832 6236
rect 14752 6177 14780 6208
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 5776 6140 9168 6168
rect 14737 6171 14795 6177
rect 5776 6128 5782 6140
rect 14737 6137 14749 6171
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 15473 6171 15531 6177
rect 15473 6137 15485 6171
rect 15519 6168 15531 6171
rect 15654 6168 15660 6180
rect 15519 6140 15660 6168
rect 15519 6137 15531 6140
rect 15473 6131 15531 6137
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 4706 6100 4712 6112
rect 4479 6072 4712 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 9122 6100 9128 6112
rect 8711 6072 9128 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 10652 6072 11805 6100
rect 10652 6060 10658 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 12710 6100 12716 6112
rect 12207 6072 12716 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15378 6100 15384 6112
rect 14875 6072 15384 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 16040 6100 16068 6199
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 17696 6245 17724 6344
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17681 6239 17739 6245
rect 17681 6205 17693 6239
rect 17727 6205 17739 6239
rect 17681 6199 17739 6205
rect 17604 6168 17632 6199
rect 17770 6196 17776 6248
rect 17828 6196 17834 6248
rect 17954 6168 17960 6180
rect 17604 6140 17960 6168
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 18046 6100 18052 6112
rect 16040 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 1104 6010 20884 6032
rect 1104 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 8367 6010
rect 8419 5958 8431 6010
rect 8483 5958 8495 6010
rect 8547 5958 8559 6010
rect 8611 5958 8623 6010
rect 8675 5958 13312 6010
rect 13364 5958 13376 6010
rect 13428 5958 13440 6010
rect 13492 5958 13504 6010
rect 13556 5958 13568 6010
rect 13620 5958 18257 6010
rect 18309 5958 18321 6010
rect 18373 5958 18385 6010
rect 18437 5958 18449 6010
rect 18501 5958 18513 6010
rect 18565 5958 20884 6010
rect 1104 5936 20884 5958
rect 2038 5856 2044 5908
rect 2096 5856 2102 5908
rect 5902 5856 5908 5908
rect 5960 5856 5966 5908
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 10505 5899 10563 5905
rect 10505 5896 10517 5899
rect 7156 5868 10517 5896
rect 7156 5856 7162 5868
rect 10505 5865 10517 5868
rect 10551 5865 10563 5899
rect 10505 5859 10563 5865
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 12618 5896 12624 5908
rect 12575 5868 12624 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 12759 5868 14289 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 14458 5856 14464 5908
rect 14516 5856 14522 5908
rect 5169 5831 5227 5837
rect 5169 5797 5181 5831
rect 5215 5828 5227 5831
rect 6822 5828 6828 5840
rect 5215 5800 6828 5828
rect 5215 5797 5227 5800
rect 5169 5791 5227 5797
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8938 5828 8944 5840
rect 8435 5800 8944 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 10594 5788 10600 5840
rect 10652 5788 10658 5840
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 13228 5800 13553 5828
rect 13228 5788 13234 5800
rect 13541 5797 13553 5800
rect 13587 5797 13599 5831
rect 13541 5791 13599 5797
rect 14366 5788 14372 5840
rect 14424 5828 14430 5840
rect 17129 5831 17187 5837
rect 14424 5800 16068 5828
rect 14424 5788 14430 5800
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2317 5763 2375 5769
rect 2317 5760 2329 5763
rect 2004 5732 2329 5760
rect 2004 5720 2010 5732
rect 2317 5729 2329 5732
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2240 5556 2268 5655
rect 2332 5624 2360 5723
rect 2498 5720 2504 5772
rect 2556 5720 2562 5772
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4709 5763 4767 5769
rect 4709 5760 4721 5763
rect 4580 5732 4721 5760
rect 4580 5720 4586 5732
rect 4709 5729 4721 5732
rect 4755 5729 4767 5763
rect 4709 5723 4767 5729
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5316 5732 6408 5760
rect 5316 5720 5322 5732
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 3234 5692 3240 5704
rect 2455 5664 3240 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 5810 5692 5816 5704
rect 4672 5664 5816 5692
rect 4672 5652 4678 5664
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6270 5692 6276 5704
rect 6043 5664 6276 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6380 5692 6408 5732
rect 6454 5720 6460 5772
rect 6512 5720 6518 5772
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 9582 5760 9588 5772
rect 8343 5732 9588 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 14568 5769 14596 5800
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10284 5732 10425 5760
rect 10284 5720 10290 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 15286 5720 15292 5772
rect 15344 5760 15350 5772
rect 16040 5769 16068 5800
rect 17129 5797 17141 5831
rect 17175 5828 17187 5831
rect 17678 5828 17684 5840
rect 17175 5800 17684 5828
rect 17175 5797 17187 5800
rect 17129 5791 17187 5797
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 15344 5732 15577 5760
rect 15344 5720 15350 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16025 5763 16083 5769
rect 16025 5729 16037 5763
rect 16071 5760 16083 5763
rect 16758 5760 16764 5772
rect 16071 5732 16764 5760
rect 16071 5729 16083 5732
rect 16025 5723 16083 5729
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 17954 5760 17960 5772
rect 17696 5732 17960 5760
rect 8205 5695 8263 5701
rect 6380 5664 8156 5692
rect 3050 5624 3056 5636
rect 2332 5596 3056 5624
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4338 5624 4344 5636
rect 3344 5596 4344 5624
rect 2958 5556 2964 5568
rect 2240 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5556 3022 5568
rect 3344 5556 3372 5596
rect 4338 5584 4344 5596
rect 4396 5584 4402 5636
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 5626 5624 5632 5636
rect 4764 5596 5632 5624
rect 4764 5584 4770 5596
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 6638 5584 6644 5636
rect 6696 5584 6702 5636
rect 7009 5627 7067 5633
rect 7009 5593 7021 5627
rect 7055 5624 7067 5627
rect 8021 5627 8079 5633
rect 8021 5624 8033 5627
rect 7055 5596 8033 5624
rect 7055 5593 7067 5596
rect 7009 5587 7067 5593
rect 8021 5593 8033 5596
rect 8067 5593 8079 5627
rect 8021 5587 8079 5593
rect 3016 5528 3372 5556
rect 3421 5559 3479 5565
rect 3016 5516 3022 5528
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 4246 5556 4252 5568
rect 3467 5528 4252 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 6730 5516 6736 5568
rect 6788 5516 6794 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 6914 5556 6920 5568
rect 6871 5528 6920 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 6914 5516 6920 5528
rect 6972 5556 6978 5568
rect 7650 5556 7656 5568
rect 6972 5528 7656 5556
rect 6972 5516 6978 5528
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8128 5556 8156 5664
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 9030 5692 9036 5704
rect 8527 5664 9036 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8220 5624 8248 5655
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 11146 5692 11152 5704
rect 10735 5664 11152 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12406 5664 13369 5692
rect 9490 5624 9496 5636
rect 8220 5596 9496 5624
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 12406 5556 12434 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 17696 5701 17724 5732
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 14936 5664 16129 5692
rect 12897 5627 12955 5633
rect 12897 5593 12909 5627
rect 12943 5624 12955 5627
rect 13170 5624 13176 5636
rect 12943 5596 13176 5624
rect 12943 5593 12955 5596
rect 12897 5587 12955 5593
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14936 5624 14964 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 17144 5624 17172 5655
rect 17862 5652 17868 5704
rect 17920 5652 17926 5704
rect 18046 5652 18052 5704
rect 18104 5692 18110 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 18104 5664 18245 5692
rect 18104 5652 18110 5664
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18138 5624 18144 5636
rect 14516 5596 14964 5624
rect 15764 5596 18144 5624
rect 14516 5584 14522 5596
rect 12710 5565 12716 5568
rect 8128 5528 12434 5556
rect 12697 5559 12716 5565
rect 12697 5525 12709 5559
rect 12697 5519 12716 5525
rect 12710 5516 12716 5519
rect 12768 5516 12774 5568
rect 15764 5565 15792 5596
rect 18138 5584 18144 5596
rect 18196 5584 18202 5636
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5525 15807 5559
rect 15749 5519 15807 5525
rect 1104 5466 21043 5488
rect 1104 5414 5894 5466
rect 5946 5414 5958 5466
rect 6010 5414 6022 5466
rect 6074 5414 6086 5466
rect 6138 5414 6150 5466
rect 6202 5414 10839 5466
rect 10891 5414 10903 5466
rect 10955 5414 10967 5466
rect 11019 5414 11031 5466
rect 11083 5414 11095 5466
rect 11147 5414 15784 5466
rect 15836 5414 15848 5466
rect 15900 5414 15912 5466
rect 15964 5414 15976 5466
rect 16028 5414 16040 5466
rect 16092 5414 20729 5466
rect 20781 5414 20793 5466
rect 20845 5414 20857 5466
rect 20909 5414 20921 5466
rect 20973 5414 20985 5466
rect 21037 5414 21043 5466
rect 1104 5392 21043 5414
rect 2133 5355 2191 5361
rect 2133 5321 2145 5355
rect 2179 5352 2191 5355
rect 2179 5324 4476 5352
rect 2179 5321 2191 5324
rect 2133 5315 2191 5321
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 4448 5284 4476 5324
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4580 5324 4813 5352
rect 4580 5312 4586 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6730 5352 6736 5364
rect 6043 5324 6736 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 6880 5324 8616 5352
rect 6880 5312 6886 5324
rect 5258 5284 5264 5296
rect 3292 5256 4200 5284
rect 4448 5256 5264 5284
rect 3292 5244 3298 5256
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1820 5188 2053 5216
rect 1820 5176 1826 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2056 5080 2084 5179
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 4172 5225 4200 5256
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5626 5244 5632 5296
rect 5684 5244 5690 5296
rect 5810 5244 5816 5296
rect 5868 5244 5874 5296
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 6328 5256 7512 5284
rect 6328 5244 6334 5256
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3108 5188 3985 5216
rect 3108 5176 3114 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4304 5188 4997 5216
rect 4304 5176 4310 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 7190 5216 7196 5228
rect 4985 5179 5043 5185
rect 6012 5188 7196 5216
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4430 5148 4436 5160
rect 4387 5120 4436 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4430 5108 4436 5120
rect 4488 5148 4494 5160
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4488 5120 5181 5148
rect 4488 5108 4494 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 6012 5080 6040 5188
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7484 5225 7512 5256
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 7576 5148 7604 5179
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8588 5225 8616 5324
rect 8680 5324 10885 5352
rect 8573 5219 8631 5225
rect 7708 5188 8432 5216
rect 7708 5176 7714 5188
rect 6144 5120 7604 5148
rect 6144 5108 6150 5120
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7984 5120 8309 5148
rect 7984 5108 7990 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8404 5148 8432 5188
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8680 5148 8708 5324
rect 10873 5321 10885 5324
rect 10919 5352 10931 5355
rect 17497 5355 17555 5361
rect 10919 5324 15148 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 12710 5284 12716 5296
rect 8996 5256 10364 5284
rect 8996 5244 9002 5256
rect 9122 5176 9128 5228
rect 9180 5176 9186 5228
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 10336 5225 10364 5256
rect 11900 5256 12716 5284
rect 11900 5225 11928 5256
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 13188 5256 14228 5284
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 9640 5188 10149 5216
rect 9640 5176 9646 5188
rect 10137 5185 10149 5188
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12250 5216 12256 5228
rect 12115 5188 12256 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 8404 5120 8708 5148
rect 8297 5111 8355 5117
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 10888 5148 10916 5179
rect 12250 5176 12256 5188
rect 12308 5216 12314 5228
rect 13188 5216 13216 5256
rect 14200 5228 14228 5256
rect 12308 5188 13216 5216
rect 13265 5219 13323 5225
rect 12308 5176 12314 5188
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 13630 5216 13636 5228
rect 13311 5188 13636 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13630 5176 13636 5188
rect 13688 5216 13694 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13688 5188 14105 5216
rect 13688 5176 13694 5188
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14093 5179 14151 5185
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14292 5188 15025 5216
rect 9548 5120 10916 5148
rect 9548 5108 9554 5120
rect 12158 5108 12164 5160
rect 12216 5148 12222 5160
rect 12345 5151 12403 5157
rect 12345 5148 12357 5151
rect 12216 5120 12357 5148
rect 12216 5108 12222 5120
rect 12345 5117 12357 5120
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12483 5120 13001 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 13354 5108 13360 5160
rect 13412 5108 13418 5160
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 13722 5148 13728 5160
rect 13495 5120 13728 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 2056 5052 6040 5080
rect 9214 5040 9220 5092
rect 9272 5040 9278 5092
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 14292 5080 14320 5188
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15120 5148 15148 5324
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 18785 5355 18843 5361
rect 18785 5352 18797 5355
rect 17543 5324 18797 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 18785 5321 18797 5324
rect 18831 5352 18843 5355
rect 19610 5352 19616 5364
rect 18831 5324 19616 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 16574 5244 16580 5296
rect 16632 5284 16638 5296
rect 17589 5287 17647 5293
rect 17589 5284 17601 5287
rect 16632 5256 17601 5284
rect 16632 5244 16638 5256
rect 17589 5253 17601 5256
rect 17635 5253 17647 5287
rect 17589 5247 17647 5253
rect 18138 5244 18144 5296
rect 18196 5244 18202 5296
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15436 5188 15485 5216
rect 15436 5176 15442 5188
rect 15473 5185 15485 5188
rect 15519 5216 15531 5219
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 15519 5188 17417 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 16853 5151 16911 5157
rect 15120 5120 15424 5148
rect 15396 5089 15424 5120
rect 16853 5117 16865 5151
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 12032 5052 14320 5080
rect 15381 5083 15439 5089
rect 12032 5040 12038 5052
rect 15381 5049 15393 5083
rect 15427 5080 15439 5083
rect 16114 5080 16120 5092
rect 15427 5052 16120 5080
rect 15427 5049 15439 5052
rect 15381 5043 15439 5049
rect 16114 5040 16120 5052
rect 16172 5040 16178 5092
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 8110 5012 8116 5024
rect 7791 4984 8116 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 14458 5012 14464 5024
rect 13412 4984 14464 5012
rect 13412 4972 13418 4984
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 16868 5012 16896 5111
rect 17034 5108 17040 5160
rect 17092 5108 17098 5160
rect 17420 5080 17448 5179
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18288 5219 18346 5225
rect 18288 5216 18300 5219
rect 18012 5188 18300 5216
rect 18012 5176 18018 5188
rect 18288 5185 18300 5188
rect 18334 5185 18346 5219
rect 18288 5179 18346 5185
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18104 5120 18521 5148
rect 18104 5108 18110 5120
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 17954 5080 17960 5092
rect 17420 5052 17960 5080
rect 17954 5040 17960 5052
rect 18012 5080 18018 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 18012 5052 18429 5080
rect 18012 5040 18018 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 17494 5012 17500 5024
rect 16868 4984 17500 5012
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 1104 4922 20884 4944
rect 1104 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 8367 4922
rect 8419 4870 8431 4922
rect 8483 4870 8495 4922
rect 8547 4870 8559 4922
rect 8611 4870 8623 4922
rect 8675 4870 13312 4922
rect 13364 4870 13376 4922
rect 13428 4870 13440 4922
rect 13492 4870 13504 4922
rect 13556 4870 13568 4922
rect 13620 4870 18257 4922
rect 18309 4870 18321 4922
rect 18373 4870 18385 4922
rect 18437 4870 18449 4922
rect 18501 4870 18513 4922
rect 18565 4870 20884 4922
rect 1104 4848 20884 4870
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6638 4808 6644 4820
rect 6227 4780 6644 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12768 4780 13277 4808
rect 12768 4768 12774 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 15194 4768 15200 4820
rect 15252 4768 15258 4820
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 14734 4740 14740 4752
rect 7340 4712 14740 4740
rect 7340 4700 7346 4712
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 4387 4644 6132 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 6104 4616 6132 4644
rect 7926 4632 7932 4684
rect 7984 4632 7990 4684
rect 8110 4632 8116 4684
rect 8168 4632 8174 4684
rect 9582 4672 9588 4684
rect 8312 4644 9588 4672
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 8312 4613 8340 4644
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 14642 4672 14648 4684
rect 13188 4644 14648 4672
rect 13188 4616 13216 4644
rect 14642 4632 14648 4644
rect 14700 4672 14706 4684
rect 17034 4672 17040 4684
rect 14700 4644 17040 4672
rect 14700 4632 14706 4644
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9490 4604 9496 4616
rect 8619 4576 9496 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 14458 4604 14464 4616
rect 13403 4576 14464 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15212 4613 15240 4644
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 16482 4604 16488 4616
rect 15427 4576 16488 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 15396 4536 15424 4567
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 13780 4508 15424 4536
rect 13780 4496 13786 4508
rect 1104 4378 21043 4400
rect 1104 4326 5894 4378
rect 5946 4326 5958 4378
rect 6010 4326 6022 4378
rect 6074 4326 6086 4378
rect 6138 4326 6150 4378
rect 6202 4326 10839 4378
rect 10891 4326 10903 4378
rect 10955 4326 10967 4378
rect 11019 4326 11031 4378
rect 11083 4326 11095 4378
rect 11147 4326 15784 4378
rect 15836 4326 15848 4378
rect 15900 4326 15912 4378
rect 15964 4326 15976 4378
rect 16028 4326 16040 4378
rect 16092 4326 20729 4378
rect 20781 4326 20793 4378
rect 20845 4326 20857 4378
rect 20909 4326 20921 4378
rect 20973 4326 20985 4378
rect 21037 4326 21043 4378
rect 1104 4304 21043 4326
rect 4436 4140 4488 4146
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 6270 4128 6276 4140
rect 5399 4100 6276 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 4436 4082 4488 4088
rect 1104 3834 20884 3856
rect 1104 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 8367 3834
rect 8419 3782 8431 3834
rect 8483 3782 8495 3834
rect 8547 3782 8559 3834
rect 8611 3782 8623 3834
rect 8675 3782 13312 3834
rect 13364 3782 13376 3834
rect 13428 3782 13440 3834
rect 13492 3782 13504 3834
rect 13556 3782 13568 3834
rect 13620 3782 18257 3834
rect 18309 3782 18321 3834
rect 18373 3782 18385 3834
rect 18437 3782 18449 3834
rect 18501 3782 18513 3834
rect 18565 3782 20884 3834
rect 1104 3760 20884 3782
rect 1104 3290 21043 3312
rect 1104 3238 5894 3290
rect 5946 3238 5958 3290
rect 6010 3238 6022 3290
rect 6074 3238 6086 3290
rect 6138 3238 6150 3290
rect 6202 3238 10839 3290
rect 10891 3238 10903 3290
rect 10955 3238 10967 3290
rect 11019 3238 11031 3290
rect 11083 3238 11095 3290
rect 11147 3238 15784 3290
rect 15836 3238 15848 3290
rect 15900 3238 15912 3290
rect 15964 3238 15976 3290
rect 16028 3238 16040 3290
rect 16092 3238 20729 3290
rect 20781 3238 20793 3290
rect 20845 3238 20857 3290
rect 20909 3238 20921 3290
rect 20973 3238 20985 3290
rect 21037 3238 21043 3290
rect 1104 3216 21043 3238
rect 1104 2746 20884 2768
rect 1104 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 8367 2746
rect 8419 2694 8431 2746
rect 8483 2694 8495 2746
rect 8547 2694 8559 2746
rect 8611 2694 8623 2746
rect 8675 2694 13312 2746
rect 13364 2694 13376 2746
rect 13428 2694 13440 2746
rect 13492 2694 13504 2746
rect 13556 2694 13568 2746
rect 13620 2694 18257 2746
rect 18309 2694 18321 2746
rect 18373 2694 18385 2746
rect 18437 2694 18449 2746
rect 18501 2694 18513 2746
rect 18565 2694 20884 2746
rect 1104 2672 20884 2694
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 7892 2604 15056 2632
rect 7892 2592 7898 2604
rect 6362 2496 6368 2508
rect 2148 2468 6368 2496
rect 2148 2437 2176 2468
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 8076 2468 9812 2496
rect 8076 2456 8082 2468
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 9674 2388 9680 2440
rect 9732 2388 9738 2440
rect 9784 2428 9812 2468
rect 15028 2437 15056 2604
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 9784 2400 12357 2428
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2397 15071 2431
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 15013 2391 15071 2397
rect 16546 2400 17693 2428
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1636 2332 1869 2360
rect 1636 2320 1642 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 4246 2320 4252 2372
rect 4304 2360 4310 2372
rect 4525 2363 4583 2369
rect 4525 2360 4537 2363
rect 4304 2332 4537 2360
rect 4304 2320 4310 2332
rect 4525 2329 4537 2332
rect 4571 2329 4583 2363
rect 4525 2323 4583 2329
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 7193 2363 7251 2369
rect 7193 2360 7205 2363
rect 6972 2332 7205 2360
rect 6972 2320 6978 2332
rect 7193 2329 7205 2332
rect 7239 2329 7251 2363
rect 7193 2323 7251 2329
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2329 10011 2363
rect 9953 2323 10011 2329
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9968 2292 9996 2323
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12492 2332 12633 2360
rect 12492 2320 12498 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 15289 2363 15347 2369
rect 15289 2360 15301 2363
rect 15252 2332 15301 2360
rect 15252 2320 15258 2332
rect 15289 2329 15301 2332
rect 15335 2329 15347 2363
rect 15289 2323 15347 2329
rect 9732 2264 9996 2292
rect 9732 2252 9738 2264
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 16546 2292 16574 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 19886 2388 19892 2440
rect 19944 2388 19950 2440
rect 17954 2320 17960 2372
rect 18012 2320 18018 2372
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 20254 2360 20260 2372
rect 20211 2332 20260 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 10376 2264 16574 2292
rect 10376 2252 10382 2264
rect 1104 2202 21043 2224
rect 1104 2150 5894 2202
rect 5946 2150 5958 2202
rect 6010 2150 6022 2202
rect 6074 2150 6086 2202
rect 6138 2150 6150 2202
rect 6202 2150 10839 2202
rect 10891 2150 10903 2202
rect 10955 2150 10967 2202
rect 11019 2150 11031 2202
rect 11083 2150 11095 2202
rect 11147 2150 15784 2202
rect 15836 2150 15848 2202
rect 15900 2150 15912 2202
rect 15964 2150 15976 2202
rect 16028 2150 16040 2202
rect 16092 2150 20729 2202
rect 20781 2150 20793 2202
rect 20845 2150 20857 2202
rect 20909 2150 20921 2202
rect 20973 2150 20985 2202
rect 21037 2150 21043 2202
rect 1104 2128 21043 2150
<< via1 >>
rect 8024 19660 8076 19712
rect 14648 19660 14700 19712
rect 15660 19660 15712 19712
rect 5894 19558 5946 19610
rect 5958 19558 6010 19610
rect 6022 19558 6074 19610
rect 6086 19558 6138 19610
rect 6150 19558 6202 19610
rect 10839 19558 10891 19610
rect 10903 19558 10955 19610
rect 10967 19558 11019 19610
rect 11031 19558 11083 19610
rect 11095 19558 11147 19610
rect 15784 19558 15836 19610
rect 15848 19558 15900 19610
rect 15912 19558 15964 19610
rect 15976 19558 16028 19610
rect 16040 19558 16092 19610
rect 20729 19558 20781 19610
rect 20793 19558 20845 19610
rect 20857 19558 20909 19610
rect 20921 19558 20973 19610
rect 20985 19558 21037 19610
rect 2780 19456 2832 19508
rect 13728 19456 13780 19508
rect 11244 19388 11296 19440
rect 4160 19320 4212 19372
rect 5264 19320 5316 19372
rect 11888 19320 11940 19372
rect 17132 19388 17184 19440
rect 17776 19431 17828 19440
rect 17776 19397 17803 19431
rect 17803 19397 17828 19431
rect 17776 19388 17828 19397
rect 17960 19431 18012 19440
rect 17960 19397 17969 19431
rect 17969 19397 18003 19431
rect 18003 19397 18012 19431
rect 17960 19388 18012 19397
rect 18236 19388 18288 19440
rect 8024 19295 8076 19304
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 14648 19363 14700 19372
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 15292 19252 15344 19304
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 18052 19116 18104 19168
rect 3422 19014 3474 19066
rect 3486 19014 3538 19066
rect 3550 19014 3602 19066
rect 3614 19014 3666 19066
rect 3678 19014 3730 19066
rect 8367 19014 8419 19066
rect 8431 19014 8483 19066
rect 8495 19014 8547 19066
rect 8559 19014 8611 19066
rect 8623 19014 8675 19066
rect 13312 19014 13364 19066
rect 13376 19014 13428 19066
rect 13440 19014 13492 19066
rect 13504 19014 13556 19066
rect 13568 19014 13620 19066
rect 18257 19014 18309 19066
rect 18321 19014 18373 19066
rect 18385 19014 18437 19066
rect 18449 19014 18501 19066
rect 18513 19014 18565 19066
rect 4160 18912 4212 18964
rect 14832 18955 14884 18964
rect 14832 18921 14841 18955
rect 14841 18921 14875 18955
rect 14875 18921 14884 18955
rect 14832 18912 14884 18921
rect 16120 18912 16172 18964
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 2412 18776 2464 18828
rect 4068 18708 4120 18760
rect 5264 18708 5316 18760
rect 14832 18776 14884 18828
rect 8024 18708 8076 18760
rect 9220 18708 9272 18760
rect 11888 18708 11940 18760
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 15476 18819 15528 18828
rect 15476 18785 15485 18819
rect 15485 18785 15519 18819
rect 15519 18785 15528 18819
rect 15476 18776 15528 18785
rect 17132 18776 17184 18828
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17776 18776 17828 18828
rect 3148 18683 3200 18692
rect 3148 18649 3157 18683
rect 3157 18649 3191 18683
rect 3191 18649 3200 18683
rect 3148 18640 3200 18649
rect 3792 18640 3844 18692
rect 2136 18615 2188 18624
rect 2136 18581 2145 18615
rect 2145 18581 2179 18615
rect 2179 18581 2188 18615
rect 2136 18572 2188 18581
rect 2228 18572 2280 18624
rect 7288 18640 7340 18692
rect 17040 18708 17092 18760
rect 13728 18640 13780 18692
rect 14924 18640 14976 18692
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 15016 18572 15068 18624
rect 15200 18615 15252 18624
rect 15200 18581 15209 18615
rect 15209 18581 15243 18615
rect 15243 18581 15252 18615
rect 15200 18572 15252 18581
rect 17960 18572 18012 18624
rect 19248 18572 19300 18624
rect 5894 18470 5946 18522
rect 5958 18470 6010 18522
rect 6022 18470 6074 18522
rect 6086 18470 6138 18522
rect 6150 18470 6202 18522
rect 10839 18470 10891 18522
rect 10903 18470 10955 18522
rect 10967 18470 11019 18522
rect 11031 18470 11083 18522
rect 11095 18470 11147 18522
rect 15784 18470 15836 18522
rect 15848 18470 15900 18522
rect 15912 18470 15964 18522
rect 15976 18470 16028 18522
rect 16040 18470 16092 18522
rect 20729 18470 20781 18522
rect 20793 18470 20845 18522
rect 20857 18470 20909 18522
rect 20921 18470 20973 18522
rect 20985 18470 21037 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 2136 18300 2188 18352
rect 7104 18343 7156 18352
rect 7104 18309 7113 18343
rect 7113 18309 7147 18343
rect 7147 18309 7156 18343
rect 7104 18300 7156 18309
rect 7288 18343 7340 18352
rect 7288 18309 7297 18343
rect 7297 18309 7331 18343
rect 7331 18309 7340 18343
rect 7288 18300 7340 18309
rect 2412 18275 2464 18284
rect 2412 18241 2421 18275
rect 2421 18241 2455 18275
rect 2455 18241 2464 18275
rect 2412 18232 2464 18241
rect 3884 18232 3936 18284
rect 3148 18164 3200 18216
rect 12256 18275 12308 18284
rect 12256 18241 12290 18275
rect 12290 18241 12308 18275
rect 12256 18232 12308 18241
rect 15384 18300 15436 18352
rect 15844 18411 15896 18420
rect 15844 18377 15853 18411
rect 15853 18377 15887 18411
rect 15887 18377 15896 18411
rect 15844 18368 15896 18377
rect 18052 18411 18104 18420
rect 18052 18377 18061 18411
rect 18061 18377 18095 18411
rect 18095 18377 18104 18411
rect 18052 18368 18104 18377
rect 16120 18300 16172 18352
rect 17040 18300 17092 18352
rect 5264 18164 5316 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 11888 18164 11940 18216
rect 13636 18164 13688 18216
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 16120 18164 16172 18216
rect 17592 18232 17644 18284
rect 16212 18096 16264 18148
rect 16948 18096 17000 18148
rect 14372 18028 14424 18080
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 15476 18071 15528 18080
rect 15476 18037 15485 18071
rect 15485 18037 15519 18071
rect 15519 18037 15528 18071
rect 15476 18028 15528 18037
rect 15568 18028 15620 18080
rect 3422 17926 3474 17978
rect 3486 17926 3538 17978
rect 3550 17926 3602 17978
rect 3614 17926 3666 17978
rect 3678 17926 3730 17978
rect 8367 17926 8419 17978
rect 8431 17926 8483 17978
rect 8495 17926 8547 17978
rect 8559 17926 8611 17978
rect 8623 17926 8675 17978
rect 13312 17926 13364 17978
rect 13376 17926 13428 17978
rect 13440 17926 13492 17978
rect 13504 17926 13556 17978
rect 13568 17926 13620 17978
rect 18257 17926 18309 17978
rect 18321 17926 18373 17978
rect 18385 17926 18437 17978
rect 18449 17926 18501 17978
rect 18513 17926 18565 17978
rect 3884 17824 3936 17876
rect 4068 17824 4120 17876
rect 10968 17867 11020 17876
rect 10968 17833 10977 17867
rect 10977 17833 11011 17867
rect 11011 17833 11020 17867
rect 10968 17824 11020 17833
rect 15568 17824 15620 17876
rect 17224 17824 17276 17876
rect 15752 17756 15804 17808
rect 2044 17620 2096 17672
rect 2780 17620 2832 17672
rect 5264 17620 5316 17672
rect 9220 17620 9272 17672
rect 2412 17552 2464 17604
rect 7932 17552 7984 17604
rect 14556 17620 14608 17672
rect 15476 17688 15528 17740
rect 15568 17688 15620 17740
rect 17132 17620 17184 17672
rect 4988 17484 5040 17536
rect 15476 17552 15528 17604
rect 17040 17552 17092 17604
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 5894 17382 5946 17434
rect 5958 17382 6010 17434
rect 6022 17382 6074 17434
rect 6086 17382 6138 17434
rect 6150 17382 6202 17434
rect 10839 17382 10891 17434
rect 10903 17382 10955 17434
rect 10967 17382 11019 17434
rect 11031 17382 11083 17434
rect 11095 17382 11147 17434
rect 15784 17382 15836 17434
rect 15848 17382 15900 17434
rect 15912 17382 15964 17434
rect 15976 17382 16028 17434
rect 16040 17382 16092 17434
rect 20729 17382 20781 17434
rect 20793 17382 20845 17434
rect 20857 17382 20909 17434
rect 20921 17382 20973 17434
rect 20985 17382 21037 17434
rect 2412 17323 2464 17332
rect 2412 17289 2421 17323
rect 2421 17289 2455 17323
rect 2455 17289 2464 17323
rect 2412 17280 2464 17289
rect 15200 17280 15252 17332
rect 2044 17212 2096 17264
rect 3976 17212 4028 17264
rect 8760 17212 8812 17264
rect 15292 17212 15344 17264
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 9220 17144 9272 17196
rect 9404 17187 9456 17196
rect 9404 17153 9438 17187
rect 9438 17153 9456 17187
rect 9404 17144 9456 17153
rect 11888 17144 11940 17196
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 15476 17144 15528 17196
rect 17500 17212 17552 17264
rect 16396 17144 16448 17196
rect 16580 17144 16632 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 16672 17076 16724 17128
rect 15200 17008 15252 17060
rect 12348 16940 12400 16992
rect 15016 16940 15068 16992
rect 16764 16940 16816 16992
rect 3422 16838 3474 16890
rect 3486 16838 3538 16890
rect 3550 16838 3602 16890
rect 3614 16838 3666 16890
rect 3678 16838 3730 16890
rect 8367 16838 8419 16890
rect 8431 16838 8483 16890
rect 8495 16838 8547 16890
rect 8559 16838 8611 16890
rect 8623 16838 8675 16890
rect 13312 16838 13364 16890
rect 13376 16838 13428 16890
rect 13440 16838 13492 16890
rect 13504 16838 13556 16890
rect 13568 16838 13620 16890
rect 18257 16838 18309 16890
rect 18321 16838 18373 16890
rect 18385 16838 18437 16890
rect 18449 16838 18501 16890
rect 18513 16838 18565 16890
rect 3056 16736 3108 16788
rect 9404 16736 9456 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 15200 16668 15252 16720
rect 16580 16668 16632 16720
rect 16764 16711 16816 16720
rect 16764 16677 16773 16711
rect 16773 16677 16807 16711
rect 16807 16677 16816 16711
rect 16764 16668 16816 16677
rect 1768 16532 1820 16584
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 5264 16532 5316 16584
rect 15016 16600 15068 16652
rect 11888 16532 11940 16584
rect 15568 16600 15620 16652
rect 1860 16507 1912 16516
rect 1860 16473 1869 16507
rect 1869 16473 1903 16507
rect 1903 16473 1912 16507
rect 1860 16464 1912 16473
rect 2228 16464 2280 16516
rect 2320 16464 2372 16516
rect 13176 16464 13228 16516
rect 1952 16439 2004 16448
rect 1952 16405 1967 16439
rect 1967 16405 2001 16439
rect 2001 16405 2004 16439
rect 1952 16396 2004 16405
rect 12716 16396 12768 16448
rect 16304 16600 16356 16652
rect 17500 16600 17552 16652
rect 19248 16600 19300 16652
rect 16120 16532 16172 16584
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 16672 16464 16724 16516
rect 17776 16507 17828 16516
rect 17776 16473 17785 16507
rect 17785 16473 17819 16507
rect 17819 16473 17828 16507
rect 17776 16464 17828 16473
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 19708 16396 19760 16448
rect 20076 16439 20128 16448
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 5894 16294 5946 16346
rect 5958 16294 6010 16346
rect 6022 16294 6074 16346
rect 6086 16294 6138 16346
rect 6150 16294 6202 16346
rect 10839 16294 10891 16346
rect 10903 16294 10955 16346
rect 10967 16294 11019 16346
rect 11031 16294 11083 16346
rect 11095 16294 11147 16346
rect 15784 16294 15836 16346
rect 15848 16294 15900 16346
rect 15912 16294 15964 16346
rect 15976 16294 16028 16346
rect 16040 16294 16092 16346
rect 20729 16294 20781 16346
rect 20793 16294 20845 16346
rect 20857 16294 20909 16346
rect 20921 16294 20973 16346
rect 20985 16294 21037 16346
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 16396 16192 16448 16244
rect 16580 16192 16632 16244
rect 17316 16192 17368 16244
rect 17592 16192 17644 16244
rect 19800 16192 19852 16244
rect 2044 16124 2096 16176
rect 2228 16124 2280 16176
rect 4988 16167 5040 16176
rect 4988 16133 5006 16167
rect 5006 16133 5040 16167
rect 4988 16124 5040 16133
rect 9588 16124 9640 16176
rect 12348 16124 12400 16176
rect 1952 16056 2004 16108
rect 2504 16056 2556 16108
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 13728 16056 13780 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 15660 16056 15712 16108
rect 16856 16056 16908 16108
rect 17408 16056 17460 16108
rect 18880 16056 18932 16108
rect 1768 15988 1820 16040
rect 2044 15988 2096 16040
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 11888 15988 11940 16040
rect 2136 15920 2188 15972
rect 17500 15988 17552 16040
rect 2320 15852 2372 15904
rect 6736 15852 6788 15904
rect 7932 15852 7984 15904
rect 14832 15920 14884 15972
rect 16304 15963 16356 15972
rect 16304 15929 16313 15963
rect 16313 15929 16347 15963
rect 16347 15929 16356 15963
rect 16304 15920 16356 15929
rect 16396 15920 16448 15972
rect 19892 15988 19944 16040
rect 14464 15852 14516 15904
rect 15384 15852 15436 15904
rect 3422 15750 3474 15802
rect 3486 15750 3538 15802
rect 3550 15750 3602 15802
rect 3614 15750 3666 15802
rect 3678 15750 3730 15802
rect 8367 15750 8419 15802
rect 8431 15750 8483 15802
rect 8495 15750 8547 15802
rect 8559 15750 8611 15802
rect 8623 15750 8675 15802
rect 13312 15750 13364 15802
rect 13376 15750 13428 15802
rect 13440 15750 13492 15802
rect 13504 15750 13556 15802
rect 13568 15750 13620 15802
rect 18257 15750 18309 15802
rect 18321 15750 18373 15802
rect 18385 15750 18437 15802
rect 18449 15750 18501 15802
rect 18513 15750 18565 15802
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 5264 15648 5316 15700
rect 6736 15648 6788 15700
rect 16856 15648 16908 15700
rect 17316 15691 17368 15700
rect 17316 15657 17325 15691
rect 17325 15657 17359 15691
rect 17359 15657 17368 15691
rect 17316 15648 17368 15657
rect 19708 15648 19760 15700
rect 16672 15580 16724 15632
rect 17776 15580 17828 15632
rect 14464 15512 14516 15564
rect 17316 15512 17368 15564
rect 19340 15512 19392 15564
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 5816 15444 5868 15496
rect 17408 15444 17460 15496
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 9956 15376 10008 15428
rect 17500 15419 17552 15428
rect 17500 15385 17509 15419
rect 17509 15385 17543 15419
rect 17543 15385 17552 15419
rect 17500 15376 17552 15385
rect 19524 15376 19576 15428
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 18144 15308 18196 15360
rect 19708 15351 19760 15360
rect 19708 15317 19717 15351
rect 19717 15317 19751 15351
rect 19751 15317 19760 15351
rect 19708 15308 19760 15317
rect 5894 15206 5946 15258
rect 5958 15206 6010 15258
rect 6022 15206 6074 15258
rect 6086 15206 6138 15258
rect 6150 15206 6202 15258
rect 10839 15206 10891 15258
rect 10903 15206 10955 15258
rect 10967 15206 11019 15258
rect 11031 15206 11083 15258
rect 11095 15206 11147 15258
rect 15784 15206 15836 15258
rect 15848 15206 15900 15258
rect 15912 15206 15964 15258
rect 15976 15206 16028 15258
rect 16040 15206 16092 15258
rect 20729 15206 20781 15258
rect 20793 15206 20845 15258
rect 20857 15206 20909 15258
rect 20921 15206 20973 15258
rect 20985 15206 21037 15258
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 14556 15104 14608 15156
rect 15660 15104 15712 15156
rect 7104 15036 7156 15088
rect 8760 15036 8812 15088
rect 19524 15104 19576 15156
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 1952 14943 2004 14952
rect 1952 14909 1961 14943
rect 1961 14909 1995 14943
rect 1995 14909 2004 14943
rect 1952 14900 2004 14909
rect 6736 14943 6788 14952
rect 6736 14909 6745 14943
rect 6745 14909 6779 14943
rect 6779 14909 6788 14943
rect 6736 14900 6788 14909
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 15016 14968 15068 15020
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 17960 15079 18012 15088
rect 17960 15045 17969 15079
rect 17969 15045 18003 15079
rect 18003 15045 18012 15079
rect 17960 15036 18012 15045
rect 19340 15079 19392 15088
rect 19340 15045 19349 15079
rect 19349 15045 19383 15079
rect 19383 15045 19392 15079
rect 19340 15036 19392 15045
rect 15200 14968 15252 14977
rect 15660 14900 15712 14952
rect 17684 15011 17736 15020
rect 17684 14977 17693 15011
rect 17693 14977 17727 15011
rect 17727 14977 17736 15011
rect 17684 14968 17736 14977
rect 19524 14968 19576 15020
rect 16396 14900 16448 14952
rect 14924 14832 14976 14884
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 6920 14764 6972 14816
rect 14004 14764 14056 14816
rect 14740 14807 14792 14816
rect 14740 14773 14749 14807
rect 14749 14773 14783 14807
rect 14783 14773 14792 14807
rect 14740 14764 14792 14773
rect 14832 14764 14884 14816
rect 18144 14832 18196 14884
rect 19708 14900 19760 14952
rect 17132 14764 17184 14816
rect 19156 14807 19208 14816
rect 19156 14773 19165 14807
rect 19165 14773 19199 14807
rect 19199 14773 19208 14807
rect 19156 14764 19208 14773
rect 19800 14807 19852 14816
rect 19800 14773 19809 14807
rect 19809 14773 19843 14807
rect 19843 14773 19852 14807
rect 19800 14764 19852 14773
rect 3422 14662 3474 14714
rect 3486 14662 3538 14714
rect 3550 14662 3602 14714
rect 3614 14662 3666 14714
rect 3678 14662 3730 14714
rect 8367 14662 8419 14714
rect 8431 14662 8483 14714
rect 8495 14662 8547 14714
rect 8559 14662 8611 14714
rect 8623 14662 8675 14714
rect 13312 14662 13364 14714
rect 13376 14662 13428 14714
rect 13440 14662 13492 14714
rect 13504 14662 13556 14714
rect 13568 14662 13620 14714
rect 18257 14662 18309 14714
rect 18321 14662 18373 14714
rect 18385 14662 18437 14714
rect 18449 14662 18501 14714
rect 18513 14662 18565 14714
rect 2228 14560 2280 14612
rect 5816 14560 5868 14612
rect 14832 14560 14884 14612
rect 15660 14560 15712 14612
rect 13084 14492 13136 14544
rect 10692 14424 10744 14476
rect 2044 14356 2096 14408
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 5540 14356 5592 14408
rect 6736 14356 6788 14408
rect 11888 14356 11940 14408
rect 14372 14424 14424 14476
rect 15476 14424 15528 14476
rect 15660 14424 15712 14476
rect 16948 14356 17000 14408
rect 4160 14288 4212 14340
rect 6920 14288 6972 14340
rect 12256 14288 12308 14340
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 18052 14560 18104 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 19800 14424 19852 14476
rect 19340 14356 19392 14408
rect 18144 14288 18196 14340
rect 14556 14220 14608 14272
rect 17132 14220 17184 14272
rect 17960 14220 18012 14272
rect 19340 14220 19392 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 19708 14220 19760 14272
rect 5894 14118 5946 14170
rect 5958 14118 6010 14170
rect 6022 14118 6074 14170
rect 6086 14118 6138 14170
rect 6150 14118 6202 14170
rect 10839 14118 10891 14170
rect 10903 14118 10955 14170
rect 10967 14118 11019 14170
rect 11031 14118 11083 14170
rect 11095 14118 11147 14170
rect 15784 14118 15836 14170
rect 15848 14118 15900 14170
rect 15912 14118 15964 14170
rect 15976 14118 16028 14170
rect 16040 14118 16092 14170
rect 20729 14118 20781 14170
rect 20793 14118 20845 14170
rect 20857 14118 20909 14170
rect 20921 14118 20973 14170
rect 20985 14118 21037 14170
rect 10692 14016 10744 14068
rect 13084 14016 13136 14068
rect 14832 14016 14884 14068
rect 19432 14016 19484 14068
rect 19524 14016 19576 14068
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 5724 13880 5776 13932
rect 12072 13923 12124 13932
rect 12072 13889 12106 13923
rect 12106 13889 12124 13923
rect 12072 13880 12124 13889
rect 3976 13812 4028 13864
rect 4068 13812 4120 13864
rect 5448 13812 5500 13864
rect 2688 13744 2740 13796
rect 3240 13676 3292 13728
rect 9312 13812 9364 13864
rect 10416 13812 10468 13864
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 17408 13948 17460 14000
rect 16948 13880 17000 13932
rect 13728 13812 13780 13864
rect 17224 13880 17276 13932
rect 18604 13880 18656 13932
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 19524 13744 19576 13796
rect 19892 13744 19944 13796
rect 7932 13676 7984 13728
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 3422 13574 3474 13626
rect 3486 13574 3538 13626
rect 3550 13574 3602 13626
rect 3614 13574 3666 13626
rect 3678 13574 3730 13626
rect 8367 13574 8419 13626
rect 8431 13574 8483 13626
rect 8495 13574 8547 13626
rect 8559 13574 8611 13626
rect 8623 13574 8675 13626
rect 13312 13574 13364 13626
rect 13376 13574 13428 13626
rect 13440 13574 13492 13626
rect 13504 13574 13556 13626
rect 13568 13574 13620 13626
rect 18257 13574 18309 13626
rect 18321 13574 18373 13626
rect 18385 13574 18437 13626
rect 18449 13574 18501 13626
rect 18513 13574 18565 13626
rect 3976 13515 4028 13524
rect 3976 13481 3985 13515
rect 3985 13481 4019 13515
rect 4019 13481 4028 13515
rect 3976 13472 4028 13481
rect 15292 13472 15344 13524
rect 4160 13404 4212 13456
rect 2044 13336 2096 13388
rect 3240 13336 3292 13388
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 16948 13336 17000 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 2688 13268 2740 13320
rect 5448 13268 5500 13320
rect 5724 13268 5776 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 14648 13268 14700 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 17040 13268 17092 13320
rect 17224 13268 17276 13320
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 19340 13268 19392 13320
rect 19432 13200 19484 13252
rect 2228 13132 2280 13184
rect 15016 13132 15068 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 17132 13132 17184 13184
rect 19524 13132 19576 13184
rect 5894 13030 5946 13082
rect 5958 13030 6010 13082
rect 6022 13030 6074 13082
rect 6086 13030 6138 13082
rect 6150 13030 6202 13082
rect 10839 13030 10891 13082
rect 10903 13030 10955 13082
rect 10967 13030 11019 13082
rect 11031 13030 11083 13082
rect 11095 13030 11147 13082
rect 15784 13030 15836 13082
rect 15848 13030 15900 13082
rect 15912 13030 15964 13082
rect 15976 13030 16028 13082
rect 16040 13030 16092 13082
rect 20729 13030 20781 13082
rect 20793 13030 20845 13082
rect 20857 13030 20909 13082
rect 20921 13030 20973 13082
rect 20985 13030 21037 13082
rect 2136 12928 2188 12980
rect 15292 12928 15344 12980
rect 1860 12903 1912 12912
rect 1860 12869 1869 12903
rect 1869 12869 1903 12903
rect 1903 12869 1912 12903
rect 1860 12860 1912 12869
rect 2044 12903 2096 12912
rect 2044 12869 2053 12903
rect 2053 12869 2087 12903
rect 2087 12869 2096 12903
rect 2044 12860 2096 12869
rect 6920 12860 6972 12912
rect 16764 12860 16816 12912
rect 2228 12792 2280 12844
rect 14648 12792 14700 12844
rect 16948 12792 17000 12844
rect 17408 12860 17460 12912
rect 17684 12928 17736 12980
rect 18604 12860 18656 12912
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 16120 12724 16172 12776
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17960 12835 18012 12844
rect 17224 12792 17276 12801
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 17960 12792 18012 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 8024 12588 8076 12640
rect 14096 12588 14148 12640
rect 15108 12588 15160 12640
rect 16948 12588 17000 12640
rect 19616 12724 19668 12776
rect 19432 12699 19484 12708
rect 19432 12665 19441 12699
rect 19441 12665 19475 12699
rect 19475 12665 19484 12699
rect 19432 12656 19484 12665
rect 19984 12588 20036 12640
rect 3422 12486 3474 12538
rect 3486 12486 3538 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 8367 12486 8419 12538
rect 8431 12486 8483 12538
rect 8495 12486 8547 12538
rect 8559 12486 8611 12538
rect 8623 12486 8675 12538
rect 13312 12486 13364 12538
rect 13376 12486 13428 12538
rect 13440 12486 13492 12538
rect 13504 12486 13556 12538
rect 13568 12486 13620 12538
rect 18257 12486 18309 12538
rect 18321 12486 18373 12538
rect 18385 12486 18437 12538
rect 18449 12486 18501 12538
rect 18513 12486 18565 12538
rect 14648 12384 14700 12436
rect 15200 12384 15252 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 2228 12316 2280 12368
rect 2320 12180 2372 12232
rect 3148 12316 3200 12368
rect 15108 12359 15160 12368
rect 15108 12325 15117 12359
rect 15117 12325 15151 12359
rect 15151 12325 15160 12359
rect 15108 12316 15160 12325
rect 5448 12248 5500 12300
rect 6552 12248 6604 12300
rect 2044 12112 2096 12164
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 9312 12180 9364 12232
rect 12348 12180 12400 12232
rect 17960 12248 18012 12300
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17408 12180 17460 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 10508 12112 10560 12164
rect 14556 12112 14608 12164
rect 14924 12112 14976 12164
rect 17868 12112 17920 12164
rect 17040 12044 17092 12096
rect 17500 12087 17552 12096
rect 17500 12053 17509 12087
rect 17509 12053 17543 12087
rect 17543 12053 17552 12087
rect 17500 12044 17552 12053
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 19708 12044 19760 12096
rect 5894 11942 5946 11994
rect 5958 11942 6010 11994
rect 6022 11942 6074 11994
rect 6086 11942 6138 11994
rect 6150 11942 6202 11994
rect 10839 11942 10891 11994
rect 10903 11942 10955 11994
rect 10967 11942 11019 11994
rect 11031 11942 11083 11994
rect 11095 11942 11147 11994
rect 15784 11942 15836 11994
rect 15848 11942 15900 11994
rect 15912 11942 15964 11994
rect 15976 11942 16028 11994
rect 16040 11942 16092 11994
rect 20729 11942 20781 11994
rect 20793 11942 20845 11994
rect 20857 11942 20909 11994
rect 20921 11942 20973 11994
rect 20985 11942 21037 11994
rect 4068 11840 4120 11892
rect 2688 11772 2740 11824
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 19524 11840 19576 11892
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 14280 11772 14332 11824
rect 2320 11704 2372 11756
rect 5448 11704 5500 11756
rect 6552 11704 6604 11756
rect 7196 11747 7248 11756
rect 7196 11713 7230 11747
rect 7230 11713 7248 11747
rect 7196 11704 7248 11713
rect 9312 11704 9364 11756
rect 12716 11704 12768 11756
rect 14648 11704 14700 11756
rect 16672 11704 16724 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 19340 11704 19392 11756
rect 2872 11636 2924 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 11796 11636 11848 11688
rect 17500 11636 17552 11688
rect 15384 11611 15436 11620
rect 15384 11577 15393 11611
rect 15393 11577 15427 11611
rect 15427 11577 15436 11611
rect 15384 11568 15436 11577
rect 15568 11568 15620 11620
rect 16856 11568 16908 11620
rect 9128 11500 9180 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 14648 11500 14700 11552
rect 17224 11500 17276 11552
rect 3422 11398 3474 11450
rect 3486 11398 3538 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 8367 11398 8419 11450
rect 8431 11398 8483 11450
rect 8495 11398 8547 11450
rect 8559 11398 8611 11450
rect 8623 11398 8675 11450
rect 13312 11398 13364 11450
rect 13376 11398 13428 11450
rect 13440 11398 13492 11450
rect 13504 11398 13556 11450
rect 13568 11398 13620 11450
rect 18257 11398 18309 11450
rect 18321 11398 18373 11450
rect 18385 11398 18437 11450
rect 18449 11398 18501 11450
rect 18513 11398 18565 11450
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 2136 11228 2188 11280
rect 10324 11228 10376 11280
rect 15016 11228 15068 11280
rect 17224 11160 17276 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 9220 11092 9272 11144
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 14004 11092 14056 11144
rect 6828 11024 6880 11076
rect 8944 11024 8996 11076
rect 12072 11067 12124 11076
rect 12072 11033 12106 11067
rect 12106 11033 12124 11067
rect 12072 11024 12124 11033
rect 15200 11024 15252 11076
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 17408 11092 17460 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 19340 11092 19392 11144
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 19616 11024 19668 11033
rect 19432 10999 19484 11008
rect 19432 10965 19441 10999
rect 19441 10965 19475 10999
rect 19475 10965 19484 10999
rect 19432 10956 19484 10965
rect 5894 10854 5946 10906
rect 5958 10854 6010 10906
rect 6022 10854 6074 10906
rect 6086 10854 6138 10906
rect 6150 10854 6202 10906
rect 10839 10854 10891 10906
rect 10903 10854 10955 10906
rect 10967 10854 11019 10906
rect 11031 10854 11083 10906
rect 11095 10854 11147 10906
rect 15784 10854 15836 10906
rect 15848 10854 15900 10906
rect 15912 10854 15964 10906
rect 15976 10854 16028 10906
rect 16040 10854 16092 10906
rect 20729 10854 20781 10906
rect 20793 10854 20845 10906
rect 20857 10854 20909 10906
rect 20921 10854 20973 10906
rect 20985 10854 21037 10906
rect 1860 10752 1912 10804
rect 1860 10616 1912 10668
rect 7012 10684 7064 10736
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 15200 10752 15252 10804
rect 15016 10684 15068 10736
rect 16764 10752 16816 10804
rect 17040 10684 17092 10736
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 4160 10548 4212 10600
rect 5264 10548 5316 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 15476 10616 15528 10668
rect 17776 10684 17828 10736
rect 18052 10727 18104 10736
rect 18052 10693 18079 10727
rect 18079 10693 18104 10727
rect 18052 10684 18104 10693
rect 19340 10795 19392 10804
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 18696 10684 18748 10736
rect 17316 10616 17368 10668
rect 17500 10616 17552 10668
rect 20076 10616 20128 10668
rect 15108 10548 15160 10600
rect 17776 10548 17828 10600
rect 19616 10548 19668 10600
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 14188 10412 14240 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 14556 10412 14608 10464
rect 15660 10412 15712 10464
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 18696 10412 18748 10464
rect 3422 10310 3474 10362
rect 3486 10310 3538 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 8367 10310 8419 10362
rect 8431 10310 8483 10362
rect 8495 10310 8547 10362
rect 8559 10310 8611 10362
rect 8623 10310 8675 10362
rect 13312 10310 13364 10362
rect 13376 10310 13428 10362
rect 13440 10310 13492 10362
rect 13504 10310 13556 10362
rect 13568 10310 13620 10362
rect 18257 10310 18309 10362
rect 18321 10310 18373 10362
rect 18385 10310 18437 10362
rect 18449 10310 18501 10362
rect 18513 10310 18565 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 14188 10208 14240 10260
rect 15200 10208 15252 10260
rect 17500 10208 17552 10260
rect 1952 10072 2004 10124
rect 9312 10072 9364 10124
rect 11796 10072 11848 10124
rect 15108 10072 15160 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2136 10004 2188 10056
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 10600 9936 10652 9988
rect 15200 9979 15252 9988
rect 15200 9945 15209 9979
rect 15209 9945 15243 9979
rect 15243 9945 15252 9979
rect 15200 9936 15252 9945
rect 17040 10004 17092 10056
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 19248 10140 19300 10192
rect 19616 10004 19668 10056
rect 19340 9936 19392 9988
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 15108 9868 15160 9920
rect 19800 9911 19852 9920
rect 19800 9877 19809 9911
rect 19809 9877 19843 9911
rect 19843 9877 19852 9911
rect 19800 9868 19852 9877
rect 5894 9766 5946 9818
rect 5958 9766 6010 9818
rect 6022 9766 6074 9818
rect 6086 9766 6138 9818
rect 6150 9766 6202 9818
rect 10839 9766 10891 9818
rect 10903 9766 10955 9818
rect 10967 9766 11019 9818
rect 11031 9766 11083 9818
rect 11095 9766 11147 9818
rect 15784 9766 15836 9818
rect 15848 9766 15900 9818
rect 15912 9766 15964 9818
rect 15976 9766 16028 9818
rect 16040 9766 16092 9818
rect 20729 9766 20781 9818
rect 20793 9766 20845 9818
rect 20857 9766 20909 9818
rect 20921 9766 20973 9818
rect 20985 9766 21037 9818
rect 3976 9460 4028 9512
rect 5264 9664 5316 9716
rect 6552 9664 6604 9716
rect 14740 9596 14792 9648
rect 19800 9664 19852 9716
rect 20076 9707 20128 9716
rect 20076 9673 20085 9707
rect 20085 9673 20119 9707
rect 20119 9673 20128 9707
rect 20076 9664 20128 9673
rect 4712 9528 4764 9580
rect 8852 9528 8904 9580
rect 9220 9528 9272 9580
rect 11796 9528 11848 9580
rect 12164 9571 12216 9580
rect 12164 9537 12198 9571
rect 12198 9537 12216 9571
rect 12164 9528 12216 9537
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 14464 9528 14516 9580
rect 17132 9596 17184 9648
rect 19156 9596 19208 9648
rect 8760 9460 8812 9512
rect 9312 9460 9364 9512
rect 14556 9460 14608 9512
rect 7472 9324 7524 9376
rect 15108 9435 15160 9444
rect 15108 9401 15117 9435
rect 15117 9401 15151 9435
rect 15151 9401 15160 9435
rect 15108 9392 15160 9401
rect 9772 9324 9824 9376
rect 10692 9324 10744 9376
rect 13820 9324 13872 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14464 9324 14516 9376
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 17500 9528 17552 9580
rect 16856 9460 16908 9512
rect 17684 9503 17736 9512
rect 17684 9469 17693 9503
rect 17693 9469 17727 9503
rect 17727 9469 17736 9503
rect 17684 9460 17736 9469
rect 19248 9460 19300 9512
rect 19616 9528 19668 9580
rect 17592 9392 17644 9444
rect 18052 9392 18104 9444
rect 3422 9222 3474 9274
rect 3486 9222 3538 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 8367 9222 8419 9274
rect 8431 9222 8483 9274
rect 8495 9222 8547 9274
rect 8559 9222 8611 9274
rect 8623 9222 8675 9274
rect 13312 9222 13364 9274
rect 13376 9222 13428 9274
rect 13440 9222 13492 9274
rect 13504 9222 13556 9274
rect 13568 9222 13620 9274
rect 18257 9222 18309 9274
rect 18321 9222 18373 9274
rect 18385 9222 18437 9274
rect 18449 9222 18501 9274
rect 18513 9222 18565 9274
rect 8944 9120 8996 9172
rect 14280 9120 14332 9172
rect 17040 9120 17092 9172
rect 17500 9120 17552 9172
rect 17684 9120 17736 9172
rect 10508 9052 10560 9104
rect 17592 9052 17644 9104
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 8760 8984 8812 9036
rect 14556 8984 14608 9036
rect 15016 8984 15068 9036
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 6736 8916 6788 8968
rect 8944 8916 8996 8968
rect 9496 8916 9548 8968
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 19248 8984 19300 9036
rect 4528 8848 4580 8900
rect 5724 8848 5776 8900
rect 14004 8848 14056 8900
rect 14648 8848 14700 8900
rect 1860 8780 1912 8832
rect 4804 8780 4856 8832
rect 6368 8780 6420 8832
rect 15016 8823 15068 8832
rect 15016 8789 15025 8823
rect 15025 8789 15059 8823
rect 15059 8789 15068 8823
rect 15016 8780 15068 8789
rect 15292 8848 15344 8900
rect 16580 8848 16632 8900
rect 17500 8916 17552 8968
rect 19156 8916 19208 8968
rect 17868 8780 17920 8832
rect 5894 8678 5946 8730
rect 5958 8678 6010 8730
rect 6022 8678 6074 8730
rect 6086 8678 6138 8730
rect 6150 8678 6202 8730
rect 10839 8678 10891 8730
rect 10903 8678 10955 8730
rect 10967 8678 11019 8730
rect 11031 8678 11083 8730
rect 11095 8678 11147 8730
rect 15784 8678 15836 8730
rect 15848 8678 15900 8730
rect 15912 8678 15964 8730
rect 15976 8678 16028 8730
rect 16040 8678 16092 8730
rect 20729 8678 20781 8730
rect 20793 8678 20845 8730
rect 20857 8678 20909 8730
rect 20921 8678 20973 8730
rect 20985 8678 21037 8730
rect 4160 8576 4212 8628
rect 4712 8576 4764 8628
rect 7196 8576 7248 8628
rect 12164 8576 12216 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17592 8576 17644 8628
rect 5540 8508 5592 8560
rect 9588 8508 9640 8560
rect 14464 8508 14516 8560
rect 1952 8440 2004 8492
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 4528 8440 4580 8492
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 5632 8440 5684 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 2044 8304 2096 8356
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 14924 8508 14976 8560
rect 16672 8508 16724 8560
rect 8760 8236 8812 8288
rect 10968 8236 11020 8288
rect 13728 8372 13780 8424
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 12808 8236 12860 8288
rect 14648 8440 14700 8492
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 16856 8440 16908 8492
rect 14740 8372 14792 8424
rect 17040 8372 17092 8424
rect 19248 8508 19300 8560
rect 19340 8508 19392 8560
rect 19800 8508 19852 8560
rect 17316 8440 17368 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 17592 8372 17644 8424
rect 17684 8372 17736 8424
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 19616 8372 19668 8424
rect 17132 8304 17184 8356
rect 17960 8236 18012 8288
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 8367 8134 8419 8186
rect 8431 8134 8483 8186
rect 8495 8134 8547 8186
rect 8559 8134 8611 8186
rect 8623 8134 8675 8186
rect 13312 8134 13364 8186
rect 13376 8134 13428 8186
rect 13440 8134 13492 8186
rect 13504 8134 13556 8186
rect 13568 8134 13620 8186
rect 18257 8134 18309 8186
rect 18321 8134 18373 8186
rect 18385 8134 18437 8186
rect 18449 8134 18501 8186
rect 18513 8134 18565 8186
rect 2320 8032 2372 8084
rect 5724 8032 5776 8084
rect 6920 8032 6972 8084
rect 8852 8032 8904 8084
rect 9036 8032 9088 8084
rect 10600 8032 10652 8084
rect 8484 7964 8536 8016
rect 10968 7964 11020 8016
rect 4620 7896 4672 7948
rect 10232 7896 10284 7948
rect 12348 7964 12400 8016
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 13176 8032 13228 8084
rect 14648 8075 14700 8084
rect 14648 8041 14657 8075
rect 14657 8041 14691 8075
rect 14691 8041 14700 8075
rect 14648 8032 14700 8041
rect 15384 8032 15436 8084
rect 16120 8032 16172 8084
rect 12808 7964 12860 8016
rect 17040 8032 17092 8084
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 19800 8075 19852 8084
rect 19800 8041 19809 8075
rect 19809 8041 19843 8075
rect 19843 8041 19852 8075
rect 19800 8032 19852 8041
rect 2044 7828 2096 7880
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 1768 7760 1820 7812
rect 4712 7828 4764 7880
rect 5540 7828 5592 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 6000 7828 6052 7880
rect 6460 7828 6512 7880
rect 6644 7828 6696 7880
rect 7380 7760 7432 7812
rect 8300 7828 8352 7880
rect 8944 7828 8996 7880
rect 9864 7828 9916 7880
rect 10600 7828 10652 7880
rect 11060 7828 11112 7880
rect 12624 7896 12676 7948
rect 12072 7828 12124 7880
rect 17592 7964 17644 8016
rect 13268 7896 13320 7948
rect 13636 7896 13688 7948
rect 9220 7760 9272 7812
rect 9680 7803 9732 7812
rect 9680 7769 9689 7803
rect 9689 7769 9723 7803
rect 9723 7769 9732 7803
rect 9680 7760 9732 7769
rect 12256 7803 12308 7812
rect 12256 7769 12265 7803
rect 12265 7769 12299 7803
rect 12299 7769 12308 7803
rect 12256 7760 12308 7769
rect 12440 7803 12492 7812
rect 12440 7769 12481 7803
rect 12481 7769 12492 7803
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13544 7828 13596 7880
rect 15660 7896 15712 7948
rect 15292 7828 15344 7880
rect 12440 7760 12492 7769
rect 13728 7760 13780 7812
rect 16488 7896 16540 7948
rect 18144 7896 18196 7948
rect 17960 7828 18012 7880
rect 18880 7828 18932 7880
rect 17316 7803 17368 7812
rect 17316 7769 17343 7803
rect 17343 7769 17368 7803
rect 17316 7760 17368 7769
rect 17592 7760 17644 7812
rect 19616 7803 19668 7812
rect 19616 7769 19625 7803
rect 19625 7769 19659 7803
rect 19659 7769 19668 7803
rect 19616 7760 19668 7769
rect 1952 7692 2004 7744
rect 2136 7692 2188 7744
rect 3148 7692 3200 7744
rect 4712 7692 4764 7744
rect 6644 7692 6696 7744
rect 10140 7692 10192 7744
rect 12624 7692 12676 7744
rect 17684 7692 17736 7744
rect 5894 7590 5946 7642
rect 5958 7590 6010 7642
rect 6022 7590 6074 7642
rect 6086 7590 6138 7642
rect 6150 7590 6202 7642
rect 10839 7590 10891 7642
rect 10903 7590 10955 7642
rect 10967 7590 11019 7642
rect 11031 7590 11083 7642
rect 11095 7590 11147 7642
rect 15784 7590 15836 7642
rect 15848 7590 15900 7642
rect 15912 7590 15964 7642
rect 15976 7590 16028 7642
rect 16040 7590 16092 7642
rect 20729 7590 20781 7642
rect 20793 7590 20845 7642
rect 20857 7590 20909 7642
rect 20921 7590 20973 7642
rect 20985 7590 21037 7642
rect 2780 7488 2832 7540
rect 2964 7420 3016 7472
rect 5632 7488 5684 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 8300 7488 8352 7540
rect 10600 7488 10652 7540
rect 12256 7488 12308 7540
rect 13176 7488 13228 7540
rect 13728 7488 13780 7540
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 5264 7352 5316 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 6460 7352 6512 7404
rect 6092 7284 6144 7336
rect 6644 7352 6696 7404
rect 7196 7352 7248 7404
rect 7380 7352 7432 7404
rect 9496 7420 9548 7472
rect 9680 7420 9732 7472
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8760 7352 8812 7404
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10692 7352 10744 7404
rect 12348 7463 12400 7472
rect 12348 7429 12357 7463
rect 12357 7429 12391 7463
rect 12391 7429 12400 7463
rect 12348 7420 12400 7429
rect 15384 7488 15436 7540
rect 17776 7488 17828 7540
rect 19340 7488 19392 7540
rect 13544 7395 13596 7404
rect 6736 7284 6788 7336
rect 9036 7284 9088 7336
rect 12256 7284 12308 7336
rect 12440 7284 12492 7336
rect 12808 7284 12860 7336
rect 13544 7361 13550 7395
rect 13550 7361 13584 7395
rect 13584 7361 13596 7395
rect 13544 7352 13596 7361
rect 15200 7420 15252 7472
rect 16488 7420 16540 7472
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15292 7352 15344 7404
rect 16120 7352 16172 7404
rect 13820 7284 13872 7336
rect 15016 7284 15068 7336
rect 9588 7216 9640 7268
rect 9864 7259 9916 7268
rect 9864 7225 9873 7259
rect 9873 7225 9907 7259
rect 9907 7225 9916 7259
rect 9864 7216 9916 7225
rect 12532 7216 12584 7268
rect 14924 7259 14976 7268
rect 14924 7225 14933 7259
rect 14933 7225 14967 7259
rect 14967 7225 14976 7259
rect 14924 7216 14976 7225
rect 6460 7148 6512 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 9680 7148 9732 7200
rect 15108 7148 15160 7200
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 8367 7046 8419 7098
rect 8431 7046 8483 7098
rect 8495 7046 8547 7098
rect 8559 7046 8611 7098
rect 8623 7046 8675 7098
rect 13312 7046 13364 7098
rect 13376 7046 13428 7098
rect 13440 7046 13492 7098
rect 13504 7046 13556 7098
rect 13568 7046 13620 7098
rect 18257 7046 18309 7098
rect 18321 7046 18373 7098
rect 18385 7046 18437 7098
rect 18449 7046 18501 7098
rect 18513 7046 18565 7098
rect 4528 6987 4580 6996
rect 4528 6953 4537 6987
rect 4537 6953 4571 6987
rect 4571 6953 4580 6987
rect 4528 6944 4580 6953
rect 6736 6944 6788 6996
rect 12256 6944 12308 6996
rect 14188 6944 14240 6996
rect 2872 6808 2924 6860
rect 2136 6740 2188 6792
rect 4712 6808 4764 6860
rect 7380 6808 7432 6860
rect 10600 6808 10652 6860
rect 5724 6740 5776 6792
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6460 6740 6512 6792
rect 11244 6740 11296 6792
rect 12808 6808 12860 6860
rect 16856 6876 16908 6928
rect 15016 6808 15068 6860
rect 17224 6808 17276 6860
rect 13728 6740 13780 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 15108 6740 15160 6792
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 16856 6783 16908 6792
rect 16856 6749 16866 6783
rect 16866 6749 16900 6783
rect 16900 6749 16908 6783
rect 16856 6740 16908 6749
rect 12900 6672 12952 6724
rect 13452 6672 13504 6724
rect 17408 6672 17460 6724
rect 2504 6604 2556 6656
rect 10692 6647 10744 6656
rect 10692 6613 10707 6647
rect 10707 6613 10741 6647
rect 10741 6613 10744 6647
rect 10692 6604 10744 6613
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 15292 6604 15344 6656
rect 5894 6502 5946 6554
rect 5958 6502 6010 6554
rect 6022 6502 6074 6554
rect 6086 6502 6138 6554
rect 6150 6502 6202 6554
rect 10839 6502 10891 6554
rect 10903 6502 10955 6554
rect 10967 6502 11019 6554
rect 11031 6502 11083 6554
rect 11095 6502 11147 6554
rect 15784 6502 15836 6554
rect 15848 6502 15900 6554
rect 15912 6502 15964 6554
rect 15976 6502 16028 6554
rect 16040 6502 16092 6554
rect 20729 6502 20781 6554
rect 20793 6502 20845 6554
rect 20857 6502 20909 6554
rect 20921 6502 20973 6554
rect 20985 6502 21037 6554
rect 7380 6375 7432 6384
rect 7380 6341 7389 6375
rect 7389 6341 7423 6375
rect 7423 6341 7432 6375
rect 7380 6332 7432 6341
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 6920 6264 6972 6316
rect 4620 6196 4672 6248
rect 5908 6196 5960 6248
rect 6736 6196 6788 6248
rect 8116 6264 8168 6316
rect 7196 6196 7248 6248
rect 9588 6400 9640 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 9496 6332 9548 6384
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 5724 6128 5776 6180
rect 9680 6264 9732 6316
rect 10232 6264 10284 6316
rect 10692 6264 10744 6316
rect 11244 6264 11296 6316
rect 13452 6400 13504 6452
rect 13636 6400 13688 6452
rect 14004 6400 14056 6452
rect 16856 6400 16908 6452
rect 17776 6400 17828 6452
rect 13728 6332 13780 6384
rect 14280 6332 14332 6384
rect 14464 6332 14516 6384
rect 14556 6332 14608 6384
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 13084 6264 13136 6316
rect 14004 6264 14056 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 16764 6332 16816 6384
rect 11152 6196 11204 6205
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14832 6196 14884 6248
rect 15660 6128 15712 6180
rect 4712 6060 4764 6112
rect 9128 6060 9180 6112
rect 10600 6060 10652 6112
rect 12716 6060 12768 6112
rect 15384 6060 15436 6112
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 18144 6332 18196 6384
rect 17776 6239 17828 6248
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 17960 6128 18012 6180
rect 18052 6060 18104 6112
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 8367 5958 8419 6010
rect 8431 5958 8483 6010
rect 8495 5958 8547 6010
rect 8559 5958 8611 6010
rect 8623 5958 8675 6010
rect 13312 5958 13364 6010
rect 13376 5958 13428 6010
rect 13440 5958 13492 6010
rect 13504 5958 13556 6010
rect 13568 5958 13620 6010
rect 18257 5958 18309 6010
rect 18321 5958 18373 6010
rect 18385 5958 18437 6010
rect 18449 5958 18501 6010
rect 18513 5958 18565 6010
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 7104 5856 7156 5908
rect 12624 5856 12676 5908
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 6828 5788 6880 5840
rect 8944 5788 8996 5840
rect 10600 5831 10652 5840
rect 10600 5797 10609 5831
rect 10609 5797 10643 5831
rect 10643 5797 10652 5831
rect 10600 5788 10652 5797
rect 13176 5788 13228 5840
rect 14372 5788 14424 5840
rect 1952 5720 2004 5772
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 4528 5720 4580 5772
rect 5264 5720 5316 5772
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 5816 5695 5868 5704
rect 4620 5652 4672 5661
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6276 5652 6328 5704
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 9588 5720 9640 5772
rect 10232 5720 10284 5772
rect 15292 5720 15344 5772
rect 17684 5788 17736 5840
rect 16764 5720 16816 5772
rect 3056 5627 3108 5636
rect 3056 5593 3065 5627
rect 3065 5593 3099 5627
rect 3099 5593 3108 5627
rect 3056 5584 3108 5593
rect 2964 5516 3016 5568
rect 4344 5584 4396 5636
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 5632 5584 5684 5636
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 4252 5516 4304 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 6920 5516 6972 5568
rect 7656 5516 7708 5568
rect 9036 5652 9088 5704
rect 11152 5652 11204 5704
rect 9496 5584 9548 5636
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 17960 5720 18012 5772
rect 13176 5584 13228 5636
rect 14464 5584 14516 5636
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18052 5652 18104 5704
rect 12716 5559 12768 5568
rect 12716 5525 12743 5559
rect 12743 5525 12768 5559
rect 12716 5516 12768 5525
rect 18144 5584 18196 5636
rect 5894 5414 5946 5466
rect 5958 5414 6010 5466
rect 6022 5414 6074 5466
rect 6086 5414 6138 5466
rect 6150 5414 6202 5466
rect 10839 5414 10891 5466
rect 10903 5414 10955 5466
rect 10967 5414 11019 5466
rect 11031 5414 11083 5466
rect 11095 5414 11147 5466
rect 15784 5414 15836 5466
rect 15848 5414 15900 5466
rect 15912 5414 15964 5466
rect 15976 5414 16028 5466
rect 16040 5414 16092 5466
rect 20729 5414 20781 5466
rect 20793 5414 20845 5466
rect 20857 5414 20909 5466
rect 20921 5414 20973 5466
rect 20985 5414 21037 5466
rect 3240 5244 3292 5296
rect 4528 5312 4580 5364
rect 6736 5312 6788 5364
rect 6828 5312 6880 5364
rect 1768 5176 1820 5228
rect 3056 5176 3108 5228
rect 5264 5244 5316 5296
rect 5632 5287 5684 5296
rect 5632 5253 5641 5287
rect 5641 5253 5675 5287
rect 5675 5253 5684 5287
rect 5632 5244 5684 5253
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 6276 5244 6328 5296
rect 4252 5176 4304 5228
rect 7196 5219 7248 5228
rect 4436 5108 4488 5160
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 6092 5108 6144 5160
rect 7656 5176 7708 5228
rect 7932 5108 7984 5160
rect 8944 5244 8996 5296
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9588 5176 9640 5228
rect 12716 5244 12768 5296
rect 9496 5108 9548 5160
rect 12256 5176 12308 5228
rect 13636 5176 13688 5228
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 12164 5108 12216 5160
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 13728 5108 13780 5160
rect 9220 5083 9272 5092
rect 9220 5049 9229 5083
rect 9229 5049 9263 5083
rect 9263 5049 9272 5083
rect 9220 5040 9272 5049
rect 11980 5040 12032 5092
rect 19616 5312 19668 5364
rect 16580 5244 16632 5296
rect 18144 5287 18196 5296
rect 18144 5253 18153 5287
rect 18153 5253 18187 5287
rect 18187 5253 18196 5287
rect 18144 5244 18196 5253
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 15384 5176 15436 5228
rect 16120 5040 16172 5092
rect 8116 4972 8168 5024
rect 13360 4972 13412 5024
rect 14464 4972 14516 5024
rect 17040 5151 17092 5160
rect 17040 5117 17049 5151
rect 17049 5117 17083 5151
rect 17083 5117 17092 5151
rect 17040 5108 17092 5117
rect 17960 5176 18012 5228
rect 18052 5108 18104 5160
rect 17960 5040 18012 5092
rect 17500 4972 17552 5024
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 8367 4870 8419 4922
rect 8431 4870 8483 4922
rect 8495 4870 8547 4922
rect 8559 4870 8611 4922
rect 8623 4870 8675 4922
rect 13312 4870 13364 4922
rect 13376 4870 13428 4922
rect 13440 4870 13492 4922
rect 13504 4870 13556 4922
rect 13568 4870 13620 4922
rect 18257 4870 18309 4922
rect 18321 4870 18373 4922
rect 18385 4870 18437 4922
rect 18449 4870 18501 4922
rect 18513 4870 18565 4922
rect 6644 4768 6696 4820
rect 12716 4768 12768 4820
rect 15200 4811 15252 4820
rect 15200 4777 15209 4811
rect 15209 4777 15243 4811
rect 15243 4777 15252 4811
rect 15200 4768 15252 4777
rect 7288 4700 7340 4752
rect 14740 4700 14792 4752
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 8116 4675 8168 4684
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8116 4632 8168 4641
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 9588 4632 9640 4684
rect 14648 4632 14700 4684
rect 9496 4564 9548 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 14464 4564 14516 4616
rect 17040 4632 17092 4684
rect 13728 4496 13780 4548
rect 16488 4564 16540 4616
rect 5894 4326 5946 4378
rect 5958 4326 6010 4378
rect 6022 4326 6074 4378
rect 6086 4326 6138 4378
rect 6150 4326 6202 4378
rect 10839 4326 10891 4378
rect 10903 4326 10955 4378
rect 10967 4326 11019 4378
rect 11031 4326 11083 4378
rect 11095 4326 11147 4378
rect 15784 4326 15836 4378
rect 15848 4326 15900 4378
rect 15912 4326 15964 4378
rect 15976 4326 16028 4378
rect 16040 4326 16092 4378
rect 20729 4326 20781 4378
rect 20793 4326 20845 4378
rect 20857 4326 20909 4378
rect 20921 4326 20973 4378
rect 20985 4326 21037 4378
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4436 4088 4488 4140
rect 6276 4088 6328 4140
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 8367 3782 8419 3834
rect 8431 3782 8483 3834
rect 8495 3782 8547 3834
rect 8559 3782 8611 3834
rect 8623 3782 8675 3834
rect 13312 3782 13364 3834
rect 13376 3782 13428 3834
rect 13440 3782 13492 3834
rect 13504 3782 13556 3834
rect 13568 3782 13620 3834
rect 18257 3782 18309 3834
rect 18321 3782 18373 3834
rect 18385 3782 18437 3834
rect 18449 3782 18501 3834
rect 18513 3782 18565 3834
rect 5894 3238 5946 3290
rect 5958 3238 6010 3290
rect 6022 3238 6074 3290
rect 6086 3238 6138 3290
rect 6150 3238 6202 3290
rect 10839 3238 10891 3290
rect 10903 3238 10955 3290
rect 10967 3238 11019 3290
rect 11031 3238 11083 3290
rect 11095 3238 11147 3290
rect 15784 3238 15836 3290
rect 15848 3238 15900 3290
rect 15912 3238 15964 3290
rect 15976 3238 16028 3290
rect 16040 3238 16092 3290
rect 20729 3238 20781 3290
rect 20793 3238 20845 3290
rect 20857 3238 20909 3290
rect 20921 3238 20973 3290
rect 20985 3238 21037 3290
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 8367 2694 8419 2746
rect 8431 2694 8483 2746
rect 8495 2694 8547 2746
rect 8559 2694 8611 2746
rect 8623 2694 8675 2746
rect 13312 2694 13364 2746
rect 13376 2694 13428 2746
rect 13440 2694 13492 2746
rect 13504 2694 13556 2746
rect 13568 2694 13620 2746
rect 18257 2694 18309 2746
rect 18321 2694 18373 2746
rect 18385 2694 18437 2746
rect 18449 2694 18501 2746
rect 18513 2694 18565 2746
rect 7840 2592 7892 2644
rect 6368 2456 6420 2508
rect 8024 2456 8076 2508
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 1584 2320 1636 2372
rect 4252 2320 4304 2372
rect 6920 2320 6972 2372
rect 9680 2252 9732 2304
rect 12440 2320 12492 2372
rect 15200 2320 15252 2372
rect 10324 2252 10376 2304
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 17960 2363 18012 2372
rect 17960 2329 17969 2363
rect 17969 2329 18003 2363
rect 18003 2329 18012 2363
rect 17960 2320 18012 2329
rect 20260 2320 20312 2372
rect 5894 2150 5946 2202
rect 5958 2150 6010 2202
rect 6022 2150 6074 2202
rect 6086 2150 6138 2202
rect 6150 2150 6202 2202
rect 10839 2150 10891 2202
rect 10903 2150 10955 2202
rect 10967 2150 11019 2202
rect 11031 2150 11083 2202
rect 11095 2150 11147 2202
rect 15784 2150 15836 2202
rect 15848 2150 15900 2202
rect 15912 2150 15964 2202
rect 15976 2150 16028 2202
rect 16040 2150 16092 2202
rect 20729 2150 20781 2202
rect 20793 2150 20845 2202
rect 20857 2150 20909 2202
rect 20921 2150 20973 2202
rect 20985 2150 21037 2202
<< metal2 >>
rect 3698 21298 3754 22000
rect 10966 21298 11022 22000
rect 3698 21270 4016 21298
rect 3698 21200 3754 21270
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2148 18358 2176 18566
rect 2240 18426 2268 18566
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 2424 18290 2452 18770
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 17898 2452 18226
rect 2240 17870 2452 17898
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2056 17270 2084 17614
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 2056 17134 2084 17206
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1780 16046 1808 16526
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1872 14346 1900 16458
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16114 1992 16390
rect 2056 16182 2084 17070
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2044 16040 2096 16046
rect 1964 15988 2044 15994
rect 1964 15982 2096 15988
rect 1964 15966 2084 15982
rect 2148 15978 2176 16526
rect 2240 16522 2268 17870
rect 2792 17678 2820 19450
rect 3422 19068 3730 19077
rect 3422 19066 3428 19068
rect 3484 19066 3508 19068
rect 3564 19066 3588 19068
rect 3644 19066 3668 19068
rect 3724 19066 3730 19068
rect 3484 19014 3486 19066
rect 3666 19014 3668 19066
rect 3422 19012 3428 19014
rect 3484 19012 3508 19014
rect 3564 19012 3588 19014
rect 3644 19012 3668 19014
rect 3724 19012 3730 19014
rect 3422 19003 3730 19012
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 3160 18222 3188 18634
rect 3804 18426 3832 18634
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2424 17338 2452 17546
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3068 16794 3096 17138
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 16250 2360 16458
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2136 15972 2188 15978
rect 1964 14958 1992 15966
rect 2136 15914 2188 15920
rect 2240 15858 2268 16118
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2148 15830 2268 15858
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2148 15502 2176 15830
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1872 12918 1900 14282
rect 1964 14226 1992 14894
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2056 14414 2084 14758
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2044 14272 2096 14278
rect 1964 14220 2044 14226
rect 1964 14214 2096 14220
rect 1964 14198 2084 14214
rect 2056 13394 2084 14198
rect 2148 13870 2176 15438
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2240 14618 2268 14962
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12918 2084 13330
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 12986 2176 13262
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 2240 12850 2268 13126
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2056 11234 2084 12106
rect 1964 11206 2084 11234
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1872 10810 1900 11086
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 10062 1900 10610
rect 1964 10606 1992 11206
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10130 1992 10542
rect 2056 10266 2084 11086
rect 2148 10674 2176 11222
rect 2240 10674 2268 12310
rect 2332 12238 2360 15846
rect 2516 15706 2544 16050
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2700 13326 2728 13738
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2320 12232 2372 12238
rect 2372 12180 2452 12186
rect 2320 12174 2452 12180
rect 2332 12158 2452 12174
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11762 2360 12038
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 8922 1900 9998
rect 1964 9058 1992 10066
rect 2148 10062 2176 10610
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1964 9030 2084 9058
rect 2148 9042 2176 9998
rect 1872 8894 1992 8922
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 5234 1808 7754
rect 1872 6322 1900 8774
rect 1964 8498 1992 8894
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 7750 1992 8434
rect 2056 8362 2084 9030
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2056 7886 2084 8298
rect 2240 7886 2268 10610
rect 2424 8974 2452 12158
rect 2700 11830 2728 13262
rect 3160 12374 3188 18158
rect 3422 17980 3730 17989
rect 3422 17978 3428 17980
rect 3484 17978 3508 17980
rect 3564 17978 3588 17980
rect 3644 17978 3668 17980
rect 3724 17978 3730 17980
rect 3484 17926 3486 17978
rect 3666 17926 3668 17978
rect 3422 17924 3428 17926
rect 3484 17924 3508 17926
rect 3564 17924 3588 17926
rect 3644 17924 3668 17926
rect 3724 17924 3730 17926
rect 3422 17915 3730 17924
rect 3896 17882 3924 18226
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17270 4016 21270
rect 10966 21270 11284 21298
rect 10966 21200 11022 21270
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 5894 19612 6202 19621
rect 5894 19610 5900 19612
rect 5956 19610 5980 19612
rect 6036 19610 6060 19612
rect 6116 19610 6140 19612
rect 6196 19610 6202 19612
rect 5956 19558 5958 19610
rect 6138 19558 6140 19610
rect 5894 19556 5900 19558
rect 5956 19556 5980 19558
rect 6036 19556 6060 19558
rect 6116 19556 6140 19558
rect 6196 19556 6202 19558
rect 5894 19547 6202 19556
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 4172 18970 4200 19314
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 5276 18766 5304 19314
rect 8036 19310 8064 19654
rect 10839 19612 11147 19621
rect 10839 19610 10845 19612
rect 10901 19610 10925 19612
rect 10981 19610 11005 19612
rect 11061 19610 11085 19612
rect 11141 19610 11147 19612
rect 10901 19558 10903 19610
rect 11083 19558 11085 19610
rect 10839 19556 10845 19558
rect 10901 19556 10925 19558
rect 10981 19556 11005 19558
rect 11061 19556 11085 19558
rect 11141 19556 11147 19558
rect 10839 19547 11147 19556
rect 11256 19446 11284 21270
rect 18234 21200 18290 22000
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8036 18766 8064 19246
rect 8367 19068 8675 19077
rect 8367 19066 8373 19068
rect 8429 19066 8453 19068
rect 8509 19066 8533 19068
rect 8589 19066 8613 19068
rect 8669 19066 8675 19068
rect 8429 19014 8431 19066
rect 8611 19014 8613 19066
rect 8367 19012 8373 19014
rect 8429 19012 8453 19014
rect 8509 19012 8533 19014
rect 8589 19012 8613 19014
rect 8669 19012 8675 19014
rect 8367 19003 8675 19012
rect 11900 18766 11928 19314
rect 13312 19068 13620 19077
rect 13312 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13558 19068
rect 13614 19066 13620 19068
rect 13374 19014 13376 19066
rect 13556 19014 13558 19066
rect 13312 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13558 19014
rect 13614 19012 13620 19014
rect 13312 19003 13620 19012
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 4080 17882 4108 18702
rect 5276 18222 5304 18702
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 5894 18524 6202 18533
rect 5894 18522 5900 18524
rect 5956 18522 5980 18524
rect 6036 18522 6060 18524
rect 6116 18522 6140 18524
rect 6196 18522 6202 18524
rect 5956 18470 5958 18522
rect 6138 18470 6140 18522
rect 5894 18468 5900 18470
rect 5956 18468 5980 18470
rect 6036 18468 6060 18470
rect 6116 18468 6140 18470
rect 6196 18468 6202 18470
rect 5894 18459 6202 18468
rect 7116 18358 7144 18566
rect 7300 18358 7328 18634
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 5276 17678 5304 18158
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3422 16892 3730 16901
rect 3422 16890 3428 16892
rect 3484 16890 3508 16892
rect 3564 16890 3588 16892
rect 3644 16890 3668 16892
rect 3724 16890 3730 16892
rect 3484 16838 3486 16890
rect 3666 16838 3668 16890
rect 3422 16836 3428 16838
rect 3484 16836 3508 16838
rect 3564 16836 3588 16838
rect 3644 16836 3668 16838
rect 3724 16836 3730 16838
rect 3422 16827 3730 16836
rect 5000 16182 5028 17478
rect 5276 16590 5304 17614
rect 7944 17610 7972 18158
rect 8367 17980 8675 17989
rect 8367 17978 8373 17980
rect 8429 17978 8453 17980
rect 8509 17978 8533 17980
rect 8589 17978 8613 17980
rect 8669 17978 8675 17980
rect 8429 17926 8431 17978
rect 8611 17926 8613 17978
rect 8367 17924 8373 17926
rect 8429 17924 8453 17926
rect 8509 17924 8533 17926
rect 8589 17924 8613 17926
rect 8669 17924 8675 17926
rect 8367 17915 8675 17924
rect 9232 17678 9260 18702
rect 10839 18524 11147 18533
rect 10839 18522 10845 18524
rect 10901 18522 10925 18524
rect 10981 18522 11005 18524
rect 11061 18522 11085 18524
rect 11141 18522 11147 18524
rect 10901 18470 10903 18522
rect 11083 18470 11085 18522
rect 10839 18468 10845 18470
rect 10901 18468 10925 18470
rect 10981 18468 11005 18470
rect 11061 18468 11085 18470
rect 11141 18468 11147 18470
rect 10839 18459 11147 18468
rect 11900 18222 11928 18702
rect 13740 18698 13768 19450
rect 14660 19378 14688 19654
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14844 18970 14872 19314
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 15304 18834 15332 19246
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11888 18216 11940 18222
rect 10966 18184 11022 18193
rect 11888 18158 11940 18164
rect 10966 18119 11022 18128
rect 10980 17882 11008 18119
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 5894 17436 6202 17445
rect 5894 17434 5900 17436
rect 5956 17434 5980 17436
rect 6036 17434 6060 17436
rect 6116 17434 6140 17436
rect 6196 17434 6202 17436
rect 5956 17382 5958 17434
rect 6138 17382 6140 17434
rect 5894 17380 5900 17382
rect 5956 17380 5980 17382
rect 6036 17380 6060 17382
rect 6116 17380 6140 17382
rect 6196 17380 6202 17382
rect 5894 17371 6202 17380
rect 7944 17134 7972 17546
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 5276 16046 5304 16526
rect 5894 16348 6202 16357
rect 5894 16346 5900 16348
rect 5956 16346 5980 16348
rect 6036 16346 6060 16348
rect 6116 16346 6140 16348
rect 6196 16346 6202 16348
rect 5956 16294 5958 16346
rect 6138 16294 6140 16346
rect 5894 16292 5900 16294
rect 5956 16292 5980 16294
rect 6036 16292 6060 16294
rect 6116 16292 6140 16294
rect 6196 16292 6202 16294
rect 5894 16283 6202 16292
rect 7944 16114 7972 17070
rect 8367 16892 8675 16901
rect 8367 16890 8373 16892
rect 8429 16890 8453 16892
rect 8509 16890 8533 16892
rect 8589 16890 8613 16892
rect 8669 16890 8675 16892
rect 8429 16838 8431 16890
rect 8611 16838 8613 16890
rect 8367 16836 8373 16838
rect 8429 16836 8453 16838
rect 8509 16836 8533 16838
rect 8589 16836 8613 16838
rect 8669 16836 8675 16838
rect 8367 16827 8675 16836
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 3422 15804 3730 15813
rect 3422 15802 3428 15804
rect 3484 15802 3508 15804
rect 3564 15802 3588 15804
rect 3644 15802 3668 15804
rect 3724 15802 3730 15804
rect 3484 15750 3486 15802
rect 3666 15750 3668 15802
rect 3422 15748 3428 15750
rect 3484 15748 3508 15750
rect 3564 15748 3588 15750
rect 3644 15748 3668 15750
rect 3724 15748 3730 15750
rect 3422 15739 3730 15748
rect 5276 15706 5304 15982
rect 7944 15910 7972 16050
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 6748 15706 6776 15846
rect 8367 15804 8675 15813
rect 8367 15802 8373 15804
rect 8429 15802 8453 15804
rect 8509 15802 8533 15804
rect 8589 15802 8613 15804
rect 8669 15802 8675 15804
rect 8429 15750 8431 15802
rect 8611 15750 8613 15802
rect 8367 15748 8373 15750
rect 8429 15748 8453 15750
rect 8509 15748 8533 15750
rect 8589 15748 8613 15750
rect 8669 15748 8675 15750
rect 8367 15739 8675 15748
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 3422 14716 3730 14725
rect 3422 14714 3428 14716
rect 3484 14714 3508 14716
rect 3564 14714 3588 14716
rect 3644 14714 3668 14716
rect 3724 14714 3730 14716
rect 3484 14662 3486 14714
rect 3666 14662 3668 14714
rect 3422 14660 3428 14662
rect 3484 14660 3508 14662
rect 3564 14660 3588 14662
rect 3644 14660 3668 14662
rect 3724 14660 3730 14662
rect 3422 14651 3730 14660
rect 5828 14618 5856 15438
rect 5894 15260 6202 15269
rect 5894 15258 5900 15260
rect 5956 15258 5980 15260
rect 6036 15258 6060 15260
rect 6116 15258 6140 15260
rect 6196 15258 6202 15260
rect 5956 15206 5958 15258
rect 6138 15206 6140 15258
rect 5894 15204 5900 15206
rect 5956 15204 5980 15206
rect 6036 15204 6060 15206
rect 6116 15204 6140 15206
rect 6196 15204 6202 15206
rect 5894 15195 6202 15204
rect 6748 14958 6776 15642
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6748 14414 6776 14894
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 13394 3280 13670
rect 3422 13628 3730 13637
rect 3422 13626 3428 13628
rect 3484 13626 3508 13628
rect 3564 13626 3588 13628
rect 3644 13626 3668 13628
rect 3724 13626 3730 13628
rect 3484 13574 3486 13626
rect 3666 13574 3668 13626
rect 3422 13572 3428 13574
rect 3484 13572 3508 13574
rect 3564 13572 3588 13574
rect 3644 13572 3668 13574
rect 3724 13572 3730 13574
rect 3422 13563 3730 13572
rect 3988 13530 4016 13806
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 2688 11824 2740 11830
rect 2740 11772 2820 11778
rect 2688 11766 2820 11772
rect 2700 11750 2820 11766
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2332 8090 2360 8434
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 2056 6914 2084 7822
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 1964 6886 2084 6914
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1964 5778 1992 6886
rect 2148 6798 2176 7686
rect 2792 7546 2820 11750
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2884 7410 2912 11630
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 6866 2912 7346
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5914 2084 6258
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2516 5778 2544 6598
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2976 5574 3004 7414
rect 3160 7410 3188 7686
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3252 5710 3280 13330
rect 3422 12540 3730 12549
rect 3422 12538 3428 12540
rect 3484 12538 3508 12540
rect 3564 12538 3588 12540
rect 3644 12538 3668 12540
rect 3724 12538 3730 12540
rect 3484 12486 3486 12538
rect 3666 12486 3668 12538
rect 3422 12484 3428 12486
rect 3484 12484 3508 12486
rect 3564 12484 3588 12486
rect 3644 12484 3668 12486
rect 3724 12484 3730 12486
rect 3422 12475 3730 12484
rect 4080 11898 4108 13806
rect 4172 13462 4200 14282
rect 5448 13864 5500 13870
rect 5552 13818 5580 14350
rect 6932 14346 6960 14758
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 5894 14172 6202 14181
rect 5894 14170 5900 14172
rect 5956 14170 5980 14172
rect 6036 14170 6060 14172
rect 6116 14170 6140 14172
rect 6196 14170 6202 14172
rect 5956 14118 5958 14170
rect 6138 14118 6140 14170
rect 5894 14116 5900 14118
rect 5956 14116 5980 14118
rect 6036 14116 6060 14118
rect 6116 14116 6140 14118
rect 6196 14116 6202 14118
rect 5894 14107 6202 14116
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5500 13812 5580 13818
rect 5448 13806 5580 13812
rect 5460 13790 5580 13806
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 5460 13326 5488 13790
rect 5736 13326 5764 13874
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5460 12306 5488 13262
rect 5894 13084 6202 13093
rect 5894 13082 5900 13084
rect 5956 13082 5980 13084
rect 6036 13082 6060 13084
rect 6116 13082 6140 13084
rect 6196 13082 6202 13084
rect 5956 13030 5958 13082
rect 6138 13030 6140 13082
rect 5894 13028 5900 13030
rect 5956 13028 5980 13030
rect 6036 13028 6060 13030
rect 6116 13028 6140 13030
rect 6196 13028 6202 13030
rect 5894 13019 6202 13028
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12306 6592 12718
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 5460 11762 5488 12242
rect 5894 11996 6202 12005
rect 5894 11994 5900 11996
rect 5956 11994 5980 11996
rect 6036 11994 6060 11996
rect 6116 11994 6140 11996
rect 6196 11994 6202 11996
rect 5956 11942 5958 11994
rect 6138 11942 6140 11994
rect 5894 11940 5900 11942
rect 5956 11940 5980 11942
rect 6036 11940 6060 11942
rect 6116 11940 6140 11942
rect 6196 11940 6202 11942
rect 5894 11931 6202 11940
rect 6564 11762 6592 12242
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 3422 11452 3730 11461
rect 3422 11450 3428 11452
rect 3484 11450 3508 11452
rect 3564 11450 3588 11452
rect 3644 11450 3668 11452
rect 3724 11450 3730 11452
rect 3484 11398 3486 11450
rect 3666 11398 3668 11450
rect 3422 11396 3428 11398
rect 3484 11396 3508 11398
rect 3564 11396 3588 11398
rect 3644 11396 3668 11398
rect 3724 11396 3730 11398
rect 3422 11387 3730 11396
rect 5460 11150 5488 11698
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10606 5488 11086
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 5894 10908 6202 10917
rect 5894 10906 5900 10908
rect 5956 10906 5980 10908
rect 6036 10906 6060 10908
rect 6116 10906 6140 10908
rect 6196 10906 6202 10908
rect 5956 10854 5958 10906
rect 6138 10854 6140 10906
rect 5894 10852 5900 10854
rect 5956 10852 5980 10854
rect 6036 10852 6060 10854
rect 6116 10852 6140 10854
rect 6196 10852 6202 10854
rect 5894 10843 6202 10852
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 3422 10364 3730 10373
rect 3422 10362 3428 10364
rect 3484 10362 3508 10364
rect 3564 10362 3588 10364
rect 3644 10362 3668 10364
rect 3724 10362 3730 10364
rect 3484 10310 3486 10362
rect 3666 10310 3668 10362
rect 3422 10308 3428 10310
rect 3484 10308 3508 10310
rect 3564 10308 3588 10310
rect 3644 10308 3668 10310
rect 3724 10308 3730 10310
rect 3422 10299 3730 10308
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3422 9276 3730 9285
rect 3422 9274 3428 9276
rect 3484 9274 3508 9276
rect 3564 9274 3588 9276
rect 3644 9274 3668 9276
rect 3724 9274 3730 9276
rect 3484 9222 3486 9274
rect 3666 9222 3668 9274
rect 3422 9220 3428 9222
rect 3484 9220 3508 9222
rect 3564 9220 3588 9222
rect 3644 9220 3668 9222
rect 3724 9220 3730 9222
rect 3422 9211 3730 9220
rect 3988 9042 4016 9454
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4172 8634 4200 10542
rect 5276 9994 5304 10542
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9722 5304 9930
rect 5894 9820 6202 9829
rect 5894 9818 5900 9820
rect 5956 9818 5980 9820
rect 6036 9818 6060 9820
rect 6116 9818 6140 9820
rect 6196 9818 6202 9820
rect 5956 9766 5958 9818
rect 6138 9766 6140 9818
rect 5894 9764 5900 9766
rect 5956 9764 5980 9766
rect 6036 9764 6060 9766
rect 6116 9764 6140 9766
rect 6196 9764 6202 9766
rect 5894 9755 6202 9764
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4540 8498 4568 8842
rect 4724 8634 4752 9522
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 3422 8188 3730 8197
rect 3422 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3588 8188
rect 3644 8186 3668 8188
rect 3724 8186 3730 8188
rect 3484 8134 3486 8186
rect 3666 8134 3668 8186
rect 3422 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3588 8134
rect 3644 8132 3668 8134
rect 3724 8132 3730 8134
rect 3422 8123 3730 8132
rect 3422 7100 3730 7109
rect 3422 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3588 7100
rect 3644 7098 3668 7100
rect 3724 7098 3730 7100
rect 3484 7046 3486 7098
rect 3666 7046 3668 7098
rect 3422 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3588 7046
rect 3644 7044 3668 7046
rect 3724 7044 3730 7046
rect 3422 7035 3730 7044
rect 4540 7002 4568 8434
rect 4632 7954 4660 8434
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7750 4752 7822
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 4724 6866 4752 7686
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 3422 6012 3730 6021
rect 3422 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3588 6012
rect 3644 6010 3668 6012
rect 3724 6010 3730 6012
rect 3484 5958 3486 6010
rect 3666 5958 3668 6010
rect 3422 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3588 5958
rect 3644 5956 3668 5958
rect 3724 5956 3730 5958
rect 3422 5947 3730 5956
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 3068 5234 3096 5578
rect 3252 5302 3280 5646
rect 4356 5642 4384 6258
rect 4540 5778 4568 6258
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 4264 5234 4292 5510
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 3422 4924 3730 4933
rect 3422 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3588 4924
rect 3644 4922 3668 4924
rect 3724 4922 3730 4924
rect 3484 4870 3486 4922
rect 3666 4870 3668 4922
rect 3422 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3588 4870
rect 3644 4868 3668 4870
rect 3724 4868 3730 4870
rect 3422 4859 3730 4868
rect 4264 4622 4292 5170
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4356 4146 4384 5578
rect 4540 5370 4568 5714
rect 4632 5710 4660 6190
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4724 5642 4752 6054
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4448 4622 4476 5102
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 4146 4476 4558
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 3422 3836 3730 3845
rect 3422 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3588 3836
rect 3644 3834 3668 3836
rect 3724 3834 3730 3836
rect 3484 3782 3486 3834
rect 3666 3782 3668 3834
rect 3422 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3588 3782
rect 3644 3780 3668 3782
rect 3724 3780 3730 3782
rect 3422 3771 3730 3780
rect 3422 2748 3730 2757
rect 3422 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3588 2748
rect 3644 2746 3668 2748
rect 3724 2746 3730 2748
rect 3484 2694 3486 2746
rect 3666 2694 3668 2746
rect 3422 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3588 2694
rect 3644 2692 3668 2694
rect 3724 2692 3730 2694
rect 3422 2683 3730 2692
rect 4816 2446 4844 8774
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 7886 5580 8502
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 7886 5672 8434
rect 5736 8090 5764 8842
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 5894 8732 6202 8741
rect 5894 8730 5900 8732
rect 5956 8730 5980 8732
rect 6036 8730 6060 8732
rect 6116 8730 6140 8732
rect 6196 8730 6202 8732
rect 5956 8678 5958 8730
rect 6138 8678 6140 8730
rect 5894 8676 5900 8678
rect 5956 8676 5980 8678
rect 6036 8676 6060 8678
rect 6116 8676 6140 8678
rect 6196 8676 6202 8678
rect 5894 8667 6202 8676
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 6012 7886 6040 8434
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5644 7546 5672 7822
rect 5894 7644 6202 7653
rect 5894 7642 5900 7644
rect 5956 7642 5980 7644
rect 6036 7642 6060 7644
rect 6116 7642 6140 7644
rect 6196 7642 6202 7644
rect 5956 7590 5958 7642
rect 6138 7590 6140 7642
rect 5894 7588 5900 7590
rect 5956 7588 5980 7590
rect 6036 7588 6060 7590
rect 6116 7588 6140 7590
rect 6196 7588 6202 7590
rect 5894 7579 6202 7588
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5276 5778 5304 7346
rect 5736 6798 5764 7346
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 6798 6132 7278
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5736 6186 5764 6734
rect 5894 6556 6202 6565
rect 5894 6554 5900 6556
rect 5956 6554 5980 6556
rect 6036 6554 6060 6556
rect 6116 6554 6140 6556
rect 6196 6554 6202 6556
rect 5956 6502 5958 6554
rect 6138 6502 6140 6554
rect 5894 6500 5900 6502
rect 5956 6500 5980 6502
rect 6036 6500 6060 6502
rect 6116 6500 6140 6502
rect 6196 6500 6202 6502
rect 5894 6491 6202 6500
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5920 5914 5948 6190
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5276 5302 5304 5714
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5302 5672 5578
rect 5828 5302 5856 5646
rect 5894 5468 6202 5477
rect 5894 5466 5900 5468
rect 5956 5466 5980 5468
rect 6036 5466 6060 5468
rect 6116 5466 6140 5468
rect 6196 5466 6202 5468
rect 5956 5414 5958 5466
rect 6138 5414 6140 5466
rect 5894 5412 5900 5414
rect 5956 5412 5980 5414
rect 6036 5412 6060 5414
rect 6116 5412 6140 5414
rect 6196 5412 6202 5414
rect 5894 5403 6202 5412
rect 6288 5302 6316 5646
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 4622 6132 5102
rect 6288 4622 6316 5238
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5894 4380 6202 4389
rect 5894 4378 5900 4380
rect 5956 4378 5980 4380
rect 6036 4378 6060 4380
rect 6116 4378 6140 4380
rect 6196 4378 6202 4380
rect 5956 4326 5958 4378
rect 6138 4326 6140 4378
rect 5894 4324 5900 4326
rect 5956 4324 5980 4326
rect 6036 4324 6060 4326
rect 6116 4324 6140 4326
rect 6196 4324 6202 4326
rect 5894 4315 6202 4324
rect 6288 4146 6316 4558
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 5894 3292 6202 3301
rect 5894 3290 5900 3292
rect 5956 3290 5980 3292
rect 6036 3290 6060 3292
rect 6116 3290 6140 3292
rect 6196 3290 6202 3292
rect 5956 3238 5958 3290
rect 6138 3238 6140 3290
rect 5894 3236 5900 3238
rect 5956 3236 5980 3238
rect 6036 3236 6060 3238
rect 6116 3236 6140 3238
rect 6196 3236 6202 3238
rect 5894 3227 6202 3236
rect 6380 2514 6408 8774
rect 6564 8498 6592 9658
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6472 7410 6500 7822
rect 6656 7750 6684 7822
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7410 6684 7686
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6472 7206 6500 7346
rect 6748 7342 6776 8910
rect 6840 7546 6868 11018
rect 6932 8090 6960 12854
rect 7024 10742 7052 15370
rect 8772 15094 8800 17206
rect 9232 17202 9260 17614
rect 10839 17436 11147 17445
rect 10839 17434 10845 17436
rect 10901 17434 10925 17436
rect 10981 17434 11005 17436
rect 11061 17434 11085 17436
rect 11141 17434 11147 17436
rect 10901 17382 10903 17434
rect 11083 17382 11085 17434
rect 10839 17380 10845 17382
rect 10901 17380 10925 17382
rect 10981 17380 11005 17382
rect 11061 17380 11085 17382
rect 11141 17380 11147 17382
rect 10839 17371 11147 17380
rect 11900 17202 11928 18158
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 9232 16114 9260 17138
rect 9416 16794 9444 17138
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 11900 16590 11928 17138
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 10839 16348 11147 16357
rect 10839 16346 10845 16348
rect 10901 16346 10925 16348
rect 10981 16346 11005 16348
rect 11061 16346 11085 16348
rect 11141 16346 11147 16348
rect 10901 16294 10903 16346
rect 11083 16294 11085 16346
rect 10839 16292 10845 16294
rect 10901 16292 10925 16294
rect 10981 16292 11005 16294
rect 11061 16292 11085 16294
rect 11141 16292 11147 16294
rect 10839 16283 11147 16292
rect 9588 16176 9640 16182
rect 9586 16144 9588 16153
rect 9640 16144 9642 16153
rect 9220 16108 9272 16114
rect 9586 16079 9642 16088
rect 9220 16050 9272 16056
rect 11900 16046 11928 16526
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9968 15162 9996 15370
rect 11900 15366 11928 15982
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 10839 15260 11147 15269
rect 10839 15258 10845 15260
rect 10901 15258 10925 15260
rect 10981 15258 11005 15260
rect 11061 15258 11085 15260
rect 11141 15258 11147 15260
rect 10901 15206 10903 15258
rect 11083 15206 11085 15258
rect 10839 15204 10845 15206
rect 10901 15204 10925 15206
rect 10981 15204 11005 15206
rect 11061 15204 11085 15206
rect 11141 15204 11147 15206
rect 10839 15195 11147 15204
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7024 10062 7052 10678
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6798 6500 7142
rect 6748 7002 6776 7278
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 5778 6500 6734
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6656 4826 6684 5578
rect 6748 5574 6776 6190
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5370 6776 5510
rect 6840 5370 6868 5782
rect 6932 5574 6960 6258
rect 7116 5914 7144 15030
rect 11900 14958 11928 15302
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 8367 14716 8675 14725
rect 8367 14714 8373 14716
rect 8429 14714 8453 14716
rect 8509 14714 8533 14716
rect 8589 14714 8613 14716
rect 8669 14714 8675 14716
rect 8429 14662 8431 14714
rect 8611 14662 8613 14714
rect 8367 14660 8373 14662
rect 8429 14660 8453 14662
rect 8509 14660 8533 14662
rect 8589 14660 8613 14662
rect 8669 14660 8675 14662
rect 8367 14651 8675 14660
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10704 14074 10732 14418
rect 11900 14414 11928 14894
rect 12268 14464 12296 18226
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 14646 18184 14702 18193
rect 13312 17980 13620 17989
rect 13312 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13558 17980
rect 13614 17978 13620 17980
rect 13374 17926 13376 17978
rect 13556 17926 13558 17978
rect 13312 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13558 17926
rect 13614 17924 13620 17926
rect 13312 17915 13620 17924
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 16182 12388 16934
rect 13312 16892 13620 16901
rect 13312 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13558 16892
rect 13614 16890 13620 16892
rect 13374 16838 13376 16890
rect 13556 16838 13558 16890
rect 13312 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13558 16838
rect 13614 16836 13620 16838
rect 13312 16827 13620 16836
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12268 14436 12388 14464
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 10839 14172 11147 14181
rect 10839 14170 10845 14172
rect 10901 14170 10925 14172
rect 10981 14170 11005 14172
rect 11061 14170 11085 14172
rect 11141 14170 11147 14172
rect 10901 14118 10903 14170
rect 11083 14118 11085 14170
rect 10839 14116 10845 14118
rect 10901 14116 10925 14118
rect 10981 14116 11005 14118
rect 11061 14116 11085 14118
rect 11141 14116 11147 14118
rect 10839 14107 11147 14116
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 13394 7972 13670
rect 8367 13628 8675 13637
rect 8367 13626 8373 13628
rect 8429 13626 8453 13628
rect 8509 13626 8533 13628
rect 8589 13626 8613 13628
rect 8669 13626 8675 13628
rect 8429 13574 8431 13626
rect 8611 13574 8613 13626
rect 8367 13572 8373 13574
rect 8429 13572 8453 13574
rect 8509 13572 8533 13574
rect 8589 13572 8613 13574
rect 8669 13572 8675 13574
rect 8367 13563 8675 13572
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 8634 7236 11698
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7208 7410 7236 8570
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7410 7420 7754
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 6866 7420 7346
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6390 7420 6802
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7208 5234 7236 6190
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 7300 4758 7328 5170
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 7484 2446 7512 9318
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 5234 7696 5510
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7852 2650 7880 10950
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7944 4690 7972 5102
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8036 2514 8064 12582
rect 8367 12540 8675 12549
rect 8367 12538 8373 12540
rect 8429 12538 8453 12540
rect 8509 12538 8533 12540
rect 8589 12538 8613 12540
rect 8669 12538 8675 12540
rect 8429 12486 8431 12538
rect 8611 12486 8613 12538
rect 8367 12484 8373 12486
rect 8429 12484 8453 12486
rect 8509 12484 8533 12486
rect 8589 12484 8613 12486
rect 8669 12484 8675 12486
rect 8367 12475 8675 12484
rect 9324 12238 9352 13806
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9324 11762 9352 12174
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8367 11452 8675 11461
rect 8367 11450 8373 11452
rect 8429 11450 8453 11452
rect 8509 11450 8533 11452
rect 8589 11450 8613 11452
rect 8669 11450 8675 11452
rect 8429 11398 8431 11450
rect 8611 11398 8613 11450
rect 8367 11396 8373 11398
rect 8429 11396 8453 11398
rect 8509 11396 8533 11398
rect 8589 11396 8613 11398
rect 8669 11396 8675 11398
rect 8367 11387 8675 11396
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8367 10364 8675 10373
rect 8367 10362 8373 10364
rect 8429 10362 8453 10364
rect 8509 10362 8533 10364
rect 8589 10362 8613 10364
rect 8669 10362 8675 10364
rect 8429 10310 8431 10362
rect 8611 10310 8613 10362
rect 8367 10308 8373 10310
rect 8429 10308 8453 10310
rect 8509 10308 8533 10310
rect 8589 10308 8613 10310
rect 8669 10308 8675 10310
rect 8367 10299 8675 10308
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8367 9276 8675 9285
rect 8367 9274 8373 9276
rect 8429 9274 8453 9276
rect 8509 9274 8533 9276
rect 8589 9274 8613 9276
rect 8669 9274 8675 9276
rect 8429 9222 8431 9274
rect 8611 9222 8613 9274
rect 8367 9220 8373 9222
rect 8429 9220 8453 9222
rect 8509 9220 8533 9222
rect 8589 9220 8613 9222
rect 8669 9220 8675 9222
rect 8367 9211 8675 9220
rect 8772 9042 8800 9454
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8367 8188 8675 8197
rect 8367 8186 8373 8188
rect 8429 8186 8453 8188
rect 8509 8186 8533 8188
rect 8589 8186 8613 8188
rect 8669 8186 8675 8188
rect 8429 8134 8431 8186
rect 8611 8134 8613 8186
rect 8367 8132 8373 8134
rect 8429 8132 8453 8134
rect 8509 8132 8533 8134
rect 8589 8132 8613 8134
rect 8669 8132 8675 8134
rect 8367 8123 8675 8132
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7546 8340 7822
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8496 7410 8524 7958
rect 8772 7410 8800 8230
rect 8864 8090 8892 9522
rect 8956 9178 8984 11018
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8956 7886 8984 8910
rect 9048 8090 9076 11630
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6322 8156 7142
rect 8367 7100 8675 7109
rect 8367 7098 8373 7100
rect 8429 7098 8453 7100
rect 8509 7098 8533 7100
rect 8589 7098 8613 7100
rect 8669 7098 8675 7100
rect 8429 7046 8431 7098
rect 8611 7046 8613 7098
rect 8367 7044 8373 7046
rect 8429 7044 8453 7046
rect 8509 7044 8533 7046
rect 8589 7044 8613 7046
rect 8669 7044 8675 7046
rect 8367 7035 8675 7044
rect 9048 6338 9076 7278
rect 8956 6322 9076 6338
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8956 6316 9088 6322
rect 8956 6310 9036 6316
rect 8367 6012 8675 6021
rect 8367 6010 8373 6012
rect 8429 6010 8453 6012
rect 8509 6010 8533 6012
rect 8589 6010 8613 6012
rect 8669 6010 8675 6012
rect 8429 5958 8431 6010
rect 8611 5958 8613 6010
rect 8367 5956 8373 5958
rect 8429 5956 8453 5958
rect 8509 5956 8533 5958
rect 8589 5956 8613 5958
rect 8669 5956 8675 5958
rect 8367 5947 8675 5956
rect 8956 5846 8984 6310
rect 9036 6258 9088 6264
rect 9140 6202 9168 11494
rect 9220 11144 9272 11150
rect 9324 11098 9352 11698
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9272 11092 9352 11098
rect 9220 11086 9352 11092
rect 9232 11070 9352 11086
rect 9324 10470 9352 11070
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10130 9352 10406
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 7818 9260 9522
rect 9324 9518 9352 10066
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9048 6174 9168 6202
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8956 5302 8984 5782
rect 9048 5710 9076 6174
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 9140 5234 9168 6054
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9232 5098 9260 7754
rect 9508 7478 9536 8910
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 6390 9536 7414
rect 9600 7274 9628 8502
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7478 9720 7754
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 6458 9628 7210
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9508 5642 9536 6326
rect 9600 5778 9628 6394
rect 9692 6322 9720 7142
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5166 9536 5578
rect 9600 5234 9628 5714
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4690 8156 4966
rect 8367 4924 8675 4933
rect 8367 4922 8373 4924
rect 8429 4922 8453 4924
rect 8509 4922 8533 4924
rect 8589 4922 8613 4924
rect 8669 4922 8675 4924
rect 8429 4870 8431 4922
rect 8611 4870 8613 4922
rect 8367 4868 8373 4870
rect 8429 4868 8453 4870
rect 8509 4868 8533 4870
rect 8589 4868 8613 4870
rect 8669 4868 8675 4870
rect 8367 4859 8675 4868
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 9508 4622 9536 5102
rect 9600 4690 9628 5170
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 8367 3836 8675 3845
rect 8367 3834 8373 3836
rect 8429 3834 8453 3836
rect 8509 3834 8533 3836
rect 8589 3834 8613 3836
rect 8669 3834 8675 3836
rect 8429 3782 8431 3834
rect 8611 3782 8613 3834
rect 8367 3780 8373 3782
rect 8429 3780 8453 3782
rect 8509 3780 8533 3782
rect 8589 3780 8613 3782
rect 8669 3780 8675 3782
rect 8367 3771 8675 3780
rect 9784 2774 9812 9318
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7274 9904 7822
rect 10152 7750 10180 11494
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7410 10180 7686
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 10244 6322 10272 7890
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5778 10272 6258
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 8367 2748 8675 2757
rect 8367 2746 8373 2748
rect 8429 2746 8453 2748
rect 8509 2746 8533 2748
rect 8589 2746 8613 2748
rect 8669 2746 8675 2748
rect 8429 2694 8431 2746
rect 8611 2694 8613 2746
rect 8367 2692 8373 2694
rect 8429 2692 8453 2694
rect 8509 2692 8533 2694
rect 8589 2692 8613 2694
rect 8669 2692 8675 2694
rect 8367 2683 8675 2692
rect 9692 2746 9812 2774
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 9692 2446 9720 2746
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 1596 800 1624 2314
rect 4264 800 4292 2314
rect 5894 2204 6202 2213
rect 5894 2202 5900 2204
rect 5956 2202 5980 2204
rect 6036 2202 6060 2204
rect 6116 2202 6140 2204
rect 6196 2202 6202 2204
rect 5956 2150 5958 2202
rect 6138 2150 6140 2202
rect 5894 2148 5900 2150
rect 5956 2148 5980 2150
rect 6036 2148 6060 2150
rect 6116 2148 6140 2150
rect 6196 2148 6202 2150
rect 5894 2139 6202 2148
rect 6932 800 6960 2314
rect 10336 2310 10364 11222
rect 10428 6458 10456 13806
rect 11808 13326 11836 13806
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 10839 13084 11147 13093
rect 10839 13082 10845 13084
rect 10901 13082 10925 13084
rect 10981 13082 11005 13084
rect 11061 13082 11085 13084
rect 11141 13082 11147 13084
rect 10901 13030 10903 13082
rect 11083 13030 11085 13082
rect 10839 13028 10845 13030
rect 10901 13028 10925 13030
rect 10981 13028 11005 13030
rect 11061 13028 11085 13030
rect 11141 13028 11147 13030
rect 10839 13019 11147 13028
rect 11808 12782 11836 13262
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 9110 10548 12106
rect 10839 11996 11147 12005
rect 10839 11994 10845 11996
rect 10901 11994 10925 11996
rect 10981 11994 11005 11996
rect 11061 11994 11085 11996
rect 11141 11994 11147 11996
rect 10901 11942 10903 11994
rect 11083 11942 11085 11994
rect 10839 11940 10845 11942
rect 10901 11940 10925 11942
rect 10981 11940 11005 11942
rect 11061 11940 11085 11942
rect 11141 11940 11147 11942
rect 10839 11931 11147 11940
rect 11808 11694 11836 12718
rect 12084 12434 12112 13874
rect 11992 12406 12112 12434
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11150 11836 11630
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 10839 10908 11147 10917
rect 10839 10906 10845 10908
rect 10901 10906 10925 10908
rect 10981 10906 11005 10908
rect 11061 10906 11085 10908
rect 11141 10906 11147 10908
rect 10901 10854 10903 10906
rect 11083 10854 11085 10906
rect 10839 10852 10845 10854
rect 10901 10852 10925 10854
rect 10981 10852 11005 10854
rect 11061 10852 11085 10854
rect 11141 10852 11147 10854
rect 10839 10843 11147 10852
rect 11808 10130 11836 11086
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10612 8090 10640 9930
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 10839 9820 11147 9829
rect 10839 9818 10845 9820
rect 10901 9818 10925 9820
rect 10981 9818 11005 9820
rect 11061 9818 11085 9820
rect 11141 9818 11147 9820
rect 10901 9766 10903 9818
rect 11083 9766 11085 9818
rect 10839 9764 10845 9766
rect 10901 9764 10925 9766
rect 10981 9764 11005 9766
rect 11061 9764 11085 9766
rect 11141 9764 11147 9766
rect 10839 9755 11147 9764
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7546 10640 7822
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10612 6866 10640 7482
rect 10704 7410 10732 9318
rect 10839 8732 11147 8741
rect 10839 8730 10845 8732
rect 10901 8730 10925 8732
rect 10981 8730 11005 8732
rect 11061 8730 11085 8732
rect 11141 8730 11147 8732
rect 10901 8678 10903 8730
rect 11083 8678 11085 8730
rect 10839 8676 10845 8678
rect 10901 8676 10925 8678
rect 10981 8676 11005 8678
rect 11061 8676 11085 8678
rect 11141 8676 11147 8678
rect 10839 8667 11147 8676
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8022 11008 8230
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11060 7880 11112 7886
rect 11058 7848 11060 7857
rect 11440 7857 11468 9862
rect 11808 9586 11836 10066
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11112 7848 11114 7857
rect 11058 7783 11114 7792
rect 11426 7848 11482 7857
rect 11426 7783 11482 7792
rect 10839 7644 11147 7653
rect 10839 7642 10845 7644
rect 10901 7642 10925 7644
rect 10981 7642 11005 7644
rect 11061 7642 11085 7644
rect 11141 7642 11147 7644
rect 10901 7590 10903 7642
rect 11083 7590 11085 7642
rect 10839 7588 10845 7590
rect 10901 7588 10925 7590
rect 10981 7588 11005 7590
rect 11061 7588 11085 7590
rect 11141 7588 11147 7590
rect 10839 7579 11147 7588
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10704 6322 10732 6598
rect 10839 6556 11147 6565
rect 10839 6554 10845 6556
rect 10901 6554 10925 6556
rect 10981 6554 11005 6556
rect 11061 6554 11085 6556
rect 11141 6554 11147 6556
rect 10901 6502 10903 6554
rect 11083 6502 11085 6554
rect 10839 6500 10845 6502
rect 10901 6500 10925 6502
rect 10981 6500 11005 6502
rect 11061 6500 11085 6502
rect 11141 6500 11147 6502
rect 10839 6491 11147 6500
rect 11256 6322 11284 6734
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5846 10640 6054
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 11164 5710 11192 6190
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10839 5468 11147 5477
rect 10839 5466 10845 5468
rect 10901 5466 10925 5468
rect 10981 5466 11005 5468
rect 11061 5466 11085 5468
rect 11141 5466 11147 5468
rect 10901 5414 10903 5466
rect 11083 5414 11085 5466
rect 10839 5412 10845 5414
rect 10901 5412 10925 5414
rect 10981 5412 11005 5414
rect 11061 5412 11085 5414
rect 11141 5412 11147 5414
rect 10839 5403 11147 5412
rect 11992 5098 12020 12406
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 7886 12112 11018
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 8634 12204 9522
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8514 12296 14282
rect 12360 12238 12388 14436
rect 12728 12434 12756 16390
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13096 14074 13124 14486
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12728 12406 12940 12434
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12176 8486 12296 8514
rect 12624 8492 12676 8498
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12176 5166 12204 8486
rect 12624 8434 12676 8440
rect 12636 8378 12664 8434
rect 12544 8350 12664 8378
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12360 7478 12388 7958
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12452 7342 12480 7754
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12268 7002 12296 7278
rect 12544 7274 12572 8350
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8090 12664 8230
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12636 7750 12664 7890
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12256 6248 12308 6254
rect 12728 6202 12756 11698
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8022 12848 8230
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12820 6866 12848 7278
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6662 12848 6802
rect 12912 6730 12940 12406
rect 13188 8090 13216 16458
rect 13312 15804 13620 15813
rect 13312 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13558 15804
rect 13614 15802 13620 15804
rect 13374 15750 13376 15802
rect 13556 15750 13558 15802
rect 13312 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13558 15750
rect 13614 15748 13620 15750
rect 13312 15739 13620 15748
rect 13312 14716 13620 14725
rect 13312 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13558 14716
rect 13614 14714 13620 14716
rect 13374 14662 13376 14714
rect 13556 14662 13558 14714
rect 13312 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13558 14662
rect 13614 14660 13620 14662
rect 13312 14651 13620 14660
rect 13312 13628 13620 13637
rect 13312 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13558 13628
rect 13614 13626 13620 13628
rect 13374 13574 13376 13626
rect 13556 13574 13558 13626
rect 13312 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13558 13574
rect 13614 13572 13620 13574
rect 13312 13563 13620 13572
rect 13312 12540 13620 12549
rect 13312 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13558 12540
rect 13614 12538 13620 12540
rect 13374 12486 13376 12538
rect 13556 12486 13558 12538
rect 13312 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13558 12486
rect 13614 12484 13620 12486
rect 13312 12475 13620 12484
rect 13312 11452 13620 11461
rect 13312 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13558 11452
rect 13614 11450 13620 11452
rect 13374 11398 13376 11450
rect 13556 11398 13558 11450
rect 13312 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13558 11398
rect 13614 11396 13620 11398
rect 13312 11387 13620 11396
rect 13312 10364 13620 10373
rect 13312 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13558 10364
rect 13614 10362 13620 10364
rect 13374 10310 13376 10362
rect 13556 10310 13558 10362
rect 13312 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13558 10310
rect 13614 10308 13620 10310
rect 13312 10299 13620 10308
rect 13312 9276 13620 9285
rect 13312 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13558 9276
rect 13614 9274 13620 9276
rect 13374 9222 13376 9274
rect 13556 9222 13558 9274
rect 13312 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13558 9222
rect 13614 9220 13620 9222
rect 13312 9211 13620 9220
rect 13312 8188 13620 8197
rect 13312 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13558 8188
rect 13614 8186 13620 8188
rect 13374 8134 13376 8186
rect 13556 8134 13558 8186
rect 13312 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13558 8134
rect 13614 8132 13620 8134
rect 13312 8123 13620 8132
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13648 7954 13676 18158
rect 14646 18119 14702 18128
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13740 13870 13768 16050
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14016 11150 14044 14758
rect 14384 14482 14412 18022
rect 14568 17678 14596 18022
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15570 14504 15846
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14568 15162 14596 16050
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7546 13216 7822
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13280 7256 13308 7890
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7410 13584 7822
rect 13740 7818 13768 8366
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13188 7228 13308 7256
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12256 6190 12308 6196
rect 12268 5234 12296 6190
rect 12636 6174 12756 6202
rect 12636 5914 12664 6174
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12728 5574 12756 6054
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5302 12756 5510
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 12728 4826 12756 5238
rect 13096 5148 13124 6258
rect 13188 5846 13216 7228
rect 13312 7100 13620 7109
rect 13312 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13558 7100
rect 13614 7098 13620 7100
rect 13374 7046 13376 7098
rect 13556 7046 13558 7098
rect 13312 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13558 7046
rect 13614 7044 13620 7046
rect 13312 7035 13620 7044
rect 13740 6798 13768 7482
rect 13832 7342 13860 9318
rect 14016 8906 14044 11086
rect 14108 9586 14136 12582
rect 14568 12170 14596 14214
rect 14660 13326 14688 18119
rect 14844 15978 14872 18770
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14936 18222 14964 18634
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 15028 17202 15056 18566
rect 15212 17338 15240 18566
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15304 17270 15332 18770
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15396 17626 15424 18294
rect 15488 18086 15516 18770
rect 15672 18272 15700 19654
rect 15784 19612 16092 19621
rect 15784 19610 15790 19612
rect 15846 19610 15870 19612
rect 15926 19610 15950 19612
rect 16006 19610 16030 19612
rect 16086 19610 16092 19612
rect 15846 19558 15848 19610
rect 16028 19558 16030 19610
rect 15784 19556 15790 19558
rect 15846 19556 15870 19558
rect 15926 19556 15950 19558
rect 16006 19556 16030 19558
rect 16086 19556 16092 19558
rect 15784 19547 16092 19556
rect 18248 19446 18276 21200
rect 20729 19612 21037 19621
rect 20729 19610 20735 19612
rect 20791 19610 20815 19612
rect 20871 19610 20895 19612
rect 20951 19610 20975 19612
rect 21031 19610 21037 19612
rect 20791 19558 20793 19610
rect 20973 19558 20975 19610
rect 20729 19556 20735 19558
rect 20791 19556 20815 19558
rect 20871 19556 20895 19558
rect 20951 19556 20975 19558
rect 21031 19556 21037 19558
rect 20729 19547 21037 19556
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15784 18524 16092 18533
rect 15784 18522 15790 18524
rect 15846 18522 15870 18524
rect 15926 18522 15950 18524
rect 16006 18522 16030 18524
rect 16086 18522 16092 18524
rect 15846 18470 15848 18522
rect 16028 18470 16030 18522
rect 15784 18468 15790 18470
rect 15846 18468 15870 18470
rect 15926 18468 15950 18470
rect 16006 18468 16030 18470
rect 16086 18468 16092 18470
rect 15784 18459 16092 18468
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15672 18244 15792 18272
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15488 17746 15516 18022
rect 15580 17882 15608 18022
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15764 17814 15792 18244
rect 15856 18193 15884 18362
rect 16132 18358 16160 18906
rect 16120 18352 16172 18358
rect 16172 18312 16252 18340
rect 16120 18294 16172 18300
rect 16120 18216 16172 18222
rect 15842 18184 15898 18193
rect 16120 18158 16172 18164
rect 15842 18119 15898 18128
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15396 17610 15516 17626
rect 15396 17604 15528 17610
rect 15396 17598 15476 17604
rect 15476 17546 15528 17552
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 17082 15056 17138
rect 14936 17054 15056 17082
rect 15200 17060 15252 17066
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14936 14890 14964 17054
rect 15200 17002 15252 17008
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16658 15056 16934
rect 15212 16726 15240 17002
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 15026 15056 16594
rect 15212 15026 15240 16662
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14660 12442 14688 12786
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10266 14228 10406
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13464 6458 13492 6666
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13312 6012 13620 6021
rect 13312 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13558 6012
rect 13614 6010 13620 6012
rect 13374 5958 13376 6010
rect 13556 5958 13558 6010
rect 13312 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13558 5958
rect 13614 5956 13620 5958
rect 13312 5947 13620 5956
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13188 5642 13216 5782
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13648 5234 13676 6394
rect 13740 6390 13768 6734
rect 14016 6458 14044 8842
rect 14200 7002 14228 9318
rect 14292 9178 14320 11766
rect 14660 11762 14688 12378
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14476 9586 14504 10406
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14568 9518 14596 10406
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 14016 6322 14044 6394
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14200 5234 14228 6938
rect 14292 6390 14320 9114
rect 14476 8566 14504 9318
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14568 6798 14596 8978
rect 14660 8906 14688 11494
rect 14752 9654 14780 14758
rect 14844 14618 14872 14758
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 12782 14872 14010
rect 15212 13410 15240 14962
rect 15304 13530 15332 17206
rect 15488 17202 15516 17546
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15580 16658 15608 17682
rect 15784 17436 16092 17445
rect 15784 17434 15790 17436
rect 15846 17434 15870 17436
rect 15926 17434 15950 17436
rect 16006 17434 16030 17436
rect 16086 17434 16092 17436
rect 15846 17382 15848 17434
rect 16028 17382 16030 17434
rect 15784 17380 15790 17382
rect 15846 17380 15870 17382
rect 15926 17380 15950 17382
rect 16006 17380 16030 17382
rect 16086 17380 16092 17382
rect 15784 17371 16092 17380
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 16132 16590 16160 18158
rect 16224 18154 16252 18312
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16868 18193 16896 18226
rect 16854 18184 16910 18193
rect 16212 18148 16264 18154
rect 16960 18154 16988 19314
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17052 18970 17080 19110
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17052 18766 17080 18906
rect 17144 18834 17172 19382
rect 17788 18834 17816 19382
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16854 18119 16910 18128
rect 16948 18148 17000 18154
rect 16212 18090 16264 18096
rect 16948 18090 17000 18096
rect 17052 17610 17080 18294
rect 17144 17678 17172 18770
rect 17236 17882 17264 18770
rect 17972 18630 18000 19382
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 18064 18426 18092 19110
rect 18257 19068 18565 19077
rect 18257 19066 18263 19068
rect 18319 19066 18343 19068
rect 18399 19066 18423 19068
rect 18479 19066 18503 19068
rect 18559 19066 18565 19068
rect 18319 19014 18321 19066
rect 18501 19014 18503 19066
rect 18257 19012 18263 19014
rect 18319 19012 18343 19014
rect 18399 19012 18423 19014
rect 18479 19012 18503 19014
rect 18559 19012 18565 19014
rect 18257 19003 18565 19012
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17604 17678 17632 18226
rect 18257 17980 18565 17989
rect 18257 17978 18263 17980
rect 18319 17978 18343 17980
rect 18399 17978 18423 17980
rect 18479 17978 18503 17980
rect 18559 17978 18565 17980
rect 18319 17926 18321 17978
rect 18501 17926 18503 17978
rect 18257 17924 18263 17926
rect 18319 17924 18343 17926
rect 18399 17924 18423 17926
rect 18479 17924 18503 17926
rect 18559 17924 18565 17926
rect 18257 17915 18565 17924
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15784 16348 16092 16357
rect 15784 16346 15790 16348
rect 15846 16346 15870 16348
rect 15926 16346 15950 16348
rect 16006 16346 16030 16348
rect 16086 16346 16092 16348
rect 15846 16294 15848 16346
rect 16028 16294 16030 16346
rect 15784 16292 15790 16294
rect 15846 16292 15870 16294
rect 15926 16292 15950 16294
rect 16006 16292 16030 16294
rect 16086 16292 16092 16294
rect 15784 16283 16092 16292
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15212 13382 15332 13410
rect 15304 13326 15332 13382
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14844 8974 14872 12718
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14936 10554 14964 12106
rect 15028 11286 15056 13126
rect 15120 12782 15148 13262
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 12374 15148 12582
rect 15212 12442 15240 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15304 11354 15332 12922
rect 15396 11626 15424 15846
rect 15672 15162 15700 16050
rect 16316 15978 16344 16594
rect 16408 16250 16436 17138
rect 16592 16726 16620 17138
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16794 16712 17070
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16776 16726 16804 16934
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16592 16250 16620 16662
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16408 15978 16436 16186
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 15784 15260 16092 15269
rect 15784 15258 15790 15260
rect 15846 15258 15870 15260
rect 15926 15258 15950 15260
rect 16006 15258 16030 15260
rect 16086 15258 16092 15260
rect 15846 15206 15848 15258
rect 16028 15206 16030 15258
rect 15784 15204 15790 15206
rect 15846 15204 15870 15206
rect 15926 15204 15950 15206
rect 16006 15204 16030 15206
rect 16086 15204 16092 15206
rect 15784 15195 16092 15204
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 16408 14958 16436 15914
rect 16684 15638 16712 16458
rect 16868 16114 16896 16526
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15706 16896 16050
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 15672 14618 15700 14894
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15488 11801 15516 14418
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15028 10742 15056 11222
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10810 15240 11018
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15108 10600 15160 10606
rect 14936 10526 15056 10554
rect 15108 10542 15160 10548
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 8090 14688 8434
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14568 6390 14596 6734
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14384 5846 14412 6190
rect 14476 5914 14504 6326
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14476 5642 14504 5850
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13176 5160 13228 5166
rect 13096 5120 13176 5148
rect 13176 5102 13228 5108
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13188 4622 13216 5102
rect 13372 5030 13400 5102
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13312 4924 13620 4933
rect 13312 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13558 4924
rect 13614 4922 13620 4924
rect 13374 4870 13376 4922
rect 13556 4870 13558 4922
rect 13312 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13558 4870
rect 13614 4868 13620 4870
rect 13312 4859 13620 4868
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13740 4554 13768 5102
rect 14476 5030 14504 5578
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4622 14504 4966
rect 14660 4690 14688 5646
rect 14752 4758 14780 8366
rect 14844 6254 14872 8910
rect 14936 8566 14964 9998
rect 15028 9042 15056 10526
rect 15120 10130 15148 10542
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 9994 15240 10202
rect 15304 10130 15332 11290
rect 15488 10674 15516 11727
rect 15580 11626 15608 13126
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15672 10470 15700 14418
rect 15784 14172 16092 14181
rect 15784 14170 15790 14172
rect 15846 14170 15870 14172
rect 15926 14170 15950 14172
rect 16006 14170 16030 14172
rect 16086 14170 16092 14172
rect 15846 14118 15848 14170
rect 16028 14118 16030 14170
rect 15784 14116 15790 14118
rect 15846 14116 15870 14118
rect 15926 14116 15950 14118
rect 16006 14116 16030 14118
rect 16086 14116 16092 14118
rect 15784 14107 16092 14116
rect 15784 13084 16092 13093
rect 15784 13082 15790 13084
rect 15846 13082 15870 13084
rect 15926 13082 15950 13084
rect 16006 13082 16030 13084
rect 16086 13082 16092 13084
rect 15846 13030 15848 13082
rect 16028 13030 16030 13082
rect 15784 13028 15790 13030
rect 15846 13028 15870 13030
rect 15926 13028 15950 13030
rect 16006 13028 16030 13030
rect 16086 13028 16092 13030
rect 15784 13019 16092 13028
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 15784 11996 16092 12005
rect 15784 11994 15790 11996
rect 15846 11994 15870 11996
rect 15926 11994 15950 11996
rect 16006 11994 16030 11996
rect 16086 11994 16092 11996
rect 15846 11942 15848 11994
rect 16028 11942 16030 11994
rect 15784 11940 15790 11942
rect 15846 11940 15870 11942
rect 15926 11940 15950 11942
rect 16006 11940 16030 11942
rect 16086 11940 16092 11942
rect 15784 11931 16092 11940
rect 15784 10908 16092 10917
rect 15784 10906 15790 10908
rect 15846 10906 15870 10908
rect 15926 10906 15950 10908
rect 16006 10906 16030 10908
rect 16086 10906 16092 10908
rect 15846 10854 15848 10906
rect 16028 10854 16030 10906
rect 15784 10852 15790 10854
rect 15846 10852 15870 10854
rect 15926 10852 15950 10854
rect 16006 10852 16030 10854
rect 16086 10852 16092 10854
rect 15784 10843 16092 10852
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9450 15148 9862
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14936 7274 14964 8502
rect 15028 8498 15056 8774
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15212 7478 15240 9930
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8906 15332 9318
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15304 7410 15332 7822
rect 15396 7546 15424 8026
rect 15672 7954 15700 10406
rect 15784 9820 16092 9829
rect 15784 9818 15790 9820
rect 15846 9818 15870 9820
rect 15926 9818 15950 9820
rect 16006 9818 16030 9820
rect 16086 9818 16092 9820
rect 15846 9766 15848 9818
rect 16028 9766 16030 9818
rect 15784 9764 15790 9766
rect 15846 9764 15870 9766
rect 15926 9764 15950 9766
rect 16006 9764 16030 9766
rect 16086 9764 16092 9766
rect 15784 9755 16092 9764
rect 15784 8732 16092 8741
rect 15784 8730 15790 8732
rect 15846 8730 15870 8732
rect 15926 8730 15950 8732
rect 16006 8730 16030 8732
rect 16086 8730 16092 8732
rect 15846 8678 15848 8730
rect 16028 8678 16030 8730
rect 15784 8676 15790 8678
rect 15846 8676 15870 8678
rect 15926 8676 15950 8678
rect 16006 8676 16030 8678
rect 16086 8676 16092 8678
rect 15784 8667 16092 8676
rect 16132 8090 16160 12718
rect 16684 12434 16712 15574
rect 17144 14906 17172 17614
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17328 15706 17356 16186
rect 17420 16114 17448 17138
rect 17512 16658 17540 17206
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17052 14878 17172 14906
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13938 16988 14350
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16960 13394 16988 13874
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16592 12406 16712 12434
rect 16592 9466 16620 12406
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16500 9438 16620 9466
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16500 7954 16528 9438
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 15028 6866 15056 7278
rect 15120 7206 15148 7346
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15120 6798 15148 7142
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15304 6662 15332 7346
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 15304 5778 15332 6598
rect 15396 6322 15424 7482
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15672 6186 15700 7890
rect 15784 7644 16092 7653
rect 15784 7642 15790 7644
rect 15846 7642 15870 7644
rect 15926 7642 15950 7644
rect 16006 7642 16030 7644
rect 16086 7642 16092 7644
rect 15846 7590 15848 7642
rect 16028 7590 16030 7642
rect 15784 7588 15790 7590
rect 15846 7588 15870 7590
rect 15926 7588 15950 7590
rect 16006 7588 16030 7590
rect 16086 7588 16092 7590
rect 15784 7579 16092 7588
rect 16500 7478 16528 7890
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 15784 6556 16092 6565
rect 15784 6554 15790 6556
rect 15846 6554 15870 6556
rect 15926 6554 15950 6556
rect 16006 6554 16030 6556
rect 16086 6554 16092 6556
rect 15846 6502 15848 6554
rect 16028 6502 16030 6554
rect 15784 6500 15790 6502
rect 15846 6500 15870 6502
rect 15926 6500 15950 6502
rect 16006 6500 16030 6502
rect 16086 6500 16092 6502
rect 15784 6491 16092 6500
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15396 5234 15424 6054
rect 15784 5468 16092 5477
rect 15784 5466 15790 5468
rect 15846 5466 15870 5468
rect 15926 5466 15950 5468
rect 16006 5466 16030 5468
rect 16086 5466 16092 5468
rect 15846 5414 15848 5466
rect 16028 5414 16030 5466
rect 15784 5412 15790 5414
rect 15846 5412 15870 5414
rect 15926 5412 15950 5414
rect 16006 5412 16030 5414
rect 16086 5412 16092 5414
rect 15784 5403 16092 5412
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15212 4826 15240 5170
rect 16132 5098 16160 7346
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 16500 4622 16528 7414
rect 16592 5302 16620 8842
rect 16684 8566 16712 11698
rect 16776 10810 16804 12854
rect 16960 12850 16988 13330
rect 17052 13326 17080 14878
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14414 17172 14758
rect 17132 14408 17184 14414
rect 17184 14356 17264 14362
rect 17132 14350 17264 14356
rect 17144 14334 17264 14350
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 13734 17172 14214
rect 17236 13938 17264 14334
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12238 16988 12582
rect 17144 12238 17172 13126
rect 17236 12850 17264 13262
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11762 17080 12038
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 11354 16896 11562
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 17052 10742 17080 11698
rect 17236 11558 17264 11698
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17236 11218 17264 11494
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17052 10062 17080 10678
rect 17236 10554 17264 11154
rect 17328 10674 17356 15506
rect 17420 15502 17448 16050
rect 17512 16046 17540 16594
rect 17604 16250 17632 17614
rect 18257 16892 18565 16901
rect 18257 16890 18263 16892
rect 18319 16890 18343 16892
rect 18399 16890 18423 16892
rect 18479 16890 18503 16892
rect 18559 16890 18565 16892
rect 18319 16838 18321 16890
rect 18501 16838 18503 16890
rect 18257 16836 18263 16838
rect 18319 16836 18343 16838
rect 18399 16836 18423 16838
rect 18479 16836 18503 16838
rect 18559 16836 18565 16838
rect 18257 16827 18565 16836
rect 19260 16658 19288 18566
rect 20729 18524 21037 18533
rect 20729 18522 20735 18524
rect 20791 18522 20815 18524
rect 20871 18522 20895 18524
rect 20951 18522 20975 18524
rect 21031 18522 21037 18524
rect 20791 18470 20793 18522
rect 20973 18470 20975 18522
rect 20729 18468 20735 18470
rect 20791 18468 20815 18470
rect 20871 18468 20895 18470
rect 20951 18468 20975 18470
rect 21031 18468 21037 18470
rect 20729 18459 21037 18468
rect 20729 17436 21037 17445
rect 20729 17434 20735 17436
rect 20791 17434 20815 17436
rect 20871 17434 20895 17436
rect 20951 17434 20975 17436
rect 21031 17434 21037 17436
rect 20791 17382 20793 17434
rect 20973 17382 20975 17434
rect 20729 17380 20735 17382
rect 20791 17380 20815 17382
rect 20871 17380 20895 17382
rect 20951 17380 20975 17382
rect 21031 17380 21037 17382
rect 20729 17371 21037 17380
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17512 15434 17540 15982
rect 17788 15638 17816 16458
rect 18892 16114 18920 16526
rect 19720 16454 19748 16526
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18257 15804 18565 15813
rect 18257 15802 18263 15804
rect 18319 15802 18343 15804
rect 18399 15802 18423 15804
rect 18479 15802 18503 15804
rect 18559 15802 18565 15804
rect 18319 15750 18321 15802
rect 18501 15750 18503 15802
rect 18257 15748 18263 15750
rect 18319 15748 18343 15750
rect 18399 15748 18423 15750
rect 18479 15748 18503 15750
rect 18559 15748 18565 15750
rect 18257 15739 18565 15748
rect 19720 15706 19748 16390
rect 19812 16250 19840 16526
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 20088 16153 20116 16390
rect 20729 16348 21037 16357
rect 20729 16346 20735 16348
rect 20791 16346 20815 16348
rect 20871 16346 20895 16348
rect 20951 16346 20975 16348
rect 21031 16346 21037 16348
rect 20791 16294 20793 16346
rect 20973 16294 20975 16346
rect 20729 16292 20735 16294
rect 20791 16292 20815 16294
rect 20871 16292 20895 16294
rect 20951 16292 20975 16294
rect 21031 16292 21037 16294
rect 20729 16283 21037 16292
rect 20074 16144 20130 16153
rect 20074 16079 20130 16088
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17420 14006 17448 14350
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17420 12918 17448 13262
rect 17696 12986 17724 14962
rect 17972 14278 18000 15030
rect 18064 14618 18092 15302
rect 18156 14890 18184 15302
rect 19352 15094 19380 15506
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19536 15162 19564 15370
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18156 14346 18184 14826
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 18257 14716 18565 14725
rect 18257 14714 18263 14716
rect 18319 14714 18343 14716
rect 18399 14714 18423 14716
rect 18479 14714 18503 14716
rect 18559 14714 18565 14716
rect 18319 14662 18321 14714
rect 18501 14662 18503 14714
rect 18257 14660 18263 14662
rect 18319 14660 18343 14662
rect 18399 14660 18423 14662
rect 18479 14660 18503 14662
rect 18559 14660 18565 14662
rect 18257 14651 18565 14660
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17960 14272 18012 14278
rect 17788 14232 17960 14260
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17408 12912 17460 12918
rect 17788 12866 17816 14232
rect 17960 14214 18012 14220
rect 19168 13938 19196 14758
rect 19352 14414 19380 15030
rect 19536 15026 19564 15098
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 18257 13628 18565 13637
rect 18257 13626 18263 13628
rect 18319 13626 18343 13628
rect 18399 13626 18423 13628
rect 18479 13626 18503 13628
rect 18559 13626 18565 13628
rect 18319 13574 18321 13626
rect 18501 13574 18503 13626
rect 18257 13572 18263 13574
rect 18319 13572 18343 13574
rect 18399 13572 18423 13574
rect 18479 13572 18503 13574
rect 18559 13572 18565 13574
rect 18257 13563 18565 13572
rect 18616 12918 18644 13874
rect 17408 12854 17460 12860
rect 17696 12838 17816 12866
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 19168 12850 19196 13874
rect 19352 13326 19380 14214
rect 19444 14074 19472 14214
rect 19536 14074 19564 14962
rect 19720 14958 19748 15302
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19432 13932 19484 13938
rect 19484 13892 19564 13920
rect 19432 13874 19484 13880
rect 19536 13802 19564 13892
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 17960 12844 18012 12850
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17420 11898 17448 12174
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17512 11694 17540 12038
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17144 10526 17264 10554
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17144 9654 17172 10526
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16868 8498 16896 9454
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8634 16988 8910
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 6934 16896 8434
rect 17052 8430 17080 9114
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17052 8090 17080 8366
rect 17144 8362 17172 9590
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 17236 6866 17264 10406
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17328 7818 17356 8434
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16776 6390 16804 6734
rect 16868 6458 16896 6734
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16776 5778 16804 6326
rect 17236 6254 17264 6802
rect 17420 6730 17448 11086
rect 17512 10674 17540 11154
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17696 9602 17724 12838
rect 17960 12786 18012 12792
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 17972 12306 18000 12786
rect 19444 12714 19472 13194
rect 19536 13190 19564 13738
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 18257 12540 18565 12549
rect 18257 12538 18263 12540
rect 18319 12538 18343 12540
rect 18399 12538 18423 12540
rect 18479 12538 18503 12540
rect 18559 12538 18565 12540
rect 18319 12486 18321 12538
rect 18501 12486 18503 12538
rect 18257 12484 18263 12486
rect 18319 12484 18343 12486
rect 18399 12484 18423 12486
rect 18479 12484 18503 12486
rect 18559 12484 18565 12486
rect 18257 12475 18565 12484
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11898 17908 12106
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18064 11762 18092 12038
rect 19536 11898 19564 13126
rect 19628 12782 19656 14554
rect 19812 14482 19840 14758
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19720 14074 19748 14214
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19904 13802 19932 15982
rect 20729 15260 21037 15269
rect 20729 15258 20735 15260
rect 20791 15258 20815 15260
rect 20871 15258 20895 15260
rect 20951 15258 20975 15260
rect 21031 15258 21037 15260
rect 20791 15206 20793 15258
rect 20973 15206 20975 15258
rect 20729 15204 20735 15206
rect 20791 15204 20815 15206
rect 20871 15204 20895 15206
rect 20951 15204 20975 15206
rect 21031 15204 21037 15206
rect 20729 15195 21037 15204
rect 20729 14172 21037 14181
rect 20729 14170 20735 14172
rect 20791 14170 20815 14172
rect 20871 14170 20895 14172
rect 20951 14170 20975 14172
rect 21031 14170 21037 14172
rect 20791 14118 20793 14170
rect 20973 14118 20975 14170
rect 20729 14116 20735 14118
rect 20791 14116 20815 14118
rect 20871 14116 20895 14118
rect 20951 14116 20975 14118
rect 21031 14116 21037 14118
rect 20729 14107 21037 14116
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 20729 13084 21037 13093
rect 20729 13082 20735 13084
rect 20791 13082 20815 13084
rect 20871 13082 20895 13084
rect 20951 13082 20975 13084
rect 21031 13082 21037 13084
rect 20791 13030 20793 13082
rect 20973 13030 20975 13082
rect 20729 13028 20735 13030
rect 20791 13028 20815 13030
rect 20871 13028 20895 13030
rect 20951 13028 20975 13030
rect 21031 13028 21037 13030
rect 20729 13019 21037 13028
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 12442 19656 12718
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19246 11792 19302 11801
rect 18052 11756 18104 11762
rect 19246 11727 19248 11736
rect 18052 11698 18104 11704
rect 19300 11727 19302 11736
rect 19340 11756 19392 11762
rect 19248 11698 19300 11704
rect 19340 11698 19392 11704
rect 18064 10826 18092 11698
rect 18257 11452 18565 11461
rect 18257 11450 18263 11452
rect 18319 11450 18343 11452
rect 18399 11450 18423 11452
rect 18479 11450 18503 11452
rect 18559 11450 18565 11452
rect 18319 11398 18321 11450
rect 18501 11398 18503 11450
rect 18257 11396 18263 11398
rect 18319 11396 18343 11398
rect 18399 11396 18423 11398
rect 18479 11396 18503 11398
rect 18559 11396 18565 11398
rect 18257 11387 18565 11396
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18064 10798 18184 10826
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17788 10606 17816 10678
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17604 9574 17724 9602
rect 17512 9178 17540 9522
rect 17604 9450 17632 9574
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17696 9178 17724 9454
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17052 4690 17080 5102
rect 17512 5030 17540 8910
rect 17604 8634 17632 9046
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17604 8022 17632 8366
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17604 7818 17632 7958
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17696 7750 17724 8366
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 5846 17724 7686
rect 17788 7546 17816 10542
rect 18064 9450 18092 10678
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8498 17908 8774
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 7886 18000 8230
rect 18156 7954 18184 10798
rect 18708 10742 18736 11086
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18708 10470 18736 10678
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18257 10364 18565 10373
rect 18257 10362 18263 10364
rect 18319 10362 18343 10364
rect 18399 10362 18423 10364
rect 18479 10362 18503 10364
rect 18559 10362 18565 10364
rect 18319 10310 18321 10362
rect 18501 10310 18503 10362
rect 18257 10308 18263 10310
rect 18319 10308 18343 10310
rect 18399 10308 18423 10310
rect 18479 10308 18503 10310
rect 18559 10308 18565 10310
rect 18257 10299 18565 10308
rect 19260 10198 19288 11698
rect 19352 11150 19380 11698
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10810 19380 11086
rect 19628 11082 19656 12378
rect 19996 12238 20024 12582
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19720 11898 19748 12038
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19444 10010 19472 10950
rect 19628 10606 19656 11018
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19996 10266 20024 12174
rect 20729 11996 21037 12005
rect 20729 11994 20735 11996
rect 20791 11994 20815 11996
rect 20871 11994 20895 11996
rect 20951 11994 20975 11996
rect 21031 11994 21037 11996
rect 20791 11942 20793 11994
rect 20973 11942 20975 11994
rect 20729 11940 20735 11942
rect 20791 11940 20815 11942
rect 20871 11940 20895 11942
rect 20951 11940 20975 11942
rect 21031 11940 21037 11942
rect 20729 11931 21037 11940
rect 20729 10908 21037 10917
rect 20729 10906 20735 10908
rect 20791 10906 20815 10908
rect 20871 10906 20895 10908
rect 20951 10906 20975 10908
rect 21031 10906 21037 10908
rect 20791 10854 20793 10906
rect 20973 10854 20975 10906
rect 20729 10852 20735 10854
rect 20791 10852 20815 10854
rect 20871 10852 20895 10854
rect 20951 10852 20975 10854
rect 21031 10852 21037 10854
rect 20729 10843 21037 10852
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19352 9994 19472 10010
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19340 9988 19472 9994
rect 19392 9982 19472 9988
rect 19340 9930 19392 9936
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 18257 9276 18565 9285
rect 18257 9274 18263 9276
rect 18319 9274 18343 9276
rect 18399 9274 18423 9276
rect 18479 9274 18503 9276
rect 18559 9274 18565 9276
rect 18319 9222 18321 9274
rect 18501 9222 18503 9274
rect 18257 9220 18263 9222
rect 18319 9220 18343 9222
rect 18399 9220 18423 9222
rect 18479 9220 18503 9222
rect 18559 9220 18565 9222
rect 18257 9211 18565 9220
rect 19168 8974 19196 9590
rect 19628 9586 19656 9998
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19812 9722 19840 9862
rect 20088 9722 20116 10610
rect 20729 9820 21037 9829
rect 20729 9818 20735 9820
rect 20791 9818 20815 9820
rect 20871 9818 20895 9820
rect 20951 9818 20975 9820
rect 21031 9818 21037 9820
rect 20791 9766 20793 9818
rect 20973 9766 20975 9818
rect 20729 9764 20735 9766
rect 20791 9764 20815 9766
rect 20871 9764 20895 9766
rect 20951 9764 20975 9766
rect 21031 9764 21037 9766
rect 20729 9755 21037 9764
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9042 19288 9454
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19260 8566 19288 8978
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18257 8188 18565 8197
rect 18257 8186 18263 8188
rect 18319 8186 18343 8188
rect 18399 8186 18423 8188
rect 18479 8186 18503 8188
rect 18559 8186 18565 8188
rect 18319 8134 18321 8186
rect 18501 8134 18503 8186
rect 18257 8132 18263 8134
rect 18319 8132 18343 8134
rect 18399 8132 18423 8134
rect 18479 8132 18503 8134
rect 18559 8132 18565 8134
rect 18257 8123 18565 8132
rect 18892 8090 18920 8434
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17788 6254 17816 6394
rect 18156 6390 18184 7890
rect 18892 7886 18920 8026
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 19352 7546 19380 8502
rect 19628 8430 19656 9522
rect 20729 8732 21037 8741
rect 20729 8730 20735 8732
rect 20791 8730 20815 8732
rect 20871 8730 20895 8732
rect 20951 8730 20975 8732
rect 21031 8730 21037 8732
rect 20791 8678 20793 8730
rect 20973 8678 20975 8730
rect 20729 8676 20735 8678
rect 20791 8676 20815 8678
rect 20871 8676 20895 8678
rect 20951 8676 20975 8678
rect 21031 8676 21037 8678
rect 20729 8667 21037 8676
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 7818 19656 8366
rect 19812 8090 19840 8502
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19890 7848 19946 7857
rect 19616 7812 19668 7818
rect 19890 7783 19946 7792
rect 19616 7754 19668 7760
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 18257 7100 18565 7109
rect 18257 7098 18263 7100
rect 18319 7098 18343 7100
rect 18399 7098 18423 7100
rect 18479 7098 18503 7100
rect 18559 7098 18565 7100
rect 18319 7046 18321 7098
rect 18501 7046 18503 7098
rect 18257 7044 18263 7046
rect 18319 7044 18343 7046
rect 18399 7044 18423 7046
rect 18479 7044 18503 7046
rect 18559 7044 18565 7046
rect 18257 7035 18565 7044
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17972 5778 18000 6122
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 5114 17908 5646
rect 17972 5234 18000 5714
rect 18064 5710 18092 6054
rect 18257 6012 18565 6021
rect 18257 6010 18263 6012
rect 18319 6010 18343 6012
rect 18399 6010 18423 6012
rect 18479 6010 18503 6012
rect 18559 6010 18565 6012
rect 18319 5958 18321 6010
rect 18501 5958 18503 6010
rect 18257 5956 18263 5958
rect 18319 5956 18343 5958
rect 18399 5956 18423 5958
rect 18479 5956 18503 5958
rect 18559 5956 18565 5958
rect 18257 5947 18565 5956
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 18064 5166 18092 5646
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18156 5302 18184 5578
rect 19628 5370 19656 7754
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18052 5160 18104 5166
rect 17880 5098 18000 5114
rect 18052 5102 18104 5108
rect 17880 5092 18012 5098
rect 17880 5086 17960 5092
rect 17960 5034 18012 5040
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 18257 4924 18565 4933
rect 18257 4922 18263 4924
rect 18319 4922 18343 4924
rect 18399 4922 18423 4924
rect 18479 4922 18503 4924
rect 18559 4922 18565 4924
rect 18319 4870 18321 4922
rect 18501 4870 18503 4922
rect 18257 4868 18263 4870
rect 18319 4868 18343 4870
rect 18399 4868 18423 4870
rect 18479 4868 18503 4870
rect 18559 4868 18565 4870
rect 18257 4859 18565 4868
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 10839 4380 11147 4389
rect 10839 4378 10845 4380
rect 10901 4378 10925 4380
rect 10981 4378 11005 4380
rect 11061 4378 11085 4380
rect 11141 4378 11147 4380
rect 10901 4326 10903 4378
rect 11083 4326 11085 4378
rect 10839 4324 10845 4326
rect 10901 4324 10925 4326
rect 10981 4324 11005 4326
rect 11061 4324 11085 4326
rect 11141 4324 11147 4326
rect 10839 4315 11147 4324
rect 15784 4380 16092 4389
rect 15784 4378 15790 4380
rect 15846 4378 15870 4380
rect 15926 4378 15950 4380
rect 16006 4378 16030 4380
rect 16086 4378 16092 4380
rect 15846 4326 15848 4378
rect 16028 4326 16030 4378
rect 15784 4324 15790 4326
rect 15846 4324 15870 4326
rect 15926 4324 15950 4326
rect 16006 4324 16030 4326
rect 16086 4324 16092 4326
rect 15784 4315 16092 4324
rect 13312 3836 13620 3845
rect 13312 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13558 3836
rect 13614 3834 13620 3836
rect 13374 3782 13376 3834
rect 13556 3782 13558 3834
rect 13312 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13558 3782
rect 13614 3780 13620 3782
rect 13312 3771 13620 3780
rect 18257 3836 18565 3845
rect 18257 3834 18263 3836
rect 18319 3834 18343 3836
rect 18399 3834 18423 3836
rect 18479 3834 18503 3836
rect 18559 3834 18565 3836
rect 18319 3782 18321 3834
rect 18501 3782 18503 3834
rect 18257 3780 18263 3782
rect 18319 3780 18343 3782
rect 18399 3780 18423 3782
rect 18479 3780 18503 3782
rect 18559 3780 18565 3782
rect 18257 3771 18565 3780
rect 10839 3292 11147 3301
rect 10839 3290 10845 3292
rect 10901 3290 10925 3292
rect 10981 3290 11005 3292
rect 11061 3290 11085 3292
rect 11141 3290 11147 3292
rect 10901 3238 10903 3290
rect 11083 3238 11085 3290
rect 10839 3236 10845 3238
rect 10901 3236 10925 3238
rect 10981 3236 11005 3238
rect 11061 3236 11085 3238
rect 11141 3236 11147 3238
rect 10839 3227 11147 3236
rect 15784 3292 16092 3301
rect 15784 3290 15790 3292
rect 15846 3290 15870 3292
rect 15926 3290 15950 3292
rect 16006 3290 16030 3292
rect 16086 3290 16092 3292
rect 15846 3238 15848 3290
rect 16028 3238 16030 3290
rect 15784 3236 15790 3238
rect 15846 3236 15870 3238
rect 15926 3236 15950 3238
rect 16006 3236 16030 3238
rect 16086 3236 16092 3238
rect 15784 3227 16092 3236
rect 13312 2748 13620 2757
rect 13312 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13558 2748
rect 13614 2746 13620 2748
rect 13374 2694 13376 2746
rect 13556 2694 13558 2746
rect 13312 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13558 2694
rect 13614 2692 13620 2694
rect 13312 2683 13620 2692
rect 18257 2748 18565 2757
rect 18257 2746 18263 2748
rect 18319 2746 18343 2748
rect 18399 2746 18423 2748
rect 18479 2746 18503 2748
rect 18559 2746 18565 2748
rect 18319 2694 18321 2746
rect 18501 2694 18503 2746
rect 18257 2692 18263 2694
rect 18319 2692 18343 2694
rect 18399 2692 18423 2694
rect 18479 2692 18503 2694
rect 18559 2692 18565 2694
rect 18257 2683 18565 2692
rect 19904 2446 19932 7783
rect 20729 7644 21037 7653
rect 20729 7642 20735 7644
rect 20791 7642 20815 7644
rect 20871 7642 20895 7644
rect 20951 7642 20975 7644
rect 21031 7642 21037 7644
rect 20791 7590 20793 7642
rect 20973 7590 20975 7642
rect 20729 7588 20735 7590
rect 20791 7588 20815 7590
rect 20871 7588 20895 7590
rect 20951 7588 20975 7590
rect 21031 7588 21037 7590
rect 20729 7579 21037 7588
rect 20729 6556 21037 6565
rect 20729 6554 20735 6556
rect 20791 6554 20815 6556
rect 20871 6554 20895 6556
rect 20951 6554 20975 6556
rect 21031 6554 21037 6556
rect 20791 6502 20793 6554
rect 20973 6502 20975 6554
rect 20729 6500 20735 6502
rect 20791 6500 20815 6502
rect 20871 6500 20895 6502
rect 20951 6500 20975 6502
rect 21031 6500 21037 6502
rect 20729 6491 21037 6500
rect 20729 5468 21037 5477
rect 20729 5466 20735 5468
rect 20791 5466 20815 5468
rect 20871 5466 20895 5468
rect 20951 5466 20975 5468
rect 21031 5466 21037 5468
rect 20791 5414 20793 5466
rect 20973 5414 20975 5466
rect 20729 5412 20735 5414
rect 20791 5412 20815 5414
rect 20871 5412 20895 5414
rect 20951 5412 20975 5414
rect 21031 5412 21037 5414
rect 20729 5403 21037 5412
rect 20729 4380 21037 4389
rect 20729 4378 20735 4380
rect 20791 4378 20815 4380
rect 20871 4378 20895 4380
rect 20951 4378 20975 4380
rect 21031 4378 21037 4380
rect 20791 4326 20793 4378
rect 20973 4326 20975 4378
rect 20729 4324 20735 4326
rect 20791 4324 20815 4326
rect 20871 4324 20895 4326
rect 20951 4324 20975 4326
rect 21031 4324 21037 4326
rect 20729 4315 21037 4324
rect 20729 3292 21037 3301
rect 20729 3290 20735 3292
rect 20791 3290 20815 3292
rect 20871 3290 20895 3292
rect 20951 3290 20975 3292
rect 21031 3290 21037 3292
rect 20791 3238 20793 3290
rect 20973 3238 20975 3290
rect 20729 3236 20735 3238
rect 20791 3236 20815 3238
rect 20871 3236 20895 3238
rect 20951 3236 20975 3238
rect 21031 3236 21037 3238
rect 20729 3227 21037 3236
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9692 898 9720 2246
rect 10839 2204 11147 2213
rect 10839 2202 10845 2204
rect 10901 2202 10925 2204
rect 10981 2202 11005 2204
rect 11061 2202 11085 2204
rect 11141 2202 11147 2204
rect 10901 2150 10903 2202
rect 11083 2150 11085 2202
rect 10839 2148 10845 2150
rect 10901 2148 10925 2150
rect 10981 2148 11005 2150
rect 11061 2148 11085 2150
rect 11141 2148 11147 2150
rect 10839 2139 11147 2148
rect 12452 898 12480 2314
rect 15212 898 15240 2314
rect 15784 2204 16092 2213
rect 15784 2202 15790 2204
rect 15846 2202 15870 2204
rect 15926 2202 15950 2204
rect 16006 2202 16030 2204
rect 16086 2202 16092 2204
rect 15846 2150 15848 2202
rect 16028 2150 16030 2202
rect 15784 2148 15790 2150
rect 15846 2148 15870 2150
rect 15926 2148 15950 2150
rect 16006 2148 16030 2150
rect 16086 2148 16092 2150
rect 15784 2139 16092 2148
rect 17972 898 18000 2314
rect 9600 870 9720 898
rect 12268 870 12480 898
rect 14936 870 15240 898
rect 17604 870 18000 898
rect 9600 800 9628 870
rect 12268 800 12296 870
rect 14936 800 14964 870
rect 17604 800 17632 870
rect 20272 800 20300 2314
rect 20729 2204 21037 2213
rect 20729 2202 20735 2204
rect 20791 2202 20815 2204
rect 20871 2202 20895 2204
rect 20951 2202 20975 2204
rect 21031 2202 21037 2204
rect 20791 2150 20793 2202
rect 20973 2150 20975 2202
rect 20729 2148 20735 2150
rect 20791 2148 20815 2150
rect 20871 2148 20895 2150
rect 20951 2148 20975 2150
rect 21031 2148 21037 2150
rect 20729 2139 21037 2148
rect 1582 0 1638 800
rect 4250 0 4306 800
rect 6918 0 6974 800
rect 9586 0 9642 800
rect 12254 0 12310 800
rect 14922 0 14978 800
rect 17590 0 17646 800
rect 20258 0 20314 800
<< via2 >>
rect 3428 19066 3484 19068
rect 3508 19066 3564 19068
rect 3588 19066 3644 19068
rect 3668 19066 3724 19068
rect 3428 19014 3474 19066
rect 3474 19014 3484 19066
rect 3508 19014 3538 19066
rect 3538 19014 3550 19066
rect 3550 19014 3564 19066
rect 3588 19014 3602 19066
rect 3602 19014 3614 19066
rect 3614 19014 3644 19066
rect 3668 19014 3678 19066
rect 3678 19014 3724 19066
rect 3428 19012 3484 19014
rect 3508 19012 3564 19014
rect 3588 19012 3644 19014
rect 3668 19012 3724 19014
rect 3428 17978 3484 17980
rect 3508 17978 3564 17980
rect 3588 17978 3644 17980
rect 3668 17978 3724 17980
rect 3428 17926 3474 17978
rect 3474 17926 3484 17978
rect 3508 17926 3538 17978
rect 3538 17926 3550 17978
rect 3550 17926 3564 17978
rect 3588 17926 3602 17978
rect 3602 17926 3614 17978
rect 3614 17926 3644 17978
rect 3668 17926 3678 17978
rect 3678 17926 3724 17978
rect 3428 17924 3484 17926
rect 3508 17924 3564 17926
rect 3588 17924 3644 17926
rect 3668 17924 3724 17926
rect 5900 19610 5956 19612
rect 5980 19610 6036 19612
rect 6060 19610 6116 19612
rect 6140 19610 6196 19612
rect 5900 19558 5946 19610
rect 5946 19558 5956 19610
rect 5980 19558 6010 19610
rect 6010 19558 6022 19610
rect 6022 19558 6036 19610
rect 6060 19558 6074 19610
rect 6074 19558 6086 19610
rect 6086 19558 6116 19610
rect 6140 19558 6150 19610
rect 6150 19558 6196 19610
rect 5900 19556 5956 19558
rect 5980 19556 6036 19558
rect 6060 19556 6116 19558
rect 6140 19556 6196 19558
rect 10845 19610 10901 19612
rect 10925 19610 10981 19612
rect 11005 19610 11061 19612
rect 11085 19610 11141 19612
rect 10845 19558 10891 19610
rect 10891 19558 10901 19610
rect 10925 19558 10955 19610
rect 10955 19558 10967 19610
rect 10967 19558 10981 19610
rect 11005 19558 11019 19610
rect 11019 19558 11031 19610
rect 11031 19558 11061 19610
rect 11085 19558 11095 19610
rect 11095 19558 11141 19610
rect 10845 19556 10901 19558
rect 10925 19556 10981 19558
rect 11005 19556 11061 19558
rect 11085 19556 11141 19558
rect 8373 19066 8429 19068
rect 8453 19066 8509 19068
rect 8533 19066 8589 19068
rect 8613 19066 8669 19068
rect 8373 19014 8419 19066
rect 8419 19014 8429 19066
rect 8453 19014 8483 19066
rect 8483 19014 8495 19066
rect 8495 19014 8509 19066
rect 8533 19014 8547 19066
rect 8547 19014 8559 19066
rect 8559 19014 8589 19066
rect 8613 19014 8623 19066
rect 8623 19014 8669 19066
rect 8373 19012 8429 19014
rect 8453 19012 8509 19014
rect 8533 19012 8589 19014
rect 8613 19012 8669 19014
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13558 19066 13614 19068
rect 13318 19014 13364 19066
rect 13364 19014 13374 19066
rect 13398 19014 13428 19066
rect 13428 19014 13440 19066
rect 13440 19014 13454 19066
rect 13478 19014 13492 19066
rect 13492 19014 13504 19066
rect 13504 19014 13534 19066
rect 13558 19014 13568 19066
rect 13568 19014 13614 19066
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13558 19012 13614 19014
rect 5900 18522 5956 18524
rect 5980 18522 6036 18524
rect 6060 18522 6116 18524
rect 6140 18522 6196 18524
rect 5900 18470 5946 18522
rect 5946 18470 5956 18522
rect 5980 18470 6010 18522
rect 6010 18470 6022 18522
rect 6022 18470 6036 18522
rect 6060 18470 6074 18522
rect 6074 18470 6086 18522
rect 6086 18470 6116 18522
rect 6140 18470 6150 18522
rect 6150 18470 6196 18522
rect 5900 18468 5956 18470
rect 5980 18468 6036 18470
rect 6060 18468 6116 18470
rect 6140 18468 6196 18470
rect 3428 16890 3484 16892
rect 3508 16890 3564 16892
rect 3588 16890 3644 16892
rect 3668 16890 3724 16892
rect 3428 16838 3474 16890
rect 3474 16838 3484 16890
rect 3508 16838 3538 16890
rect 3538 16838 3550 16890
rect 3550 16838 3564 16890
rect 3588 16838 3602 16890
rect 3602 16838 3614 16890
rect 3614 16838 3644 16890
rect 3668 16838 3678 16890
rect 3678 16838 3724 16890
rect 3428 16836 3484 16838
rect 3508 16836 3564 16838
rect 3588 16836 3644 16838
rect 3668 16836 3724 16838
rect 8373 17978 8429 17980
rect 8453 17978 8509 17980
rect 8533 17978 8589 17980
rect 8613 17978 8669 17980
rect 8373 17926 8419 17978
rect 8419 17926 8429 17978
rect 8453 17926 8483 17978
rect 8483 17926 8495 17978
rect 8495 17926 8509 17978
rect 8533 17926 8547 17978
rect 8547 17926 8559 17978
rect 8559 17926 8589 17978
rect 8613 17926 8623 17978
rect 8623 17926 8669 17978
rect 8373 17924 8429 17926
rect 8453 17924 8509 17926
rect 8533 17924 8589 17926
rect 8613 17924 8669 17926
rect 10845 18522 10901 18524
rect 10925 18522 10981 18524
rect 11005 18522 11061 18524
rect 11085 18522 11141 18524
rect 10845 18470 10891 18522
rect 10891 18470 10901 18522
rect 10925 18470 10955 18522
rect 10955 18470 10967 18522
rect 10967 18470 10981 18522
rect 11005 18470 11019 18522
rect 11019 18470 11031 18522
rect 11031 18470 11061 18522
rect 11085 18470 11095 18522
rect 11095 18470 11141 18522
rect 10845 18468 10901 18470
rect 10925 18468 10981 18470
rect 11005 18468 11061 18470
rect 11085 18468 11141 18470
rect 10966 18128 11022 18184
rect 5900 17434 5956 17436
rect 5980 17434 6036 17436
rect 6060 17434 6116 17436
rect 6140 17434 6196 17436
rect 5900 17382 5946 17434
rect 5946 17382 5956 17434
rect 5980 17382 6010 17434
rect 6010 17382 6022 17434
rect 6022 17382 6036 17434
rect 6060 17382 6074 17434
rect 6074 17382 6086 17434
rect 6086 17382 6116 17434
rect 6140 17382 6150 17434
rect 6150 17382 6196 17434
rect 5900 17380 5956 17382
rect 5980 17380 6036 17382
rect 6060 17380 6116 17382
rect 6140 17380 6196 17382
rect 5900 16346 5956 16348
rect 5980 16346 6036 16348
rect 6060 16346 6116 16348
rect 6140 16346 6196 16348
rect 5900 16294 5946 16346
rect 5946 16294 5956 16346
rect 5980 16294 6010 16346
rect 6010 16294 6022 16346
rect 6022 16294 6036 16346
rect 6060 16294 6074 16346
rect 6074 16294 6086 16346
rect 6086 16294 6116 16346
rect 6140 16294 6150 16346
rect 6150 16294 6196 16346
rect 5900 16292 5956 16294
rect 5980 16292 6036 16294
rect 6060 16292 6116 16294
rect 6140 16292 6196 16294
rect 8373 16890 8429 16892
rect 8453 16890 8509 16892
rect 8533 16890 8589 16892
rect 8613 16890 8669 16892
rect 8373 16838 8419 16890
rect 8419 16838 8429 16890
rect 8453 16838 8483 16890
rect 8483 16838 8495 16890
rect 8495 16838 8509 16890
rect 8533 16838 8547 16890
rect 8547 16838 8559 16890
rect 8559 16838 8589 16890
rect 8613 16838 8623 16890
rect 8623 16838 8669 16890
rect 8373 16836 8429 16838
rect 8453 16836 8509 16838
rect 8533 16836 8589 16838
rect 8613 16836 8669 16838
rect 3428 15802 3484 15804
rect 3508 15802 3564 15804
rect 3588 15802 3644 15804
rect 3668 15802 3724 15804
rect 3428 15750 3474 15802
rect 3474 15750 3484 15802
rect 3508 15750 3538 15802
rect 3538 15750 3550 15802
rect 3550 15750 3564 15802
rect 3588 15750 3602 15802
rect 3602 15750 3614 15802
rect 3614 15750 3644 15802
rect 3668 15750 3678 15802
rect 3678 15750 3724 15802
rect 3428 15748 3484 15750
rect 3508 15748 3564 15750
rect 3588 15748 3644 15750
rect 3668 15748 3724 15750
rect 8373 15802 8429 15804
rect 8453 15802 8509 15804
rect 8533 15802 8589 15804
rect 8613 15802 8669 15804
rect 8373 15750 8419 15802
rect 8419 15750 8429 15802
rect 8453 15750 8483 15802
rect 8483 15750 8495 15802
rect 8495 15750 8509 15802
rect 8533 15750 8547 15802
rect 8547 15750 8559 15802
rect 8559 15750 8589 15802
rect 8613 15750 8623 15802
rect 8623 15750 8669 15802
rect 8373 15748 8429 15750
rect 8453 15748 8509 15750
rect 8533 15748 8589 15750
rect 8613 15748 8669 15750
rect 3428 14714 3484 14716
rect 3508 14714 3564 14716
rect 3588 14714 3644 14716
rect 3668 14714 3724 14716
rect 3428 14662 3474 14714
rect 3474 14662 3484 14714
rect 3508 14662 3538 14714
rect 3538 14662 3550 14714
rect 3550 14662 3564 14714
rect 3588 14662 3602 14714
rect 3602 14662 3614 14714
rect 3614 14662 3644 14714
rect 3668 14662 3678 14714
rect 3678 14662 3724 14714
rect 3428 14660 3484 14662
rect 3508 14660 3564 14662
rect 3588 14660 3644 14662
rect 3668 14660 3724 14662
rect 5900 15258 5956 15260
rect 5980 15258 6036 15260
rect 6060 15258 6116 15260
rect 6140 15258 6196 15260
rect 5900 15206 5946 15258
rect 5946 15206 5956 15258
rect 5980 15206 6010 15258
rect 6010 15206 6022 15258
rect 6022 15206 6036 15258
rect 6060 15206 6074 15258
rect 6074 15206 6086 15258
rect 6086 15206 6116 15258
rect 6140 15206 6150 15258
rect 6150 15206 6196 15258
rect 5900 15204 5956 15206
rect 5980 15204 6036 15206
rect 6060 15204 6116 15206
rect 6140 15204 6196 15206
rect 3428 13626 3484 13628
rect 3508 13626 3564 13628
rect 3588 13626 3644 13628
rect 3668 13626 3724 13628
rect 3428 13574 3474 13626
rect 3474 13574 3484 13626
rect 3508 13574 3538 13626
rect 3538 13574 3550 13626
rect 3550 13574 3564 13626
rect 3588 13574 3602 13626
rect 3602 13574 3614 13626
rect 3614 13574 3644 13626
rect 3668 13574 3678 13626
rect 3678 13574 3724 13626
rect 3428 13572 3484 13574
rect 3508 13572 3564 13574
rect 3588 13572 3644 13574
rect 3668 13572 3724 13574
rect 3428 12538 3484 12540
rect 3508 12538 3564 12540
rect 3588 12538 3644 12540
rect 3668 12538 3724 12540
rect 3428 12486 3474 12538
rect 3474 12486 3484 12538
rect 3508 12486 3538 12538
rect 3538 12486 3550 12538
rect 3550 12486 3564 12538
rect 3588 12486 3602 12538
rect 3602 12486 3614 12538
rect 3614 12486 3644 12538
rect 3668 12486 3678 12538
rect 3678 12486 3724 12538
rect 3428 12484 3484 12486
rect 3508 12484 3564 12486
rect 3588 12484 3644 12486
rect 3668 12484 3724 12486
rect 5900 14170 5956 14172
rect 5980 14170 6036 14172
rect 6060 14170 6116 14172
rect 6140 14170 6196 14172
rect 5900 14118 5946 14170
rect 5946 14118 5956 14170
rect 5980 14118 6010 14170
rect 6010 14118 6022 14170
rect 6022 14118 6036 14170
rect 6060 14118 6074 14170
rect 6074 14118 6086 14170
rect 6086 14118 6116 14170
rect 6140 14118 6150 14170
rect 6150 14118 6196 14170
rect 5900 14116 5956 14118
rect 5980 14116 6036 14118
rect 6060 14116 6116 14118
rect 6140 14116 6196 14118
rect 5900 13082 5956 13084
rect 5980 13082 6036 13084
rect 6060 13082 6116 13084
rect 6140 13082 6196 13084
rect 5900 13030 5946 13082
rect 5946 13030 5956 13082
rect 5980 13030 6010 13082
rect 6010 13030 6022 13082
rect 6022 13030 6036 13082
rect 6060 13030 6074 13082
rect 6074 13030 6086 13082
rect 6086 13030 6116 13082
rect 6140 13030 6150 13082
rect 6150 13030 6196 13082
rect 5900 13028 5956 13030
rect 5980 13028 6036 13030
rect 6060 13028 6116 13030
rect 6140 13028 6196 13030
rect 5900 11994 5956 11996
rect 5980 11994 6036 11996
rect 6060 11994 6116 11996
rect 6140 11994 6196 11996
rect 5900 11942 5946 11994
rect 5946 11942 5956 11994
rect 5980 11942 6010 11994
rect 6010 11942 6022 11994
rect 6022 11942 6036 11994
rect 6060 11942 6074 11994
rect 6074 11942 6086 11994
rect 6086 11942 6116 11994
rect 6140 11942 6150 11994
rect 6150 11942 6196 11994
rect 5900 11940 5956 11942
rect 5980 11940 6036 11942
rect 6060 11940 6116 11942
rect 6140 11940 6196 11942
rect 3428 11450 3484 11452
rect 3508 11450 3564 11452
rect 3588 11450 3644 11452
rect 3668 11450 3724 11452
rect 3428 11398 3474 11450
rect 3474 11398 3484 11450
rect 3508 11398 3538 11450
rect 3538 11398 3550 11450
rect 3550 11398 3564 11450
rect 3588 11398 3602 11450
rect 3602 11398 3614 11450
rect 3614 11398 3644 11450
rect 3668 11398 3678 11450
rect 3678 11398 3724 11450
rect 3428 11396 3484 11398
rect 3508 11396 3564 11398
rect 3588 11396 3644 11398
rect 3668 11396 3724 11398
rect 5900 10906 5956 10908
rect 5980 10906 6036 10908
rect 6060 10906 6116 10908
rect 6140 10906 6196 10908
rect 5900 10854 5946 10906
rect 5946 10854 5956 10906
rect 5980 10854 6010 10906
rect 6010 10854 6022 10906
rect 6022 10854 6036 10906
rect 6060 10854 6074 10906
rect 6074 10854 6086 10906
rect 6086 10854 6116 10906
rect 6140 10854 6150 10906
rect 6150 10854 6196 10906
rect 5900 10852 5956 10854
rect 5980 10852 6036 10854
rect 6060 10852 6116 10854
rect 6140 10852 6196 10854
rect 3428 10362 3484 10364
rect 3508 10362 3564 10364
rect 3588 10362 3644 10364
rect 3668 10362 3724 10364
rect 3428 10310 3474 10362
rect 3474 10310 3484 10362
rect 3508 10310 3538 10362
rect 3538 10310 3550 10362
rect 3550 10310 3564 10362
rect 3588 10310 3602 10362
rect 3602 10310 3614 10362
rect 3614 10310 3644 10362
rect 3668 10310 3678 10362
rect 3678 10310 3724 10362
rect 3428 10308 3484 10310
rect 3508 10308 3564 10310
rect 3588 10308 3644 10310
rect 3668 10308 3724 10310
rect 3428 9274 3484 9276
rect 3508 9274 3564 9276
rect 3588 9274 3644 9276
rect 3668 9274 3724 9276
rect 3428 9222 3474 9274
rect 3474 9222 3484 9274
rect 3508 9222 3538 9274
rect 3538 9222 3550 9274
rect 3550 9222 3564 9274
rect 3588 9222 3602 9274
rect 3602 9222 3614 9274
rect 3614 9222 3644 9274
rect 3668 9222 3678 9274
rect 3678 9222 3724 9274
rect 3428 9220 3484 9222
rect 3508 9220 3564 9222
rect 3588 9220 3644 9222
rect 3668 9220 3724 9222
rect 5900 9818 5956 9820
rect 5980 9818 6036 9820
rect 6060 9818 6116 9820
rect 6140 9818 6196 9820
rect 5900 9766 5946 9818
rect 5946 9766 5956 9818
rect 5980 9766 6010 9818
rect 6010 9766 6022 9818
rect 6022 9766 6036 9818
rect 6060 9766 6074 9818
rect 6074 9766 6086 9818
rect 6086 9766 6116 9818
rect 6140 9766 6150 9818
rect 6150 9766 6196 9818
rect 5900 9764 5956 9766
rect 5980 9764 6036 9766
rect 6060 9764 6116 9766
rect 6140 9764 6196 9766
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3588 8186 3644 8188
rect 3668 8186 3724 8188
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3550 8186
rect 3550 8134 3564 8186
rect 3588 8134 3602 8186
rect 3602 8134 3614 8186
rect 3614 8134 3644 8186
rect 3668 8134 3678 8186
rect 3678 8134 3724 8186
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 3588 8132 3644 8134
rect 3668 8132 3724 8134
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3588 7098 3644 7100
rect 3668 7098 3724 7100
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3550 7098
rect 3550 7046 3564 7098
rect 3588 7046 3602 7098
rect 3602 7046 3614 7098
rect 3614 7046 3644 7098
rect 3668 7046 3678 7098
rect 3678 7046 3724 7098
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 3588 7044 3644 7046
rect 3668 7044 3724 7046
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3588 6010 3644 6012
rect 3668 6010 3724 6012
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3550 6010
rect 3550 5958 3564 6010
rect 3588 5958 3602 6010
rect 3602 5958 3614 6010
rect 3614 5958 3644 6010
rect 3668 5958 3678 6010
rect 3678 5958 3724 6010
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 3588 5956 3644 5958
rect 3668 5956 3724 5958
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3588 4922 3644 4924
rect 3668 4922 3724 4924
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3550 4922
rect 3550 4870 3564 4922
rect 3588 4870 3602 4922
rect 3602 4870 3614 4922
rect 3614 4870 3644 4922
rect 3668 4870 3678 4922
rect 3678 4870 3724 4922
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3588 4868 3644 4870
rect 3668 4868 3724 4870
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3588 3834 3644 3836
rect 3668 3834 3724 3836
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3550 3834
rect 3550 3782 3564 3834
rect 3588 3782 3602 3834
rect 3602 3782 3614 3834
rect 3614 3782 3644 3834
rect 3668 3782 3678 3834
rect 3678 3782 3724 3834
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3588 3780 3644 3782
rect 3668 3780 3724 3782
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3588 2746 3644 2748
rect 3668 2746 3724 2748
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3550 2746
rect 3550 2694 3564 2746
rect 3588 2694 3602 2746
rect 3602 2694 3614 2746
rect 3614 2694 3644 2746
rect 3668 2694 3678 2746
rect 3678 2694 3724 2746
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 3588 2692 3644 2694
rect 3668 2692 3724 2694
rect 5900 8730 5956 8732
rect 5980 8730 6036 8732
rect 6060 8730 6116 8732
rect 6140 8730 6196 8732
rect 5900 8678 5946 8730
rect 5946 8678 5956 8730
rect 5980 8678 6010 8730
rect 6010 8678 6022 8730
rect 6022 8678 6036 8730
rect 6060 8678 6074 8730
rect 6074 8678 6086 8730
rect 6086 8678 6116 8730
rect 6140 8678 6150 8730
rect 6150 8678 6196 8730
rect 5900 8676 5956 8678
rect 5980 8676 6036 8678
rect 6060 8676 6116 8678
rect 6140 8676 6196 8678
rect 5900 7642 5956 7644
rect 5980 7642 6036 7644
rect 6060 7642 6116 7644
rect 6140 7642 6196 7644
rect 5900 7590 5946 7642
rect 5946 7590 5956 7642
rect 5980 7590 6010 7642
rect 6010 7590 6022 7642
rect 6022 7590 6036 7642
rect 6060 7590 6074 7642
rect 6074 7590 6086 7642
rect 6086 7590 6116 7642
rect 6140 7590 6150 7642
rect 6150 7590 6196 7642
rect 5900 7588 5956 7590
rect 5980 7588 6036 7590
rect 6060 7588 6116 7590
rect 6140 7588 6196 7590
rect 5900 6554 5956 6556
rect 5980 6554 6036 6556
rect 6060 6554 6116 6556
rect 6140 6554 6196 6556
rect 5900 6502 5946 6554
rect 5946 6502 5956 6554
rect 5980 6502 6010 6554
rect 6010 6502 6022 6554
rect 6022 6502 6036 6554
rect 6060 6502 6074 6554
rect 6074 6502 6086 6554
rect 6086 6502 6116 6554
rect 6140 6502 6150 6554
rect 6150 6502 6196 6554
rect 5900 6500 5956 6502
rect 5980 6500 6036 6502
rect 6060 6500 6116 6502
rect 6140 6500 6196 6502
rect 5900 5466 5956 5468
rect 5980 5466 6036 5468
rect 6060 5466 6116 5468
rect 6140 5466 6196 5468
rect 5900 5414 5946 5466
rect 5946 5414 5956 5466
rect 5980 5414 6010 5466
rect 6010 5414 6022 5466
rect 6022 5414 6036 5466
rect 6060 5414 6074 5466
rect 6074 5414 6086 5466
rect 6086 5414 6116 5466
rect 6140 5414 6150 5466
rect 6150 5414 6196 5466
rect 5900 5412 5956 5414
rect 5980 5412 6036 5414
rect 6060 5412 6116 5414
rect 6140 5412 6196 5414
rect 5900 4378 5956 4380
rect 5980 4378 6036 4380
rect 6060 4378 6116 4380
rect 6140 4378 6196 4380
rect 5900 4326 5946 4378
rect 5946 4326 5956 4378
rect 5980 4326 6010 4378
rect 6010 4326 6022 4378
rect 6022 4326 6036 4378
rect 6060 4326 6074 4378
rect 6074 4326 6086 4378
rect 6086 4326 6116 4378
rect 6140 4326 6150 4378
rect 6150 4326 6196 4378
rect 5900 4324 5956 4326
rect 5980 4324 6036 4326
rect 6060 4324 6116 4326
rect 6140 4324 6196 4326
rect 5900 3290 5956 3292
rect 5980 3290 6036 3292
rect 6060 3290 6116 3292
rect 6140 3290 6196 3292
rect 5900 3238 5946 3290
rect 5946 3238 5956 3290
rect 5980 3238 6010 3290
rect 6010 3238 6022 3290
rect 6022 3238 6036 3290
rect 6060 3238 6074 3290
rect 6074 3238 6086 3290
rect 6086 3238 6116 3290
rect 6140 3238 6150 3290
rect 6150 3238 6196 3290
rect 5900 3236 5956 3238
rect 5980 3236 6036 3238
rect 6060 3236 6116 3238
rect 6140 3236 6196 3238
rect 10845 17434 10901 17436
rect 10925 17434 10981 17436
rect 11005 17434 11061 17436
rect 11085 17434 11141 17436
rect 10845 17382 10891 17434
rect 10891 17382 10901 17434
rect 10925 17382 10955 17434
rect 10955 17382 10967 17434
rect 10967 17382 10981 17434
rect 11005 17382 11019 17434
rect 11019 17382 11031 17434
rect 11031 17382 11061 17434
rect 11085 17382 11095 17434
rect 11095 17382 11141 17434
rect 10845 17380 10901 17382
rect 10925 17380 10981 17382
rect 11005 17380 11061 17382
rect 11085 17380 11141 17382
rect 10845 16346 10901 16348
rect 10925 16346 10981 16348
rect 11005 16346 11061 16348
rect 11085 16346 11141 16348
rect 10845 16294 10891 16346
rect 10891 16294 10901 16346
rect 10925 16294 10955 16346
rect 10955 16294 10967 16346
rect 10967 16294 10981 16346
rect 11005 16294 11019 16346
rect 11019 16294 11031 16346
rect 11031 16294 11061 16346
rect 11085 16294 11095 16346
rect 11095 16294 11141 16346
rect 10845 16292 10901 16294
rect 10925 16292 10981 16294
rect 11005 16292 11061 16294
rect 11085 16292 11141 16294
rect 9586 16124 9588 16144
rect 9588 16124 9640 16144
rect 9640 16124 9642 16144
rect 9586 16088 9642 16124
rect 10845 15258 10901 15260
rect 10925 15258 10981 15260
rect 11005 15258 11061 15260
rect 11085 15258 11141 15260
rect 10845 15206 10891 15258
rect 10891 15206 10901 15258
rect 10925 15206 10955 15258
rect 10955 15206 10967 15258
rect 10967 15206 10981 15258
rect 11005 15206 11019 15258
rect 11019 15206 11031 15258
rect 11031 15206 11061 15258
rect 11085 15206 11095 15258
rect 11095 15206 11141 15258
rect 10845 15204 10901 15206
rect 10925 15204 10981 15206
rect 11005 15204 11061 15206
rect 11085 15204 11141 15206
rect 8373 14714 8429 14716
rect 8453 14714 8509 14716
rect 8533 14714 8589 14716
rect 8613 14714 8669 14716
rect 8373 14662 8419 14714
rect 8419 14662 8429 14714
rect 8453 14662 8483 14714
rect 8483 14662 8495 14714
rect 8495 14662 8509 14714
rect 8533 14662 8547 14714
rect 8547 14662 8559 14714
rect 8559 14662 8589 14714
rect 8613 14662 8623 14714
rect 8623 14662 8669 14714
rect 8373 14660 8429 14662
rect 8453 14660 8509 14662
rect 8533 14660 8589 14662
rect 8613 14660 8669 14662
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13558 17978 13614 17980
rect 13318 17926 13364 17978
rect 13364 17926 13374 17978
rect 13398 17926 13428 17978
rect 13428 17926 13440 17978
rect 13440 17926 13454 17978
rect 13478 17926 13492 17978
rect 13492 17926 13504 17978
rect 13504 17926 13534 17978
rect 13558 17926 13568 17978
rect 13568 17926 13614 17978
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 13558 17924 13614 17926
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13558 16890 13614 16892
rect 13318 16838 13364 16890
rect 13364 16838 13374 16890
rect 13398 16838 13428 16890
rect 13428 16838 13440 16890
rect 13440 16838 13454 16890
rect 13478 16838 13492 16890
rect 13492 16838 13504 16890
rect 13504 16838 13534 16890
rect 13558 16838 13568 16890
rect 13568 16838 13614 16890
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13558 16836 13614 16838
rect 10845 14170 10901 14172
rect 10925 14170 10981 14172
rect 11005 14170 11061 14172
rect 11085 14170 11141 14172
rect 10845 14118 10891 14170
rect 10891 14118 10901 14170
rect 10925 14118 10955 14170
rect 10955 14118 10967 14170
rect 10967 14118 10981 14170
rect 11005 14118 11019 14170
rect 11019 14118 11031 14170
rect 11031 14118 11061 14170
rect 11085 14118 11095 14170
rect 11095 14118 11141 14170
rect 10845 14116 10901 14118
rect 10925 14116 10981 14118
rect 11005 14116 11061 14118
rect 11085 14116 11141 14118
rect 8373 13626 8429 13628
rect 8453 13626 8509 13628
rect 8533 13626 8589 13628
rect 8613 13626 8669 13628
rect 8373 13574 8419 13626
rect 8419 13574 8429 13626
rect 8453 13574 8483 13626
rect 8483 13574 8495 13626
rect 8495 13574 8509 13626
rect 8533 13574 8547 13626
rect 8547 13574 8559 13626
rect 8559 13574 8589 13626
rect 8613 13574 8623 13626
rect 8623 13574 8669 13626
rect 8373 13572 8429 13574
rect 8453 13572 8509 13574
rect 8533 13572 8589 13574
rect 8613 13572 8669 13574
rect 8373 12538 8429 12540
rect 8453 12538 8509 12540
rect 8533 12538 8589 12540
rect 8613 12538 8669 12540
rect 8373 12486 8419 12538
rect 8419 12486 8429 12538
rect 8453 12486 8483 12538
rect 8483 12486 8495 12538
rect 8495 12486 8509 12538
rect 8533 12486 8547 12538
rect 8547 12486 8559 12538
rect 8559 12486 8589 12538
rect 8613 12486 8623 12538
rect 8623 12486 8669 12538
rect 8373 12484 8429 12486
rect 8453 12484 8509 12486
rect 8533 12484 8589 12486
rect 8613 12484 8669 12486
rect 8373 11450 8429 11452
rect 8453 11450 8509 11452
rect 8533 11450 8589 11452
rect 8613 11450 8669 11452
rect 8373 11398 8419 11450
rect 8419 11398 8429 11450
rect 8453 11398 8483 11450
rect 8483 11398 8495 11450
rect 8495 11398 8509 11450
rect 8533 11398 8547 11450
rect 8547 11398 8559 11450
rect 8559 11398 8589 11450
rect 8613 11398 8623 11450
rect 8623 11398 8669 11450
rect 8373 11396 8429 11398
rect 8453 11396 8509 11398
rect 8533 11396 8589 11398
rect 8613 11396 8669 11398
rect 8373 10362 8429 10364
rect 8453 10362 8509 10364
rect 8533 10362 8589 10364
rect 8613 10362 8669 10364
rect 8373 10310 8419 10362
rect 8419 10310 8429 10362
rect 8453 10310 8483 10362
rect 8483 10310 8495 10362
rect 8495 10310 8509 10362
rect 8533 10310 8547 10362
rect 8547 10310 8559 10362
rect 8559 10310 8589 10362
rect 8613 10310 8623 10362
rect 8623 10310 8669 10362
rect 8373 10308 8429 10310
rect 8453 10308 8509 10310
rect 8533 10308 8589 10310
rect 8613 10308 8669 10310
rect 8373 9274 8429 9276
rect 8453 9274 8509 9276
rect 8533 9274 8589 9276
rect 8613 9274 8669 9276
rect 8373 9222 8419 9274
rect 8419 9222 8429 9274
rect 8453 9222 8483 9274
rect 8483 9222 8495 9274
rect 8495 9222 8509 9274
rect 8533 9222 8547 9274
rect 8547 9222 8559 9274
rect 8559 9222 8589 9274
rect 8613 9222 8623 9274
rect 8623 9222 8669 9274
rect 8373 9220 8429 9222
rect 8453 9220 8509 9222
rect 8533 9220 8589 9222
rect 8613 9220 8669 9222
rect 8373 8186 8429 8188
rect 8453 8186 8509 8188
rect 8533 8186 8589 8188
rect 8613 8186 8669 8188
rect 8373 8134 8419 8186
rect 8419 8134 8429 8186
rect 8453 8134 8483 8186
rect 8483 8134 8495 8186
rect 8495 8134 8509 8186
rect 8533 8134 8547 8186
rect 8547 8134 8559 8186
rect 8559 8134 8589 8186
rect 8613 8134 8623 8186
rect 8623 8134 8669 8186
rect 8373 8132 8429 8134
rect 8453 8132 8509 8134
rect 8533 8132 8589 8134
rect 8613 8132 8669 8134
rect 8373 7098 8429 7100
rect 8453 7098 8509 7100
rect 8533 7098 8589 7100
rect 8613 7098 8669 7100
rect 8373 7046 8419 7098
rect 8419 7046 8429 7098
rect 8453 7046 8483 7098
rect 8483 7046 8495 7098
rect 8495 7046 8509 7098
rect 8533 7046 8547 7098
rect 8547 7046 8559 7098
rect 8559 7046 8589 7098
rect 8613 7046 8623 7098
rect 8623 7046 8669 7098
rect 8373 7044 8429 7046
rect 8453 7044 8509 7046
rect 8533 7044 8589 7046
rect 8613 7044 8669 7046
rect 8373 6010 8429 6012
rect 8453 6010 8509 6012
rect 8533 6010 8589 6012
rect 8613 6010 8669 6012
rect 8373 5958 8419 6010
rect 8419 5958 8429 6010
rect 8453 5958 8483 6010
rect 8483 5958 8495 6010
rect 8495 5958 8509 6010
rect 8533 5958 8547 6010
rect 8547 5958 8559 6010
rect 8559 5958 8589 6010
rect 8613 5958 8623 6010
rect 8623 5958 8669 6010
rect 8373 5956 8429 5958
rect 8453 5956 8509 5958
rect 8533 5956 8589 5958
rect 8613 5956 8669 5958
rect 8373 4922 8429 4924
rect 8453 4922 8509 4924
rect 8533 4922 8589 4924
rect 8613 4922 8669 4924
rect 8373 4870 8419 4922
rect 8419 4870 8429 4922
rect 8453 4870 8483 4922
rect 8483 4870 8495 4922
rect 8495 4870 8509 4922
rect 8533 4870 8547 4922
rect 8547 4870 8559 4922
rect 8559 4870 8589 4922
rect 8613 4870 8623 4922
rect 8623 4870 8669 4922
rect 8373 4868 8429 4870
rect 8453 4868 8509 4870
rect 8533 4868 8589 4870
rect 8613 4868 8669 4870
rect 8373 3834 8429 3836
rect 8453 3834 8509 3836
rect 8533 3834 8589 3836
rect 8613 3834 8669 3836
rect 8373 3782 8419 3834
rect 8419 3782 8429 3834
rect 8453 3782 8483 3834
rect 8483 3782 8495 3834
rect 8495 3782 8509 3834
rect 8533 3782 8547 3834
rect 8547 3782 8559 3834
rect 8559 3782 8589 3834
rect 8613 3782 8623 3834
rect 8623 3782 8669 3834
rect 8373 3780 8429 3782
rect 8453 3780 8509 3782
rect 8533 3780 8589 3782
rect 8613 3780 8669 3782
rect 8373 2746 8429 2748
rect 8453 2746 8509 2748
rect 8533 2746 8589 2748
rect 8613 2746 8669 2748
rect 8373 2694 8419 2746
rect 8419 2694 8429 2746
rect 8453 2694 8483 2746
rect 8483 2694 8495 2746
rect 8495 2694 8509 2746
rect 8533 2694 8547 2746
rect 8547 2694 8559 2746
rect 8559 2694 8589 2746
rect 8613 2694 8623 2746
rect 8623 2694 8669 2746
rect 8373 2692 8429 2694
rect 8453 2692 8509 2694
rect 8533 2692 8589 2694
rect 8613 2692 8669 2694
rect 5900 2202 5956 2204
rect 5980 2202 6036 2204
rect 6060 2202 6116 2204
rect 6140 2202 6196 2204
rect 5900 2150 5946 2202
rect 5946 2150 5956 2202
rect 5980 2150 6010 2202
rect 6010 2150 6022 2202
rect 6022 2150 6036 2202
rect 6060 2150 6074 2202
rect 6074 2150 6086 2202
rect 6086 2150 6116 2202
rect 6140 2150 6150 2202
rect 6150 2150 6196 2202
rect 5900 2148 5956 2150
rect 5980 2148 6036 2150
rect 6060 2148 6116 2150
rect 6140 2148 6196 2150
rect 10845 13082 10901 13084
rect 10925 13082 10981 13084
rect 11005 13082 11061 13084
rect 11085 13082 11141 13084
rect 10845 13030 10891 13082
rect 10891 13030 10901 13082
rect 10925 13030 10955 13082
rect 10955 13030 10967 13082
rect 10967 13030 10981 13082
rect 11005 13030 11019 13082
rect 11019 13030 11031 13082
rect 11031 13030 11061 13082
rect 11085 13030 11095 13082
rect 11095 13030 11141 13082
rect 10845 13028 10901 13030
rect 10925 13028 10981 13030
rect 11005 13028 11061 13030
rect 11085 13028 11141 13030
rect 10845 11994 10901 11996
rect 10925 11994 10981 11996
rect 11005 11994 11061 11996
rect 11085 11994 11141 11996
rect 10845 11942 10891 11994
rect 10891 11942 10901 11994
rect 10925 11942 10955 11994
rect 10955 11942 10967 11994
rect 10967 11942 10981 11994
rect 11005 11942 11019 11994
rect 11019 11942 11031 11994
rect 11031 11942 11061 11994
rect 11085 11942 11095 11994
rect 11095 11942 11141 11994
rect 10845 11940 10901 11942
rect 10925 11940 10981 11942
rect 11005 11940 11061 11942
rect 11085 11940 11141 11942
rect 10845 10906 10901 10908
rect 10925 10906 10981 10908
rect 11005 10906 11061 10908
rect 11085 10906 11141 10908
rect 10845 10854 10891 10906
rect 10891 10854 10901 10906
rect 10925 10854 10955 10906
rect 10955 10854 10967 10906
rect 10967 10854 10981 10906
rect 11005 10854 11019 10906
rect 11019 10854 11031 10906
rect 11031 10854 11061 10906
rect 11085 10854 11095 10906
rect 11095 10854 11141 10906
rect 10845 10852 10901 10854
rect 10925 10852 10981 10854
rect 11005 10852 11061 10854
rect 11085 10852 11141 10854
rect 10845 9818 10901 9820
rect 10925 9818 10981 9820
rect 11005 9818 11061 9820
rect 11085 9818 11141 9820
rect 10845 9766 10891 9818
rect 10891 9766 10901 9818
rect 10925 9766 10955 9818
rect 10955 9766 10967 9818
rect 10967 9766 10981 9818
rect 11005 9766 11019 9818
rect 11019 9766 11031 9818
rect 11031 9766 11061 9818
rect 11085 9766 11095 9818
rect 11095 9766 11141 9818
rect 10845 9764 10901 9766
rect 10925 9764 10981 9766
rect 11005 9764 11061 9766
rect 11085 9764 11141 9766
rect 10845 8730 10901 8732
rect 10925 8730 10981 8732
rect 11005 8730 11061 8732
rect 11085 8730 11141 8732
rect 10845 8678 10891 8730
rect 10891 8678 10901 8730
rect 10925 8678 10955 8730
rect 10955 8678 10967 8730
rect 10967 8678 10981 8730
rect 11005 8678 11019 8730
rect 11019 8678 11031 8730
rect 11031 8678 11061 8730
rect 11085 8678 11095 8730
rect 11095 8678 11141 8730
rect 10845 8676 10901 8678
rect 10925 8676 10981 8678
rect 11005 8676 11061 8678
rect 11085 8676 11141 8678
rect 11058 7828 11060 7848
rect 11060 7828 11112 7848
rect 11112 7828 11114 7848
rect 11058 7792 11114 7828
rect 11426 7792 11482 7848
rect 10845 7642 10901 7644
rect 10925 7642 10981 7644
rect 11005 7642 11061 7644
rect 11085 7642 11141 7644
rect 10845 7590 10891 7642
rect 10891 7590 10901 7642
rect 10925 7590 10955 7642
rect 10955 7590 10967 7642
rect 10967 7590 10981 7642
rect 11005 7590 11019 7642
rect 11019 7590 11031 7642
rect 11031 7590 11061 7642
rect 11085 7590 11095 7642
rect 11095 7590 11141 7642
rect 10845 7588 10901 7590
rect 10925 7588 10981 7590
rect 11005 7588 11061 7590
rect 11085 7588 11141 7590
rect 10845 6554 10901 6556
rect 10925 6554 10981 6556
rect 11005 6554 11061 6556
rect 11085 6554 11141 6556
rect 10845 6502 10891 6554
rect 10891 6502 10901 6554
rect 10925 6502 10955 6554
rect 10955 6502 10967 6554
rect 10967 6502 10981 6554
rect 11005 6502 11019 6554
rect 11019 6502 11031 6554
rect 11031 6502 11061 6554
rect 11085 6502 11095 6554
rect 11095 6502 11141 6554
rect 10845 6500 10901 6502
rect 10925 6500 10981 6502
rect 11005 6500 11061 6502
rect 11085 6500 11141 6502
rect 10845 5466 10901 5468
rect 10925 5466 10981 5468
rect 11005 5466 11061 5468
rect 11085 5466 11141 5468
rect 10845 5414 10891 5466
rect 10891 5414 10901 5466
rect 10925 5414 10955 5466
rect 10955 5414 10967 5466
rect 10967 5414 10981 5466
rect 11005 5414 11019 5466
rect 11019 5414 11031 5466
rect 11031 5414 11061 5466
rect 11085 5414 11095 5466
rect 11095 5414 11141 5466
rect 10845 5412 10901 5414
rect 10925 5412 10981 5414
rect 11005 5412 11061 5414
rect 11085 5412 11141 5414
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13558 15802 13614 15804
rect 13318 15750 13364 15802
rect 13364 15750 13374 15802
rect 13398 15750 13428 15802
rect 13428 15750 13440 15802
rect 13440 15750 13454 15802
rect 13478 15750 13492 15802
rect 13492 15750 13504 15802
rect 13504 15750 13534 15802
rect 13558 15750 13568 15802
rect 13568 15750 13614 15802
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13558 15748 13614 15750
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13558 14714 13614 14716
rect 13318 14662 13364 14714
rect 13364 14662 13374 14714
rect 13398 14662 13428 14714
rect 13428 14662 13440 14714
rect 13440 14662 13454 14714
rect 13478 14662 13492 14714
rect 13492 14662 13504 14714
rect 13504 14662 13534 14714
rect 13558 14662 13568 14714
rect 13568 14662 13614 14714
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 13558 14660 13614 14662
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13558 13626 13614 13628
rect 13318 13574 13364 13626
rect 13364 13574 13374 13626
rect 13398 13574 13428 13626
rect 13428 13574 13440 13626
rect 13440 13574 13454 13626
rect 13478 13574 13492 13626
rect 13492 13574 13504 13626
rect 13504 13574 13534 13626
rect 13558 13574 13568 13626
rect 13568 13574 13614 13626
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13558 13572 13614 13574
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13558 12538 13614 12540
rect 13318 12486 13364 12538
rect 13364 12486 13374 12538
rect 13398 12486 13428 12538
rect 13428 12486 13440 12538
rect 13440 12486 13454 12538
rect 13478 12486 13492 12538
rect 13492 12486 13504 12538
rect 13504 12486 13534 12538
rect 13558 12486 13568 12538
rect 13568 12486 13614 12538
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13558 12484 13614 12486
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13558 11450 13614 11452
rect 13318 11398 13364 11450
rect 13364 11398 13374 11450
rect 13398 11398 13428 11450
rect 13428 11398 13440 11450
rect 13440 11398 13454 11450
rect 13478 11398 13492 11450
rect 13492 11398 13504 11450
rect 13504 11398 13534 11450
rect 13558 11398 13568 11450
rect 13568 11398 13614 11450
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 13558 11396 13614 11398
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13558 10362 13614 10364
rect 13318 10310 13364 10362
rect 13364 10310 13374 10362
rect 13398 10310 13428 10362
rect 13428 10310 13440 10362
rect 13440 10310 13454 10362
rect 13478 10310 13492 10362
rect 13492 10310 13504 10362
rect 13504 10310 13534 10362
rect 13558 10310 13568 10362
rect 13568 10310 13614 10362
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13558 10308 13614 10310
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13558 9274 13614 9276
rect 13318 9222 13364 9274
rect 13364 9222 13374 9274
rect 13398 9222 13428 9274
rect 13428 9222 13440 9274
rect 13440 9222 13454 9274
rect 13478 9222 13492 9274
rect 13492 9222 13504 9274
rect 13504 9222 13534 9274
rect 13558 9222 13568 9274
rect 13568 9222 13614 9274
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13558 9220 13614 9222
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13558 8186 13614 8188
rect 13318 8134 13364 8186
rect 13364 8134 13374 8186
rect 13398 8134 13428 8186
rect 13428 8134 13440 8186
rect 13440 8134 13454 8186
rect 13478 8134 13492 8186
rect 13492 8134 13504 8186
rect 13504 8134 13534 8186
rect 13558 8134 13568 8186
rect 13568 8134 13614 8186
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13558 8132 13614 8134
rect 14646 18128 14702 18184
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13558 7098 13614 7100
rect 13318 7046 13364 7098
rect 13364 7046 13374 7098
rect 13398 7046 13428 7098
rect 13428 7046 13440 7098
rect 13440 7046 13454 7098
rect 13478 7046 13492 7098
rect 13492 7046 13504 7098
rect 13504 7046 13534 7098
rect 13558 7046 13568 7098
rect 13568 7046 13614 7098
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 13558 7044 13614 7046
rect 15790 19610 15846 19612
rect 15870 19610 15926 19612
rect 15950 19610 16006 19612
rect 16030 19610 16086 19612
rect 15790 19558 15836 19610
rect 15836 19558 15846 19610
rect 15870 19558 15900 19610
rect 15900 19558 15912 19610
rect 15912 19558 15926 19610
rect 15950 19558 15964 19610
rect 15964 19558 15976 19610
rect 15976 19558 16006 19610
rect 16030 19558 16040 19610
rect 16040 19558 16086 19610
rect 15790 19556 15846 19558
rect 15870 19556 15926 19558
rect 15950 19556 16006 19558
rect 16030 19556 16086 19558
rect 20735 19610 20791 19612
rect 20815 19610 20871 19612
rect 20895 19610 20951 19612
rect 20975 19610 21031 19612
rect 20735 19558 20781 19610
rect 20781 19558 20791 19610
rect 20815 19558 20845 19610
rect 20845 19558 20857 19610
rect 20857 19558 20871 19610
rect 20895 19558 20909 19610
rect 20909 19558 20921 19610
rect 20921 19558 20951 19610
rect 20975 19558 20985 19610
rect 20985 19558 21031 19610
rect 20735 19556 20791 19558
rect 20815 19556 20871 19558
rect 20895 19556 20951 19558
rect 20975 19556 21031 19558
rect 15790 18522 15846 18524
rect 15870 18522 15926 18524
rect 15950 18522 16006 18524
rect 16030 18522 16086 18524
rect 15790 18470 15836 18522
rect 15836 18470 15846 18522
rect 15870 18470 15900 18522
rect 15900 18470 15912 18522
rect 15912 18470 15926 18522
rect 15950 18470 15964 18522
rect 15964 18470 15976 18522
rect 15976 18470 16006 18522
rect 16030 18470 16040 18522
rect 16040 18470 16086 18522
rect 15790 18468 15846 18470
rect 15870 18468 15926 18470
rect 15950 18468 16006 18470
rect 16030 18468 16086 18470
rect 15842 18128 15898 18184
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13558 6010 13614 6012
rect 13318 5958 13364 6010
rect 13364 5958 13374 6010
rect 13398 5958 13428 6010
rect 13428 5958 13440 6010
rect 13440 5958 13454 6010
rect 13478 5958 13492 6010
rect 13492 5958 13504 6010
rect 13504 5958 13534 6010
rect 13558 5958 13568 6010
rect 13568 5958 13614 6010
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 13558 5956 13614 5958
rect 15790 17434 15846 17436
rect 15870 17434 15926 17436
rect 15950 17434 16006 17436
rect 16030 17434 16086 17436
rect 15790 17382 15836 17434
rect 15836 17382 15846 17434
rect 15870 17382 15900 17434
rect 15900 17382 15912 17434
rect 15912 17382 15926 17434
rect 15950 17382 15964 17434
rect 15964 17382 15976 17434
rect 15976 17382 16006 17434
rect 16030 17382 16040 17434
rect 16040 17382 16086 17434
rect 15790 17380 15846 17382
rect 15870 17380 15926 17382
rect 15950 17380 16006 17382
rect 16030 17380 16086 17382
rect 16854 18128 16910 18184
rect 18263 19066 18319 19068
rect 18343 19066 18399 19068
rect 18423 19066 18479 19068
rect 18503 19066 18559 19068
rect 18263 19014 18309 19066
rect 18309 19014 18319 19066
rect 18343 19014 18373 19066
rect 18373 19014 18385 19066
rect 18385 19014 18399 19066
rect 18423 19014 18437 19066
rect 18437 19014 18449 19066
rect 18449 19014 18479 19066
rect 18503 19014 18513 19066
rect 18513 19014 18559 19066
rect 18263 19012 18319 19014
rect 18343 19012 18399 19014
rect 18423 19012 18479 19014
rect 18503 19012 18559 19014
rect 18263 17978 18319 17980
rect 18343 17978 18399 17980
rect 18423 17978 18479 17980
rect 18503 17978 18559 17980
rect 18263 17926 18309 17978
rect 18309 17926 18319 17978
rect 18343 17926 18373 17978
rect 18373 17926 18385 17978
rect 18385 17926 18399 17978
rect 18423 17926 18437 17978
rect 18437 17926 18449 17978
rect 18449 17926 18479 17978
rect 18503 17926 18513 17978
rect 18513 17926 18559 17978
rect 18263 17924 18319 17926
rect 18343 17924 18399 17926
rect 18423 17924 18479 17926
rect 18503 17924 18559 17926
rect 15790 16346 15846 16348
rect 15870 16346 15926 16348
rect 15950 16346 16006 16348
rect 16030 16346 16086 16348
rect 15790 16294 15836 16346
rect 15836 16294 15846 16346
rect 15870 16294 15900 16346
rect 15900 16294 15912 16346
rect 15912 16294 15926 16346
rect 15950 16294 15964 16346
rect 15964 16294 15976 16346
rect 15976 16294 16006 16346
rect 16030 16294 16040 16346
rect 16040 16294 16086 16346
rect 15790 16292 15846 16294
rect 15870 16292 15926 16294
rect 15950 16292 16006 16294
rect 16030 16292 16086 16294
rect 15790 15258 15846 15260
rect 15870 15258 15926 15260
rect 15950 15258 16006 15260
rect 16030 15258 16086 15260
rect 15790 15206 15836 15258
rect 15836 15206 15846 15258
rect 15870 15206 15900 15258
rect 15900 15206 15912 15258
rect 15912 15206 15926 15258
rect 15950 15206 15964 15258
rect 15964 15206 15976 15258
rect 15976 15206 16006 15258
rect 16030 15206 16040 15258
rect 16040 15206 16086 15258
rect 15790 15204 15846 15206
rect 15870 15204 15926 15206
rect 15950 15204 16006 15206
rect 16030 15204 16086 15206
rect 15474 11736 15530 11792
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13558 4922 13614 4924
rect 13318 4870 13364 4922
rect 13364 4870 13374 4922
rect 13398 4870 13428 4922
rect 13428 4870 13440 4922
rect 13440 4870 13454 4922
rect 13478 4870 13492 4922
rect 13492 4870 13504 4922
rect 13504 4870 13534 4922
rect 13558 4870 13568 4922
rect 13568 4870 13614 4922
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13558 4868 13614 4870
rect 15790 14170 15846 14172
rect 15870 14170 15926 14172
rect 15950 14170 16006 14172
rect 16030 14170 16086 14172
rect 15790 14118 15836 14170
rect 15836 14118 15846 14170
rect 15870 14118 15900 14170
rect 15900 14118 15912 14170
rect 15912 14118 15926 14170
rect 15950 14118 15964 14170
rect 15964 14118 15976 14170
rect 15976 14118 16006 14170
rect 16030 14118 16040 14170
rect 16040 14118 16086 14170
rect 15790 14116 15846 14118
rect 15870 14116 15926 14118
rect 15950 14116 16006 14118
rect 16030 14116 16086 14118
rect 15790 13082 15846 13084
rect 15870 13082 15926 13084
rect 15950 13082 16006 13084
rect 16030 13082 16086 13084
rect 15790 13030 15836 13082
rect 15836 13030 15846 13082
rect 15870 13030 15900 13082
rect 15900 13030 15912 13082
rect 15912 13030 15926 13082
rect 15950 13030 15964 13082
rect 15964 13030 15976 13082
rect 15976 13030 16006 13082
rect 16030 13030 16040 13082
rect 16040 13030 16086 13082
rect 15790 13028 15846 13030
rect 15870 13028 15926 13030
rect 15950 13028 16006 13030
rect 16030 13028 16086 13030
rect 15790 11994 15846 11996
rect 15870 11994 15926 11996
rect 15950 11994 16006 11996
rect 16030 11994 16086 11996
rect 15790 11942 15836 11994
rect 15836 11942 15846 11994
rect 15870 11942 15900 11994
rect 15900 11942 15912 11994
rect 15912 11942 15926 11994
rect 15950 11942 15964 11994
rect 15964 11942 15976 11994
rect 15976 11942 16006 11994
rect 16030 11942 16040 11994
rect 16040 11942 16086 11994
rect 15790 11940 15846 11942
rect 15870 11940 15926 11942
rect 15950 11940 16006 11942
rect 16030 11940 16086 11942
rect 15790 10906 15846 10908
rect 15870 10906 15926 10908
rect 15950 10906 16006 10908
rect 16030 10906 16086 10908
rect 15790 10854 15836 10906
rect 15836 10854 15846 10906
rect 15870 10854 15900 10906
rect 15900 10854 15912 10906
rect 15912 10854 15926 10906
rect 15950 10854 15964 10906
rect 15964 10854 15976 10906
rect 15976 10854 16006 10906
rect 16030 10854 16040 10906
rect 16040 10854 16086 10906
rect 15790 10852 15846 10854
rect 15870 10852 15926 10854
rect 15950 10852 16006 10854
rect 16030 10852 16086 10854
rect 15790 9818 15846 9820
rect 15870 9818 15926 9820
rect 15950 9818 16006 9820
rect 16030 9818 16086 9820
rect 15790 9766 15836 9818
rect 15836 9766 15846 9818
rect 15870 9766 15900 9818
rect 15900 9766 15912 9818
rect 15912 9766 15926 9818
rect 15950 9766 15964 9818
rect 15964 9766 15976 9818
rect 15976 9766 16006 9818
rect 16030 9766 16040 9818
rect 16040 9766 16086 9818
rect 15790 9764 15846 9766
rect 15870 9764 15926 9766
rect 15950 9764 16006 9766
rect 16030 9764 16086 9766
rect 15790 8730 15846 8732
rect 15870 8730 15926 8732
rect 15950 8730 16006 8732
rect 16030 8730 16086 8732
rect 15790 8678 15836 8730
rect 15836 8678 15846 8730
rect 15870 8678 15900 8730
rect 15900 8678 15912 8730
rect 15912 8678 15926 8730
rect 15950 8678 15964 8730
rect 15964 8678 15976 8730
rect 15976 8678 16006 8730
rect 16030 8678 16040 8730
rect 16040 8678 16086 8730
rect 15790 8676 15846 8678
rect 15870 8676 15926 8678
rect 15950 8676 16006 8678
rect 16030 8676 16086 8678
rect 15790 7642 15846 7644
rect 15870 7642 15926 7644
rect 15950 7642 16006 7644
rect 16030 7642 16086 7644
rect 15790 7590 15836 7642
rect 15836 7590 15846 7642
rect 15870 7590 15900 7642
rect 15900 7590 15912 7642
rect 15912 7590 15926 7642
rect 15950 7590 15964 7642
rect 15964 7590 15976 7642
rect 15976 7590 16006 7642
rect 16030 7590 16040 7642
rect 16040 7590 16086 7642
rect 15790 7588 15846 7590
rect 15870 7588 15926 7590
rect 15950 7588 16006 7590
rect 16030 7588 16086 7590
rect 15790 6554 15846 6556
rect 15870 6554 15926 6556
rect 15950 6554 16006 6556
rect 16030 6554 16086 6556
rect 15790 6502 15836 6554
rect 15836 6502 15846 6554
rect 15870 6502 15900 6554
rect 15900 6502 15912 6554
rect 15912 6502 15926 6554
rect 15950 6502 15964 6554
rect 15964 6502 15976 6554
rect 15976 6502 16006 6554
rect 16030 6502 16040 6554
rect 16040 6502 16086 6554
rect 15790 6500 15846 6502
rect 15870 6500 15926 6502
rect 15950 6500 16006 6502
rect 16030 6500 16086 6502
rect 15790 5466 15846 5468
rect 15870 5466 15926 5468
rect 15950 5466 16006 5468
rect 16030 5466 16086 5468
rect 15790 5414 15836 5466
rect 15836 5414 15846 5466
rect 15870 5414 15900 5466
rect 15900 5414 15912 5466
rect 15912 5414 15926 5466
rect 15950 5414 15964 5466
rect 15964 5414 15976 5466
rect 15976 5414 16006 5466
rect 16030 5414 16040 5466
rect 16040 5414 16086 5466
rect 15790 5412 15846 5414
rect 15870 5412 15926 5414
rect 15950 5412 16006 5414
rect 16030 5412 16086 5414
rect 18263 16890 18319 16892
rect 18343 16890 18399 16892
rect 18423 16890 18479 16892
rect 18503 16890 18559 16892
rect 18263 16838 18309 16890
rect 18309 16838 18319 16890
rect 18343 16838 18373 16890
rect 18373 16838 18385 16890
rect 18385 16838 18399 16890
rect 18423 16838 18437 16890
rect 18437 16838 18449 16890
rect 18449 16838 18479 16890
rect 18503 16838 18513 16890
rect 18513 16838 18559 16890
rect 18263 16836 18319 16838
rect 18343 16836 18399 16838
rect 18423 16836 18479 16838
rect 18503 16836 18559 16838
rect 20735 18522 20791 18524
rect 20815 18522 20871 18524
rect 20895 18522 20951 18524
rect 20975 18522 21031 18524
rect 20735 18470 20781 18522
rect 20781 18470 20791 18522
rect 20815 18470 20845 18522
rect 20845 18470 20857 18522
rect 20857 18470 20871 18522
rect 20895 18470 20909 18522
rect 20909 18470 20921 18522
rect 20921 18470 20951 18522
rect 20975 18470 20985 18522
rect 20985 18470 21031 18522
rect 20735 18468 20791 18470
rect 20815 18468 20871 18470
rect 20895 18468 20951 18470
rect 20975 18468 21031 18470
rect 20735 17434 20791 17436
rect 20815 17434 20871 17436
rect 20895 17434 20951 17436
rect 20975 17434 21031 17436
rect 20735 17382 20781 17434
rect 20781 17382 20791 17434
rect 20815 17382 20845 17434
rect 20845 17382 20857 17434
rect 20857 17382 20871 17434
rect 20895 17382 20909 17434
rect 20909 17382 20921 17434
rect 20921 17382 20951 17434
rect 20975 17382 20985 17434
rect 20985 17382 21031 17434
rect 20735 17380 20791 17382
rect 20815 17380 20871 17382
rect 20895 17380 20951 17382
rect 20975 17380 21031 17382
rect 18263 15802 18319 15804
rect 18343 15802 18399 15804
rect 18423 15802 18479 15804
rect 18503 15802 18559 15804
rect 18263 15750 18309 15802
rect 18309 15750 18319 15802
rect 18343 15750 18373 15802
rect 18373 15750 18385 15802
rect 18385 15750 18399 15802
rect 18423 15750 18437 15802
rect 18437 15750 18449 15802
rect 18449 15750 18479 15802
rect 18503 15750 18513 15802
rect 18513 15750 18559 15802
rect 18263 15748 18319 15750
rect 18343 15748 18399 15750
rect 18423 15748 18479 15750
rect 18503 15748 18559 15750
rect 20735 16346 20791 16348
rect 20815 16346 20871 16348
rect 20895 16346 20951 16348
rect 20975 16346 21031 16348
rect 20735 16294 20781 16346
rect 20781 16294 20791 16346
rect 20815 16294 20845 16346
rect 20845 16294 20857 16346
rect 20857 16294 20871 16346
rect 20895 16294 20909 16346
rect 20909 16294 20921 16346
rect 20921 16294 20951 16346
rect 20975 16294 20985 16346
rect 20985 16294 21031 16346
rect 20735 16292 20791 16294
rect 20815 16292 20871 16294
rect 20895 16292 20951 16294
rect 20975 16292 21031 16294
rect 20074 16088 20130 16144
rect 18263 14714 18319 14716
rect 18343 14714 18399 14716
rect 18423 14714 18479 14716
rect 18503 14714 18559 14716
rect 18263 14662 18309 14714
rect 18309 14662 18319 14714
rect 18343 14662 18373 14714
rect 18373 14662 18385 14714
rect 18385 14662 18399 14714
rect 18423 14662 18437 14714
rect 18437 14662 18449 14714
rect 18449 14662 18479 14714
rect 18503 14662 18513 14714
rect 18513 14662 18559 14714
rect 18263 14660 18319 14662
rect 18343 14660 18399 14662
rect 18423 14660 18479 14662
rect 18503 14660 18559 14662
rect 18263 13626 18319 13628
rect 18343 13626 18399 13628
rect 18423 13626 18479 13628
rect 18503 13626 18559 13628
rect 18263 13574 18309 13626
rect 18309 13574 18319 13626
rect 18343 13574 18373 13626
rect 18373 13574 18385 13626
rect 18385 13574 18399 13626
rect 18423 13574 18437 13626
rect 18437 13574 18449 13626
rect 18449 13574 18479 13626
rect 18503 13574 18513 13626
rect 18513 13574 18559 13626
rect 18263 13572 18319 13574
rect 18343 13572 18399 13574
rect 18423 13572 18479 13574
rect 18503 13572 18559 13574
rect 18263 12538 18319 12540
rect 18343 12538 18399 12540
rect 18423 12538 18479 12540
rect 18503 12538 18559 12540
rect 18263 12486 18309 12538
rect 18309 12486 18319 12538
rect 18343 12486 18373 12538
rect 18373 12486 18385 12538
rect 18385 12486 18399 12538
rect 18423 12486 18437 12538
rect 18437 12486 18449 12538
rect 18449 12486 18479 12538
rect 18503 12486 18513 12538
rect 18513 12486 18559 12538
rect 18263 12484 18319 12486
rect 18343 12484 18399 12486
rect 18423 12484 18479 12486
rect 18503 12484 18559 12486
rect 20735 15258 20791 15260
rect 20815 15258 20871 15260
rect 20895 15258 20951 15260
rect 20975 15258 21031 15260
rect 20735 15206 20781 15258
rect 20781 15206 20791 15258
rect 20815 15206 20845 15258
rect 20845 15206 20857 15258
rect 20857 15206 20871 15258
rect 20895 15206 20909 15258
rect 20909 15206 20921 15258
rect 20921 15206 20951 15258
rect 20975 15206 20985 15258
rect 20985 15206 21031 15258
rect 20735 15204 20791 15206
rect 20815 15204 20871 15206
rect 20895 15204 20951 15206
rect 20975 15204 21031 15206
rect 20735 14170 20791 14172
rect 20815 14170 20871 14172
rect 20895 14170 20951 14172
rect 20975 14170 21031 14172
rect 20735 14118 20781 14170
rect 20781 14118 20791 14170
rect 20815 14118 20845 14170
rect 20845 14118 20857 14170
rect 20857 14118 20871 14170
rect 20895 14118 20909 14170
rect 20909 14118 20921 14170
rect 20921 14118 20951 14170
rect 20975 14118 20985 14170
rect 20985 14118 21031 14170
rect 20735 14116 20791 14118
rect 20815 14116 20871 14118
rect 20895 14116 20951 14118
rect 20975 14116 21031 14118
rect 20735 13082 20791 13084
rect 20815 13082 20871 13084
rect 20895 13082 20951 13084
rect 20975 13082 21031 13084
rect 20735 13030 20781 13082
rect 20781 13030 20791 13082
rect 20815 13030 20845 13082
rect 20845 13030 20857 13082
rect 20857 13030 20871 13082
rect 20895 13030 20909 13082
rect 20909 13030 20921 13082
rect 20921 13030 20951 13082
rect 20975 13030 20985 13082
rect 20985 13030 21031 13082
rect 20735 13028 20791 13030
rect 20815 13028 20871 13030
rect 20895 13028 20951 13030
rect 20975 13028 21031 13030
rect 19246 11756 19302 11792
rect 19246 11736 19248 11756
rect 19248 11736 19300 11756
rect 19300 11736 19302 11756
rect 18263 11450 18319 11452
rect 18343 11450 18399 11452
rect 18423 11450 18479 11452
rect 18503 11450 18559 11452
rect 18263 11398 18309 11450
rect 18309 11398 18319 11450
rect 18343 11398 18373 11450
rect 18373 11398 18385 11450
rect 18385 11398 18399 11450
rect 18423 11398 18437 11450
rect 18437 11398 18449 11450
rect 18449 11398 18479 11450
rect 18503 11398 18513 11450
rect 18513 11398 18559 11450
rect 18263 11396 18319 11398
rect 18343 11396 18399 11398
rect 18423 11396 18479 11398
rect 18503 11396 18559 11398
rect 18263 10362 18319 10364
rect 18343 10362 18399 10364
rect 18423 10362 18479 10364
rect 18503 10362 18559 10364
rect 18263 10310 18309 10362
rect 18309 10310 18319 10362
rect 18343 10310 18373 10362
rect 18373 10310 18385 10362
rect 18385 10310 18399 10362
rect 18423 10310 18437 10362
rect 18437 10310 18449 10362
rect 18449 10310 18479 10362
rect 18503 10310 18513 10362
rect 18513 10310 18559 10362
rect 18263 10308 18319 10310
rect 18343 10308 18399 10310
rect 18423 10308 18479 10310
rect 18503 10308 18559 10310
rect 20735 11994 20791 11996
rect 20815 11994 20871 11996
rect 20895 11994 20951 11996
rect 20975 11994 21031 11996
rect 20735 11942 20781 11994
rect 20781 11942 20791 11994
rect 20815 11942 20845 11994
rect 20845 11942 20857 11994
rect 20857 11942 20871 11994
rect 20895 11942 20909 11994
rect 20909 11942 20921 11994
rect 20921 11942 20951 11994
rect 20975 11942 20985 11994
rect 20985 11942 21031 11994
rect 20735 11940 20791 11942
rect 20815 11940 20871 11942
rect 20895 11940 20951 11942
rect 20975 11940 21031 11942
rect 20735 10906 20791 10908
rect 20815 10906 20871 10908
rect 20895 10906 20951 10908
rect 20975 10906 21031 10908
rect 20735 10854 20781 10906
rect 20781 10854 20791 10906
rect 20815 10854 20845 10906
rect 20845 10854 20857 10906
rect 20857 10854 20871 10906
rect 20895 10854 20909 10906
rect 20909 10854 20921 10906
rect 20921 10854 20951 10906
rect 20975 10854 20985 10906
rect 20985 10854 21031 10906
rect 20735 10852 20791 10854
rect 20815 10852 20871 10854
rect 20895 10852 20951 10854
rect 20975 10852 21031 10854
rect 18263 9274 18319 9276
rect 18343 9274 18399 9276
rect 18423 9274 18479 9276
rect 18503 9274 18559 9276
rect 18263 9222 18309 9274
rect 18309 9222 18319 9274
rect 18343 9222 18373 9274
rect 18373 9222 18385 9274
rect 18385 9222 18399 9274
rect 18423 9222 18437 9274
rect 18437 9222 18449 9274
rect 18449 9222 18479 9274
rect 18503 9222 18513 9274
rect 18513 9222 18559 9274
rect 18263 9220 18319 9222
rect 18343 9220 18399 9222
rect 18423 9220 18479 9222
rect 18503 9220 18559 9222
rect 20735 9818 20791 9820
rect 20815 9818 20871 9820
rect 20895 9818 20951 9820
rect 20975 9818 21031 9820
rect 20735 9766 20781 9818
rect 20781 9766 20791 9818
rect 20815 9766 20845 9818
rect 20845 9766 20857 9818
rect 20857 9766 20871 9818
rect 20895 9766 20909 9818
rect 20909 9766 20921 9818
rect 20921 9766 20951 9818
rect 20975 9766 20985 9818
rect 20985 9766 21031 9818
rect 20735 9764 20791 9766
rect 20815 9764 20871 9766
rect 20895 9764 20951 9766
rect 20975 9764 21031 9766
rect 18263 8186 18319 8188
rect 18343 8186 18399 8188
rect 18423 8186 18479 8188
rect 18503 8186 18559 8188
rect 18263 8134 18309 8186
rect 18309 8134 18319 8186
rect 18343 8134 18373 8186
rect 18373 8134 18385 8186
rect 18385 8134 18399 8186
rect 18423 8134 18437 8186
rect 18437 8134 18449 8186
rect 18449 8134 18479 8186
rect 18503 8134 18513 8186
rect 18513 8134 18559 8186
rect 18263 8132 18319 8134
rect 18343 8132 18399 8134
rect 18423 8132 18479 8134
rect 18503 8132 18559 8134
rect 20735 8730 20791 8732
rect 20815 8730 20871 8732
rect 20895 8730 20951 8732
rect 20975 8730 21031 8732
rect 20735 8678 20781 8730
rect 20781 8678 20791 8730
rect 20815 8678 20845 8730
rect 20845 8678 20857 8730
rect 20857 8678 20871 8730
rect 20895 8678 20909 8730
rect 20909 8678 20921 8730
rect 20921 8678 20951 8730
rect 20975 8678 20985 8730
rect 20985 8678 21031 8730
rect 20735 8676 20791 8678
rect 20815 8676 20871 8678
rect 20895 8676 20951 8678
rect 20975 8676 21031 8678
rect 19890 7792 19946 7848
rect 18263 7098 18319 7100
rect 18343 7098 18399 7100
rect 18423 7098 18479 7100
rect 18503 7098 18559 7100
rect 18263 7046 18309 7098
rect 18309 7046 18319 7098
rect 18343 7046 18373 7098
rect 18373 7046 18385 7098
rect 18385 7046 18399 7098
rect 18423 7046 18437 7098
rect 18437 7046 18449 7098
rect 18449 7046 18479 7098
rect 18503 7046 18513 7098
rect 18513 7046 18559 7098
rect 18263 7044 18319 7046
rect 18343 7044 18399 7046
rect 18423 7044 18479 7046
rect 18503 7044 18559 7046
rect 18263 6010 18319 6012
rect 18343 6010 18399 6012
rect 18423 6010 18479 6012
rect 18503 6010 18559 6012
rect 18263 5958 18309 6010
rect 18309 5958 18319 6010
rect 18343 5958 18373 6010
rect 18373 5958 18385 6010
rect 18385 5958 18399 6010
rect 18423 5958 18437 6010
rect 18437 5958 18449 6010
rect 18449 5958 18479 6010
rect 18503 5958 18513 6010
rect 18513 5958 18559 6010
rect 18263 5956 18319 5958
rect 18343 5956 18399 5958
rect 18423 5956 18479 5958
rect 18503 5956 18559 5958
rect 18263 4922 18319 4924
rect 18343 4922 18399 4924
rect 18423 4922 18479 4924
rect 18503 4922 18559 4924
rect 18263 4870 18309 4922
rect 18309 4870 18319 4922
rect 18343 4870 18373 4922
rect 18373 4870 18385 4922
rect 18385 4870 18399 4922
rect 18423 4870 18437 4922
rect 18437 4870 18449 4922
rect 18449 4870 18479 4922
rect 18503 4870 18513 4922
rect 18513 4870 18559 4922
rect 18263 4868 18319 4870
rect 18343 4868 18399 4870
rect 18423 4868 18479 4870
rect 18503 4868 18559 4870
rect 10845 4378 10901 4380
rect 10925 4378 10981 4380
rect 11005 4378 11061 4380
rect 11085 4378 11141 4380
rect 10845 4326 10891 4378
rect 10891 4326 10901 4378
rect 10925 4326 10955 4378
rect 10955 4326 10967 4378
rect 10967 4326 10981 4378
rect 11005 4326 11019 4378
rect 11019 4326 11031 4378
rect 11031 4326 11061 4378
rect 11085 4326 11095 4378
rect 11095 4326 11141 4378
rect 10845 4324 10901 4326
rect 10925 4324 10981 4326
rect 11005 4324 11061 4326
rect 11085 4324 11141 4326
rect 15790 4378 15846 4380
rect 15870 4378 15926 4380
rect 15950 4378 16006 4380
rect 16030 4378 16086 4380
rect 15790 4326 15836 4378
rect 15836 4326 15846 4378
rect 15870 4326 15900 4378
rect 15900 4326 15912 4378
rect 15912 4326 15926 4378
rect 15950 4326 15964 4378
rect 15964 4326 15976 4378
rect 15976 4326 16006 4378
rect 16030 4326 16040 4378
rect 16040 4326 16086 4378
rect 15790 4324 15846 4326
rect 15870 4324 15926 4326
rect 15950 4324 16006 4326
rect 16030 4324 16086 4326
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13558 3834 13614 3836
rect 13318 3782 13364 3834
rect 13364 3782 13374 3834
rect 13398 3782 13428 3834
rect 13428 3782 13440 3834
rect 13440 3782 13454 3834
rect 13478 3782 13492 3834
rect 13492 3782 13504 3834
rect 13504 3782 13534 3834
rect 13558 3782 13568 3834
rect 13568 3782 13614 3834
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 13558 3780 13614 3782
rect 18263 3834 18319 3836
rect 18343 3834 18399 3836
rect 18423 3834 18479 3836
rect 18503 3834 18559 3836
rect 18263 3782 18309 3834
rect 18309 3782 18319 3834
rect 18343 3782 18373 3834
rect 18373 3782 18385 3834
rect 18385 3782 18399 3834
rect 18423 3782 18437 3834
rect 18437 3782 18449 3834
rect 18449 3782 18479 3834
rect 18503 3782 18513 3834
rect 18513 3782 18559 3834
rect 18263 3780 18319 3782
rect 18343 3780 18399 3782
rect 18423 3780 18479 3782
rect 18503 3780 18559 3782
rect 10845 3290 10901 3292
rect 10925 3290 10981 3292
rect 11005 3290 11061 3292
rect 11085 3290 11141 3292
rect 10845 3238 10891 3290
rect 10891 3238 10901 3290
rect 10925 3238 10955 3290
rect 10955 3238 10967 3290
rect 10967 3238 10981 3290
rect 11005 3238 11019 3290
rect 11019 3238 11031 3290
rect 11031 3238 11061 3290
rect 11085 3238 11095 3290
rect 11095 3238 11141 3290
rect 10845 3236 10901 3238
rect 10925 3236 10981 3238
rect 11005 3236 11061 3238
rect 11085 3236 11141 3238
rect 15790 3290 15846 3292
rect 15870 3290 15926 3292
rect 15950 3290 16006 3292
rect 16030 3290 16086 3292
rect 15790 3238 15836 3290
rect 15836 3238 15846 3290
rect 15870 3238 15900 3290
rect 15900 3238 15912 3290
rect 15912 3238 15926 3290
rect 15950 3238 15964 3290
rect 15964 3238 15976 3290
rect 15976 3238 16006 3290
rect 16030 3238 16040 3290
rect 16040 3238 16086 3290
rect 15790 3236 15846 3238
rect 15870 3236 15926 3238
rect 15950 3236 16006 3238
rect 16030 3236 16086 3238
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13558 2746 13614 2748
rect 13318 2694 13364 2746
rect 13364 2694 13374 2746
rect 13398 2694 13428 2746
rect 13428 2694 13440 2746
rect 13440 2694 13454 2746
rect 13478 2694 13492 2746
rect 13492 2694 13504 2746
rect 13504 2694 13534 2746
rect 13558 2694 13568 2746
rect 13568 2694 13614 2746
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 13558 2692 13614 2694
rect 18263 2746 18319 2748
rect 18343 2746 18399 2748
rect 18423 2746 18479 2748
rect 18503 2746 18559 2748
rect 18263 2694 18309 2746
rect 18309 2694 18319 2746
rect 18343 2694 18373 2746
rect 18373 2694 18385 2746
rect 18385 2694 18399 2746
rect 18423 2694 18437 2746
rect 18437 2694 18449 2746
rect 18449 2694 18479 2746
rect 18503 2694 18513 2746
rect 18513 2694 18559 2746
rect 18263 2692 18319 2694
rect 18343 2692 18399 2694
rect 18423 2692 18479 2694
rect 18503 2692 18559 2694
rect 20735 7642 20791 7644
rect 20815 7642 20871 7644
rect 20895 7642 20951 7644
rect 20975 7642 21031 7644
rect 20735 7590 20781 7642
rect 20781 7590 20791 7642
rect 20815 7590 20845 7642
rect 20845 7590 20857 7642
rect 20857 7590 20871 7642
rect 20895 7590 20909 7642
rect 20909 7590 20921 7642
rect 20921 7590 20951 7642
rect 20975 7590 20985 7642
rect 20985 7590 21031 7642
rect 20735 7588 20791 7590
rect 20815 7588 20871 7590
rect 20895 7588 20951 7590
rect 20975 7588 21031 7590
rect 20735 6554 20791 6556
rect 20815 6554 20871 6556
rect 20895 6554 20951 6556
rect 20975 6554 21031 6556
rect 20735 6502 20781 6554
rect 20781 6502 20791 6554
rect 20815 6502 20845 6554
rect 20845 6502 20857 6554
rect 20857 6502 20871 6554
rect 20895 6502 20909 6554
rect 20909 6502 20921 6554
rect 20921 6502 20951 6554
rect 20975 6502 20985 6554
rect 20985 6502 21031 6554
rect 20735 6500 20791 6502
rect 20815 6500 20871 6502
rect 20895 6500 20951 6502
rect 20975 6500 21031 6502
rect 20735 5466 20791 5468
rect 20815 5466 20871 5468
rect 20895 5466 20951 5468
rect 20975 5466 21031 5468
rect 20735 5414 20781 5466
rect 20781 5414 20791 5466
rect 20815 5414 20845 5466
rect 20845 5414 20857 5466
rect 20857 5414 20871 5466
rect 20895 5414 20909 5466
rect 20909 5414 20921 5466
rect 20921 5414 20951 5466
rect 20975 5414 20985 5466
rect 20985 5414 21031 5466
rect 20735 5412 20791 5414
rect 20815 5412 20871 5414
rect 20895 5412 20951 5414
rect 20975 5412 21031 5414
rect 20735 4378 20791 4380
rect 20815 4378 20871 4380
rect 20895 4378 20951 4380
rect 20975 4378 21031 4380
rect 20735 4326 20781 4378
rect 20781 4326 20791 4378
rect 20815 4326 20845 4378
rect 20845 4326 20857 4378
rect 20857 4326 20871 4378
rect 20895 4326 20909 4378
rect 20909 4326 20921 4378
rect 20921 4326 20951 4378
rect 20975 4326 20985 4378
rect 20985 4326 21031 4378
rect 20735 4324 20791 4326
rect 20815 4324 20871 4326
rect 20895 4324 20951 4326
rect 20975 4324 21031 4326
rect 20735 3290 20791 3292
rect 20815 3290 20871 3292
rect 20895 3290 20951 3292
rect 20975 3290 21031 3292
rect 20735 3238 20781 3290
rect 20781 3238 20791 3290
rect 20815 3238 20845 3290
rect 20845 3238 20857 3290
rect 20857 3238 20871 3290
rect 20895 3238 20909 3290
rect 20909 3238 20921 3290
rect 20921 3238 20951 3290
rect 20975 3238 20985 3290
rect 20985 3238 21031 3290
rect 20735 3236 20791 3238
rect 20815 3236 20871 3238
rect 20895 3236 20951 3238
rect 20975 3236 21031 3238
rect 10845 2202 10901 2204
rect 10925 2202 10981 2204
rect 11005 2202 11061 2204
rect 11085 2202 11141 2204
rect 10845 2150 10891 2202
rect 10891 2150 10901 2202
rect 10925 2150 10955 2202
rect 10955 2150 10967 2202
rect 10967 2150 10981 2202
rect 11005 2150 11019 2202
rect 11019 2150 11031 2202
rect 11031 2150 11061 2202
rect 11085 2150 11095 2202
rect 11095 2150 11141 2202
rect 10845 2148 10901 2150
rect 10925 2148 10981 2150
rect 11005 2148 11061 2150
rect 11085 2148 11141 2150
rect 15790 2202 15846 2204
rect 15870 2202 15926 2204
rect 15950 2202 16006 2204
rect 16030 2202 16086 2204
rect 15790 2150 15836 2202
rect 15836 2150 15846 2202
rect 15870 2150 15900 2202
rect 15900 2150 15912 2202
rect 15912 2150 15926 2202
rect 15950 2150 15964 2202
rect 15964 2150 15976 2202
rect 15976 2150 16006 2202
rect 16030 2150 16040 2202
rect 16040 2150 16086 2202
rect 15790 2148 15846 2150
rect 15870 2148 15926 2150
rect 15950 2148 16006 2150
rect 16030 2148 16086 2150
rect 20735 2202 20791 2204
rect 20815 2202 20871 2204
rect 20895 2202 20951 2204
rect 20975 2202 21031 2204
rect 20735 2150 20781 2202
rect 20781 2150 20791 2202
rect 20815 2150 20845 2202
rect 20845 2150 20857 2202
rect 20857 2150 20871 2202
rect 20895 2150 20909 2202
rect 20909 2150 20921 2202
rect 20921 2150 20951 2202
rect 20975 2150 20985 2202
rect 20985 2150 21031 2202
rect 20735 2148 20791 2150
rect 20815 2148 20871 2150
rect 20895 2148 20951 2150
rect 20975 2148 21031 2150
<< metal3 >>
rect 5890 19616 6206 19617
rect 5890 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6206 19616
rect 5890 19551 6206 19552
rect 10835 19616 11151 19617
rect 10835 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11151 19616
rect 10835 19551 11151 19552
rect 15780 19616 16096 19617
rect 15780 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16096 19616
rect 15780 19551 16096 19552
rect 20725 19616 21041 19617
rect 20725 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21041 19616
rect 20725 19551 21041 19552
rect 3418 19072 3734 19073
rect 3418 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3734 19072
rect 3418 19007 3734 19008
rect 8363 19072 8679 19073
rect 8363 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8679 19072
rect 8363 19007 8679 19008
rect 13308 19072 13624 19073
rect 13308 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13624 19072
rect 13308 19007 13624 19008
rect 18253 19072 18569 19073
rect 18253 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18569 19072
rect 18253 19007 18569 19008
rect 5890 18528 6206 18529
rect 5890 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6206 18528
rect 5890 18463 6206 18464
rect 10835 18528 11151 18529
rect 10835 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11151 18528
rect 10835 18463 11151 18464
rect 15780 18528 16096 18529
rect 15780 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16096 18528
rect 15780 18463 16096 18464
rect 20725 18528 21041 18529
rect 20725 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21041 18528
rect 20725 18463 21041 18464
rect 10961 18186 11027 18189
rect 14641 18186 14707 18189
rect 15837 18186 15903 18189
rect 16849 18186 16915 18189
rect 10961 18184 16915 18186
rect 10961 18128 10966 18184
rect 11022 18128 14646 18184
rect 14702 18128 15842 18184
rect 15898 18128 16854 18184
rect 16910 18128 16915 18184
rect 10961 18126 16915 18128
rect 10961 18123 11027 18126
rect 14641 18123 14707 18126
rect 15837 18123 15903 18126
rect 16849 18123 16915 18126
rect 3418 17984 3734 17985
rect 3418 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3734 17984
rect 3418 17919 3734 17920
rect 8363 17984 8679 17985
rect 8363 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8679 17984
rect 8363 17919 8679 17920
rect 13308 17984 13624 17985
rect 13308 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13624 17984
rect 13308 17919 13624 17920
rect 18253 17984 18569 17985
rect 18253 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18569 17984
rect 18253 17919 18569 17920
rect 5890 17440 6206 17441
rect 5890 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6206 17440
rect 5890 17375 6206 17376
rect 10835 17440 11151 17441
rect 10835 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11151 17440
rect 10835 17375 11151 17376
rect 15780 17440 16096 17441
rect 15780 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16096 17440
rect 15780 17375 16096 17376
rect 20725 17440 21041 17441
rect 20725 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21041 17440
rect 20725 17375 21041 17376
rect 3418 16896 3734 16897
rect 3418 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3734 16896
rect 3418 16831 3734 16832
rect 8363 16896 8679 16897
rect 8363 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8679 16896
rect 8363 16831 8679 16832
rect 13308 16896 13624 16897
rect 13308 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13624 16896
rect 13308 16831 13624 16832
rect 18253 16896 18569 16897
rect 18253 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18569 16896
rect 18253 16831 18569 16832
rect 5890 16352 6206 16353
rect 5890 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6206 16352
rect 5890 16287 6206 16288
rect 10835 16352 11151 16353
rect 10835 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11151 16352
rect 10835 16287 11151 16288
rect 15780 16352 16096 16353
rect 15780 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16096 16352
rect 15780 16287 16096 16288
rect 20725 16352 21041 16353
rect 20725 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21041 16352
rect 20725 16287 21041 16288
rect 9581 16146 9647 16149
rect 20069 16146 20135 16149
rect 9581 16144 20135 16146
rect 9581 16088 9586 16144
rect 9642 16088 20074 16144
rect 20130 16088 20135 16144
rect 9581 16086 20135 16088
rect 9581 16083 9647 16086
rect 20069 16083 20135 16086
rect 3418 15808 3734 15809
rect 3418 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3734 15808
rect 3418 15743 3734 15744
rect 8363 15808 8679 15809
rect 8363 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8679 15808
rect 8363 15743 8679 15744
rect 13308 15808 13624 15809
rect 13308 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13624 15808
rect 13308 15743 13624 15744
rect 18253 15808 18569 15809
rect 18253 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18569 15808
rect 18253 15743 18569 15744
rect 5890 15264 6206 15265
rect 5890 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6206 15264
rect 5890 15199 6206 15200
rect 10835 15264 11151 15265
rect 10835 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11151 15264
rect 10835 15199 11151 15200
rect 15780 15264 16096 15265
rect 15780 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16096 15264
rect 15780 15199 16096 15200
rect 20725 15264 21041 15265
rect 20725 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21041 15264
rect 20725 15199 21041 15200
rect 3418 14720 3734 14721
rect 3418 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3734 14720
rect 3418 14655 3734 14656
rect 8363 14720 8679 14721
rect 8363 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8679 14720
rect 8363 14655 8679 14656
rect 13308 14720 13624 14721
rect 13308 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13624 14720
rect 13308 14655 13624 14656
rect 18253 14720 18569 14721
rect 18253 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18569 14720
rect 18253 14655 18569 14656
rect 5890 14176 6206 14177
rect 5890 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6206 14176
rect 5890 14111 6206 14112
rect 10835 14176 11151 14177
rect 10835 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11151 14176
rect 10835 14111 11151 14112
rect 15780 14176 16096 14177
rect 15780 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16096 14176
rect 15780 14111 16096 14112
rect 20725 14176 21041 14177
rect 20725 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21041 14176
rect 20725 14111 21041 14112
rect 3418 13632 3734 13633
rect 3418 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3734 13632
rect 3418 13567 3734 13568
rect 8363 13632 8679 13633
rect 8363 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8679 13632
rect 8363 13567 8679 13568
rect 13308 13632 13624 13633
rect 13308 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13624 13632
rect 13308 13567 13624 13568
rect 18253 13632 18569 13633
rect 18253 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18569 13632
rect 18253 13567 18569 13568
rect 5890 13088 6206 13089
rect 5890 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6206 13088
rect 5890 13023 6206 13024
rect 10835 13088 11151 13089
rect 10835 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11151 13088
rect 10835 13023 11151 13024
rect 15780 13088 16096 13089
rect 15780 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16096 13088
rect 15780 13023 16096 13024
rect 20725 13088 21041 13089
rect 20725 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21041 13088
rect 20725 13023 21041 13024
rect 3418 12544 3734 12545
rect 3418 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3734 12544
rect 3418 12479 3734 12480
rect 8363 12544 8679 12545
rect 8363 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8679 12544
rect 8363 12479 8679 12480
rect 13308 12544 13624 12545
rect 13308 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13624 12544
rect 13308 12479 13624 12480
rect 18253 12544 18569 12545
rect 18253 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18569 12544
rect 18253 12479 18569 12480
rect 5890 12000 6206 12001
rect 5890 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6206 12000
rect 5890 11935 6206 11936
rect 10835 12000 11151 12001
rect 10835 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11151 12000
rect 10835 11935 11151 11936
rect 15780 12000 16096 12001
rect 15780 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16096 12000
rect 15780 11935 16096 11936
rect 20725 12000 21041 12001
rect 20725 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21041 12000
rect 20725 11935 21041 11936
rect 15469 11794 15535 11797
rect 19241 11794 19307 11797
rect 15469 11792 19307 11794
rect 15469 11736 15474 11792
rect 15530 11736 19246 11792
rect 19302 11736 19307 11792
rect 15469 11734 19307 11736
rect 15469 11731 15535 11734
rect 19241 11731 19307 11734
rect 3418 11456 3734 11457
rect 3418 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3734 11456
rect 3418 11391 3734 11392
rect 8363 11456 8679 11457
rect 8363 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8679 11456
rect 8363 11391 8679 11392
rect 13308 11456 13624 11457
rect 13308 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13624 11456
rect 13308 11391 13624 11392
rect 18253 11456 18569 11457
rect 18253 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18569 11456
rect 18253 11391 18569 11392
rect 5890 10912 6206 10913
rect 5890 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6206 10912
rect 5890 10847 6206 10848
rect 10835 10912 11151 10913
rect 10835 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11151 10912
rect 10835 10847 11151 10848
rect 15780 10912 16096 10913
rect 15780 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16096 10912
rect 15780 10847 16096 10848
rect 20725 10912 21041 10913
rect 20725 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21041 10912
rect 20725 10847 21041 10848
rect 3418 10368 3734 10369
rect 3418 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3734 10368
rect 3418 10303 3734 10304
rect 8363 10368 8679 10369
rect 8363 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8679 10368
rect 8363 10303 8679 10304
rect 13308 10368 13624 10369
rect 13308 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13624 10368
rect 13308 10303 13624 10304
rect 18253 10368 18569 10369
rect 18253 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18569 10368
rect 18253 10303 18569 10304
rect 5890 9824 6206 9825
rect 5890 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6206 9824
rect 5890 9759 6206 9760
rect 10835 9824 11151 9825
rect 10835 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11151 9824
rect 10835 9759 11151 9760
rect 15780 9824 16096 9825
rect 15780 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16096 9824
rect 15780 9759 16096 9760
rect 20725 9824 21041 9825
rect 20725 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21041 9824
rect 20725 9759 21041 9760
rect 3418 9280 3734 9281
rect 3418 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3734 9280
rect 3418 9215 3734 9216
rect 8363 9280 8679 9281
rect 8363 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8679 9280
rect 8363 9215 8679 9216
rect 13308 9280 13624 9281
rect 13308 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13624 9280
rect 13308 9215 13624 9216
rect 18253 9280 18569 9281
rect 18253 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18569 9280
rect 18253 9215 18569 9216
rect 5890 8736 6206 8737
rect 5890 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6206 8736
rect 5890 8671 6206 8672
rect 10835 8736 11151 8737
rect 10835 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11151 8736
rect 10835 8671 11151 8672
rect 15780 8736 16096 8737
rect 15780 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16096 8736
rect 15780 8671 16096 8672
rect 20725 8736 21041 8737
rect 20725 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21041 8736
rect 20725 8671 21041 8672
rect 3418 8192 3734 8193
rect 3418 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3734 8192
rect 3418 8127 3734 8128
rect 8363 8192 8679 8193
rect 8363 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8679 8192
rect 8363 8127 8679 8128
rect 13308 8192 13624 8193
rect 13308 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13624 8192
rect 13308 8127 13624 8128
rect 18253 8192 18569 8193
rect 18253 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18569 8192
rect 18253 8127 18569 8128
rect 11053 7850 11119 7853
rect 11421 7850 11487 7853
rect 19885 7850 19951 7853
rect 11053 7848 19951 7850
rect 11053 7792 11058 7848
rect 11114 7792 11426 7848
rect 11482 7792 19890 7848
rect 19946 7792 19951 7848
rect 11053 7790 19951 7792
rect 11053 7787 11119 7790
rect 11421 7787 11487 7790
rect 19885 7787 19951 7790
rect 5890 7648 6206 7649
rect 5890 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6206 7648
rect 5890 7583 6206 7584
rect 10835 7648 11151 7649
rect 10835 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11151 7648
rect 10835 7583 11151 7584
rect 15780 7648 16096 7649
rect 15780 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16096 7648
rect 15780 7583 16096 7584
rect 20725 7648 21041 7649
rect 20725 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21041 7648
rect 20725 7583 21041 7584
rect 3418 7104 3734 7105
rect 3418 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3734 7104
rect 3418 7039 3734 7040
rect 8363 7104 8679 7105
rect 8363 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8679 7104
rect 8363 7039 8679 7040
rect 13308 7104 13624 7105
rect 13308 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13624 7104
rect 13308 7039 13624 7040
rect 18253 7104 18569 7105
rect 18253 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18569 7104
rect 18253 7039 18569 7040
rect 5890 6560 6206 6561
rect 5890 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6206 6560
rect 5890 6495 6206 6496
rect 10835 6560 11151 6561
rect 10835 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11151 6560
rect 10835 6495 11151 6496
rect 15780 6560 16096 6561
rect 15780 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16096 6560
rect 15780 6495 16096 6496
rect 20725 6560 21041 6561
rect 20725 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21041 6560
rect 20725 6495 21041 6496
rect 3418 6016 3734 6017
rect 3418 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3734 6016
rect 3418 5951 3734 5952
rect 8363 6016 8679 6017
rect 8363 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8679 6016
rect 8363 5951 8679 5952
rect 13308 6016 13624 6017
rect 13308 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13624 6016
rect 13308 5951 13624 5952
rect 18253 6016 18569 6017
rect 18253 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18569 6016
rect 18253 5951 18569 5952
rect 5890 5472 6206 5473
rect 5890 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6206 5472
rect 5890 5407 6206 5408
rect 10835 5472 11151 5473
rect 10835 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11151 5472
rect 10835 5407 11151 5408
rect 15780 5472 16096 5473
rect 15780 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16096 5472
rect 15780 5407 16096 5408
rect 20725 5472 21041 5473
rect 20725 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21041 5472
rect 20725 5407 21041 5408
rect 3418 4928 3734 4929
rect 3418 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3734 4928
rect 3418 4863 3734 4864
rect 8363 4928 8679 4929
rect 8363 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8679 4928
rect 8363 4863 8679 4864
rect 13308 4928 13624 4929
rect 13308 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13624 4928
rect 13308 4863 13624 4864
rect 18253 4928 18569 4929
rect 18253 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18569 4928
rect 18253 4863 18569 4864
rect 5890 4384 6206 4385
rect 5890 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6206 4384
rect 5890 4319 6206 4320
rect 10835 4384 11151 4385
rect 10835 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11151 4384
rect 10835 4319 11151 4320
rect 15780 4384 16096 4385
rect 15780 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16096 4384
rect 15780 4319 16096 4320
rect 20725 4384 21041 4385
rect 20725 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21041 4384
rect 20725 4319 21041 4320
rect 3418 3840 3734 3841
rect 3418 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3734 3840
rect 3418 3775 3734 3776
rect 8363 3840 8679 3841
rect 8363 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8679 3840
rect 8363 3775 8679 3776
rect 13308 3840 13624 3841
rect 13308 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13624 3840
rect 13308 3775 13624 3776
rect 18253 3840 18569 3841
rect 18253 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18569 3840
rect 18253 3775 18569 3776
rect 5890 3296 6206 3297
rect 5890 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6206 3296
rect 5890 3231 6206 3232
rect 10835 3296 11151 3297
rect 10835 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11151 3296
rect 10835 3231 11151 3232
rect 15780 3296 16096 3297
rect 15780 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16096 3296
rect 15780 3231 16096 3232
rect 20725 3296 21041 3297
rect 20725 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21041 3296
rect 20725 3231 21041 3232
rect 3418 2752 3734 2753
rect 3418 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3734 2752
rect 3418 2687 3734 2688
rect 8363 2752 8679 2753
rect 8363 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8679 2752
rect 8363 2687 8679 2688
rect 13308 2752 13624 2753
rect 13308 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13624 2752
rect 13308 2687 13624 2688
rect 18253 2752 18569 2753
rect 18253 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18569 2752
rect 18253 2687 18569 2688
rect 5890 2208 6206 2209
rect 5890 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6206 2208
rect 5890 2143 6206 2144
rect 10835 2208 11151 2209
rect 10835 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11151 2208
rect 10835 2143 11151 2144
rect 15780 2208 16096 2209
rect 15780 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16096 2208
rect 15780 2143 16096 2144
rect 20725 2208 21041 2209
rect 20725 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21041 2208
rect 20725 2143 21041 2144
<< via3 >>
rect 5896 19612 5960 19616
rect 5896 19556 5900 19612
rect 5900 19556 5956 19612
rect 5956 19556 5960 19612
rect 5896 19552 5960 19556
rect 5976 19612 6040 19616
rect 5976 19556 5980 19612
rect 5980 19556 6036 19612
rect 6036 19556 6040 19612
rect 5976 19552 6040 19556
rect 6056 19612 6120 19616
rect 6056 19556 6060 19612
rect 6060 19556 6116 19612
rect 6116 19556 6120 19612
rect 6056 19552 6120 19556
rect 6136 19612 6200 19616
rect 6136 19556 6140 19612
rect 6140 19556 6196 19612
rect 6196 19556 6200 19612
rect 6136 19552 6200 19556
rect 10841 19612 10905 19616
rect 10841 19556 10845 19612
rect 10845 19556 10901 19612
rect 10901 19556 10905 19612
rect 10841 19552 10905 19556
rect 10921 19612 10985 19616
rect 10921 19556 10925 19612
rect 10925 19556 10981 19612
rect 10981 19556 10985 19612
rect 10921 19552 10985 19556
rect 11001 19612 11065 19616
rect 11001 19556 11005 19612
rect 11005 19556 11061 19612
rect 11061 19556 11065 19612
rect 11001 19552 11065 19556
rect 11081 19612 11145 19616
rect 11081 19556 11085 19612
rect 11085 19556 11141 19612
rect 11141 19556 11145 19612
rect 11081 19552 11145 19556
rect 15786 19612 15850 19616
rect 15786 19556 15790 19612
rect 15790 19556 15846 19612
rect 15846 19556 15850 19612
rect 15786 19552 15850 19556
rect 15866 19612 15930 19616
rect 15866 19556 15870 19612
rect 15870 19556 15926 19612
rect 15926 19556 15930 19612
rect 15866 19552 15930 19556
rect 15946 19612 16010 19616
rect 15946 19556 15950 19612
rect 15950 19556 16006 19612
rect 16006 19556 16010 19612
rect 15946 19552 16010 19556
rect 16026 19612 16090 19616
rect 16026 19556 16030 19612
rect 16030 19556 16086 19612
rect 16086 19556 16090 19612
rect 16026 19552 16090 19556
rect 20731 19612 20795 19616
rect 20731 19556 20735 19612
rect 20735 19556 20791 19612
rect 20791 19556 20795 19612
rect 20731 19552 20795 19556
rect 20811 19612 20875 19616
rect 20811 19556 20815 19612
rect 20815 19556 20871 19612
rect 20871 19556 20875 19612
rect 20811 19552 20875 19556
rect 20891 19612 20955 19616
rect 20891 19556 20895 19612
rect 20895 19556 20951 19612
rect 20951 19556 20955 19612
rect 20891 19552 20955 19556
rect 20971 19612 21035 19616
rect 20971 19556 20975 19612
rect 20975 19556 21031 19612
rect 21031 19556 21035 19612
rect 20971 19552 21035 19556
rect 3424 19068 3488 19072
rect 3424 19012 3428 19068
rect 3428 19012 3484 19068
rect 3484 19012 3488 19068
rect 3424 19008 3488 19012
rect 3504 19068 3568 19072
rect 3504 19012 3508 19068
rect 3508 19012 3564 19068
rect 3564 19012 3568 19068
rect 3504 19008 3568 19012
rect 3584 19068 3648 19072
rect 3584 19012 3588 19068
rect 3588 19012 3644 19068
rect 3644 19012 3648 19068
rect 3584 19008 3648 19012
rect 3664 19068 3728 19072
rect 3664 19012 3668 19068
rect 3668 19012 3724 19068
rect 3724 19012 3728 19068
rect 3664 19008 3728 19012
rect 8369 19068 8433 19072
rect 8369 19012 8373 19068
rect 8373 19012 8429 19068
rect 8429 19012 8433 19068
rect 8369 19008 8433 19012
rect 8449 19068 8513 19072
rect 8449 19012 8453 19068
rect 8453 19012 8509 19068
rect 8509 19012 8513 19068
rect 8449 19008 8513 19012
rect 8529 19068 8593 19072
rect 8529 19012 8533 19068
rect 8533 19012 8589 19068
rect 8589 19012 8593 19068
rect 8529 19008 8593 19012
rect 8609 19068 8673 19072
rect 8609 19012 8613 19068
rect 8613 19012 8669 19068
rect 8669 19012 8673 19068
rect 8609 19008 8673 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 13554 19068 13618 19072
rect 13554 19012 13558 19068
rect 13558 19012 13614 19068
rect 13614 19012 13618 19068
rect 13554 19008 13618 19012
rect 18259 19068 18323 19072
rect 18259 19012 18263 19068
rect 18263 19012 18319 19068
rect 18319 19012 18323 19068
rect 18259 19008 18323 19012
rect 18339 19068 18403 19072
rect 18339 19012 18343 19068
rect 18343 19012 18399 19068
rect 18399 19012 18403 19068
rect 18339 19008 18403 19012
rect 18419 19068 18483 19072
rect 18419 19012 18423 19068
rect 18423 19012 18479 19068
rect 18479 19012 18483 19068
rect 18419 19008 18483 19012
rect 18499 19068 18563 19072
rect 18499 19012 18503 19068
rect 18503 19012 18559 19068
rect 18559 19012 18563 19068
rect 18499 19008 18563 19012
rect 5896 18524 5960 18528
rect 5896 18468 5900 18524
rect 5900 18468 5956 18524
rect 5956 18468 5960 18524
rect 5896 18464 5960 18468
rect 5976 18524 6040 18528
rect 5976 18468 5980 18524
rect 5980 18468 6036 18524
rect 6036 18468 6040 18524
rect 5976 18464 6040 18468
rect 6056 18524 6120 18528
rect 6056 18468 6060 18524
rect 6060 18468 6116 18524
rect 6116 18468 6120 18524
rect 6056 18464 6120 18468
rect 6136 18524 6200 18528
rect 6136 18468 6140 18524
rect 6140 18468 6196 18524
rect 6196 18468 6200 18524
rect 6136 18464 6200 18468
rect 10841 18524 10905 18528
rect 10841 18468 10845 18524
rect 10845 18468 10901 18524
rect 10901 18468 10905 18524
rect 10841 18464 10905 18468
rect 10921 18524 10985 18528
rect 10921 18468 10925 18524
rect 10925 18468 10981 18524
rect 10981 18468 10985 18524
rect 10921 18464 10985 18468
rect 11001 18524 11065 18528
rect 11001 18468 11005 18524
rect 11005 18468 11061 18524
rect 11061 18468 11065 18524
rect 11001 18464 11065 18468
rect 11081 18524 11145 18528
rect 11081 18468 11085 18524
rect 11085 18468 11141 18524
rect 11141 18468 11145 18524
rect 11081 18464 11145 18468
rect 15786 18524 15850 18528
rect 15786 18468 15790 18524
rect 15790 18468 15846 18524
rect 15846 18468 15850 18524
rect 15786 18464 15850 18468
rect 15866 18524 15930 18528
rect 15866 18468 15870 18524
rect 15870 18468 15926 18524
rect 15926 18468 15930 18524
rect 15866 18464 15930 18468
rect 15946 18524 16010 18528
rect 15946 18468 15950 18524
rect 15950 18468 16006 18524
rect 16006 18468 16010 18524
rect 15946 18464 16010 18468
rect 16026 18524 16090 18528
rect 16026 18468 16030 18524
rect 16030 18468 16086 18524
rect 16086 18468 16090 18524
rect 16026 18464 16090 18468
rect 20731 18524 20795 18528
rect 20731 18468 20735 18524
rect 20735 18468 20791 18524
rect 20791 18468 20795 18524
rect 20731 18464 20795 18468
rect 20811 18524 20875 18528
rect 20811 18468 20815 18524
rect 20815 18468 20871 18524
rect 20871 18468 20875 18524
rect 20811 18464 20875 18468
rect 20891 18524 20955 18528
rect 20891 18468 20895 18524
rect 20895 18468 20951 18524
rect 20951 18468 20955 18524
rect 20891 18464 20955 18468
rect 20971 18524 21035 18528
rect 20971 18468 20975 18524
rect 20975 18468 21031 18524
rect 21031 18468 21035 18524
rect 20971 18464 21035 18468
rect 3424 17980 3488 17984
rect 3424 17924 3428 17980
rect 3428 17924 3484 17980
rect 3484 17924 3488 17980
rect 3424 17920 3488 17924
rect 3504 17980 3568 17984
rect 3504 17924 3508 17980
rect 3508 17924 3564 17980
rect 3564 17924 3568 17980
rect 3504 17920 3568 17924
rect 3584 17980 3648 17984
rect 3584 17924 3588 17980
rect 3588 17924 3644 17980
rect 3644 17924 3648 17980
rect 3584 17920 3648 17924
rect 3664 17980 3728 17984
rect 3664 17924 3668 17980
rect 3668 17924 3724 17980
rect 3724 17924 3728 17980
rect 3664 17920 3728 17924
rect 8369 17980 8433 17984
rect 8369 17924 8373 17980
rect 8373 17924 8429 17980
rect 8429 17924 8433 17980
rect 8369 17920 8433 17924
rect 8449 17980 8513 17984
rect 8449 17924 8453 17980
rect 8453 17924 8509 17980
rect 8509 17924 8513 17980
rect 8449 17920 8513 17924
rect 8529 17980 8593 17984
rect 8529 17924 8533 17980
rect 8533 17924 8589 17980
rect 8589 17924 8593 17980
rect 8529 17920 8593 17924
rect 8609 17980 8673 17984
rect 8609 17924 8613 17980
rect 8613 17924 8669 17980
rect 8669 17924 8673 17980
rect 8609 17920 8673 17924
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 13554 17980 13618 17984
rect 13554 17924 13558 17980
rect 13558 17924 13614 17980
rect 13614 17924 13618 17980
rect 13554 17920 13618 17924
rect 18259 17980 18323 17984
rect 18259 17924 18263 17980
rect 18263 17924 18319 17980
rect 18319 17924 18323 17980
rect 18259 17920 18323 17924
rect 18339 17980 18403 17984
rect 18339 17924 18343 17980
rect 18343 17924 18399 17980
rect 18399 17924 18403 17980
rect 18339 17920 18403 17924
rect 18419 17980 18483 17984
rect 18419 17924 18423 17980
rect 18423 17924 18479 17980
rect 18479 17924 18483 17980
rect 18419 17920 18483 17924
rect 18499 17980 18563 17984
rect 18499 17924 18503 17980
rect 18503 17924 18559 17980
rect 18559 17924 18563 17980
rect 18499 17920 18563 17924
rect 5896 17436 5960 17440
rect 5896 17380 5900 17436
rect 5900 17380 5956 17436
rect 5956 17380 5960 17436
rect 5896 17376 5960 17380
rect 5976 17436 6040 17440
rect 5976 17380 5980 17436
rect 5980 17380 6036 17436
rect 6036 17380 6040 17436
rect 5976 17376 6040 17380
rect 6056 17436 6120 17440
rect 6056 17380 6060 17436
rect 6060 17380 6116 17436
rect 6116 17380 6120 17436
rect 6056 17376 6120 17380
rect 6136 17436 6200 17440
rect 6136 17380 6140 17436
rect 6140 17380 6196 17436
rect 6196 17380 6200 17436
rect 6136 17376 6200 17380
rect 10841 17436 10905 17440
rect 10841 17380 10845 17436
rect 10845 17380 10901 17436
rect 10901 17380 10905 17436
rect 10841 17376 10905 17380
rect 10921 17436 10985 17440
rect 10921 17380 10925 17436
rect 10925 17380 10981 17436
rect 10981 17380 10985 17436
rect 10921 17376 10985 17380
rect 11001 17436 11065 17440
rect 11001 17380 11005 17436
rect 11005 17380 11061 17436
rect 11061 17380 11065 17436
rect 11001 17376 11065 17380
rect 11081 17436 11145 17440
rect 11081 17380 11085 17436
rect 11085 17380 11141 17436
rect 11141 17380 11145 17436
rect 11081 17376 11145 17380
rect 15786 17436 15850 17440
rect 15786 17380 15790 17436
rect 15790 17380 15846 17436
rect 15846 17380 15850 17436
rect 15786 17376 15850 17380
rect 15866 17436 15930 17440
rect 15866 17380 15870 17436
rect 15870 17380 15926 17436
rect 15926 17380 15930 17436
rect 15866 17376 15930 17380
rect 15946 17436 16010 17440
rect 15946 17380 15950 17436
rect 15950 17380 16006 17436
rect 16006 17380 16010 17436
rect 15946 17376 16010 17380
rect 16026 17436 16090 17440
rect 16026 17380 16030 17436
rect 16030 17380 16086 17436
rect 16086 17380 16090 17436
rect 16026 17376 16090 17380
rect 20731 17436 20795 17440
rect 20731 17380 20735 17436
rect 20735 17380 20791 17436
rect 20791 17380 20795 17436
rect 20731 17376 20795 17380
rect 20811 17436 20875 17440
rect 20811 17380 20815 17436
rect 20815 17380 20871 17436
rect 20871 17380 20875 17436
rect 20811 17376 20875 17380
rect 20891 17436 20955 17440
rect 20891 17380 20895 17436
rect 20895 17380 20951 17436
rect 20951 17380 20955 17436
rect 20891 17376 20955 17380
rect 20971 17436 21035 17440
rect 20971 17380 20975 17436
rect 20975 17380 21031 17436
rect 21031 17380 21035 17436
rect 20971 17376 21035 17380
rect 3424 16892 3488 16896
rect 3424 16836 3428 16892
rect 3428 16836 3484 16892
rect 3484 16836 3488 16892
rect 3424 16832 3488 16836
rect 3504 16892 3568 16896
rect 3504 16836 3508 16892
rect 3508 16836 3564 16892
rect 3564 16836 3568 16892
rect 3504 16832 3568 16836
rect 3584 16892 3648 16896
rect 3584 16836 3588 16892
rect 3588 16836 3644 16892
rect 3644 16836 3648 16892
rect 3584 16832 3648 16836
rect 3664 16892 3728 16896
rect 3664 16836 3668 16892
rect 3668 16836 3724 16892
rect 3724 16836 3728 16892
rect 3664 16832 3728 16836
rect 8369 16892 8433 16896
rect 8369 16836 8373 16892
rect 8373 16836 8429 16892
rect 8429 16836 8433 16892
rect 8369 16832 8433 16836
rect 8449 16892 8513 16896
rect 8449 16836 8453 16892
rect 8453 16836 8509 16892
rect 8509 16836 8513 16892
rect 8449 16832 8513 16836
rect 8529 16892 8593 16896
rect 8529 16836 8533 16892
rect 8533 16836 8589 16892
rect 8589 16836 8593 16892
rect 8529 16832 8593 16836
rect 8609 16892 8673 16896
rect 8609 16836 8613 16892
rect 8613 16836 8669 16892
rect 8669 16836 8673 16892
rect 8609 16832 8673 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 13554 16892 13618 16896
rect 13554 16836 13558 16892
rect 13558 16836 13614 16892
rect 13614 16836 13618 16892
rect 13554 16832 13618 16836
rect 18259 16892 18323 16896
rect 18259 16836 18263 16892
rect 18263 16836 18319 16892
rect 18319 16836 18323 16892
rect 18259 16832 18323 16836
rect 18339 16892 18403 16896
rect 18339 16836 18343 16892
rect 18343 16836 18399 16892
rect 18399 16836 18403 16892
rect 18339 16832 18403 16836
rect 18419 16892 18483 16896
rect 18419 16836 18423 16892
rect 18423 16836 18479 16892
rect 18479 16836 18483 16892
rect 18419 16832 18483 16836
rect 18499 16892 18563 16896
rect 18499 16836 18503 16892
rect 18503 16836 18559 16892
rect 18559 16836 18563 16892
rect 18499 16832 18563 16836
rect 5896 16348 5960 16352
rect 5896 16292 5900 16348
rect 5900 16292 5956 16348
rect 5956 16292 5960 16348
rect 5896 16288 5960 16292
rect 5976 16348 6040 16352
rect 5976 16292 5980 16348
rect 5980 16292 6036 16348
rect 6036 16292 6040 16348
rect 5976 16288 6040 16292
rect 6056 16348 6120 16352
rect 6056 16292 6060 16348
rect 6060 16292 6116 16348
rect 6116 16292 6120 16348
rect 6056 16288 6120 16292
rect 6136 16348 6200 16352
rect 6136 16292 6140 16348
rect 6140 16292 6196 16348
rect 6196 16292 6200 16348
rect 6136 16288 6200 16292
rect 10841 16348 10905 16352
rect 10841 16292 10845 16348
rect 10845 16292 10901 16348
rect 10901 16292 10905 16348
rect 10841 16288 10905 16292
rect 10921 16348 10985 16352
rect 10921 16292 10925 16348
rect 10925 16292 10981 16348
rect 10981 16292 10985 16348
rect 10921 16288 10985 16292
rect 11001 16348 11065 16352
rect 11001 16292 11005 16348
rect 11005 16292 11061 16348
rect 11061 16292 11065 16348
rect 11001 16288 11065 16292
rect 11081 16348 11145 16352
rect 11081 16292 11085 16348
rect 11085 16292 11141 16348
rect 11141 16292 11145 16348
rect 11081 16288 11145 16292
rect 15786 16348 15850 16352
rect 15786 16292 15790 16348
rect 15790 16292 15846 16348
rect 15846 16292 15850 16348
rect 15786 16288 15850 16292
rect 15866 16348 15930 16352
rect 15866 16292 15870 16348
rect 15870 16292 15926 16348
rect 15926 16292 15930 16348
rect 15866 16288 15930 16292
rect 15946 16348 16010 16352
rect 15946 16292 15950 16348
rect 15950 16292 16006 16348
rect 16006 16292 16010 16348
rect 15946 16288 16010 16292
rect 16026 16348 16090 16352
rect 16026 16292 16030 16348
rect 16030 16292 16086 16348
rect 16086 16292 16090 16348
rect 16026 16288 16090 16292
rect 20731 16348 20795 16352
rect 20731 16292 20735 16348
rect 20735 16292 20791 16348
rect 20791 16292 20795 16348
rect 20731 16288 20795 16292
rect 20811 16348 20875 16352
rect 20811 16292 20815 16348
rect 20815 16292 20871 16348
rect 20871 16292 20875 16348
rect 20811 16288 20875 16292
rect 20891 16348 20955 16352
rect 20891 16292 20895 16348
rect 20895 16292 20951 16348
rect 20951 16292 20955 16348
rect 20891 16288 20955 16292
rect 20971 16348 21035 16352
rect 20971 16292 20975 16348
rect 20975 16292 21031 16348
rect 21031 16292 21035 16348
rect 20971 16288 21035 16292
rect 3424 15804 3488 15808
rect 3424 15748 3428 15804
rect 3428 15748 3484 15804
rect 3484 15748 3488 15804
rect 3424 15744 3488 15748
rect 3504 15804 3568 15808
rect 3504 15748 3508 15804
rect 3508 15748 3564 15804
rect 3564 15748 3568 15804
rect 3504 15744 3568 15748
rect 3584 15804 3648 15808
rect 3584 15748 3588 15804
rect 3588 15748 3644 15804
rect 3644 15748 3648 15804
rect 3584 15744 3648 15748
rect 3664 15804 3728 15808
rect 3664 15748 3668 15804
rect 3668 15748 3724 15804
rect 3724 15748 3728 15804
rect 3664 15744 3728 15748
rect 8369 15804 8433 15808
rect 8369 15748 8373 15804
rect 8373 15748 8429 15804
rect 8429 15748 8433 15804
rect 8369 15744 8433 15748
rect 8449 15804 8513 15808
rect 8449 15748 8453 15804
rect 8453 15748 8509 15804
rect 8509 15748 8513 15804
rect 8449 15744 8513 15748
rect 8529 15804 8593 15808
rect 8529 15748 8533 15804
rect 8533 15748 8589 15804
rect 8589 15748 8593 15804
rect 8529 15744 8593 15748
rect 8609 15804 8673 15808
rect 8609 15748 8613 15804
rect 8613 15748 8669 15804
rect 8669 15748 8673 15804
rect 8609 15744 8673 15748
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 13554 15804 13618 15808
rect 13554 15748 13558 15804
rect 13558 15748 13614 15804
rect 13614 15748 13618 15804
rect 13554 15744 13618 15748
rect 18259 15804 18323 15808
rect 18259 15748 18263 15804
rect 18263 15748 18319 15804
rect 18319 15748 18323 15804
rect 18259 15744 18323 15748
rect 18339 15804 18403 15808
rect 18339 15748 18343 15804
rect 18343 15748 18399 15804
rect 18399 15748 18403 15804
rect 18339 15744 18403 15748
rect 18419 15804 18483 15808
rect 18419 15748 18423 15804
rect 18423 15748 18479 15804
rect 18479 15748 18483 15804
rect 18419 15744 18483 15748
rect 18499 15804 18563 15808
rect 18499 15748 18503 15804
rect 18503 15748 18559 15804
rect 18559 15748 18563 15804
rect 18499 15744 18563 15748
rect 5896 15260 5960 15264
rect 5896 15204 5900 15260
rect 5900 15204 5956 15260
rect 5956 15204 5960 15260
rect 5896 15200 5960 15204
rect 5976 15260 6040 15264
rect 5976 15204 5980 15260
rect 5980 15204 6036 15260
rect 6036 15204 6040 15260
rect 5976 15200 6040 15204
rect 6056 15260 6120 15264
rect 6056 15204 6060 15260
rect 6060 15204 6116 15260
rect 6116 15204 6120 15260
rect 6056 15200 6120 15204
rect 6136 15260 6200 15264
rect 6136 15204 6140 15260
rect 6140 15204 6196 15260
rect 6196 15204 6200 15260
rect 6136 15200 6200 15204
rect 10841 15260 10905 15264
rect 10841 15204 10845 15260
rect 10845 15204 10901 15260
rect 10901 15204 10905 15260
rect 10841 15200 10905 15204
rect 10921 15260 10985 15264
rect 10921 15204 10925 15260
rect 10925 15204 10981 15260
rect 10981 15204 10985 15260
rect 10921 15200 10985 15204
rect 11001 15260 11065 15264
rect 11001 15204 11005 15260
rect 11005 15204 11061 15260
rect 11061 15204 11065 15260
rect 11001 15200 11065 15204
rect 11081 15260 11145 15264
rect 11081 15204 11085 15260
rect 11085 15204 11141 15260
rect 11141 15204 11145 15260
rect 11081 15200 11145 15204
rect 15786 15260 15850 15264
rect 15786 15204 15790 15260
rect 15790 15204 15846 15260
rect 15846 15204 15850 15260
rect 15786 15200 15850 15204
rect 15866 15260 15930 15264
rect 15866 15204 15870 15260
rect 15870 15204 15926 15260
rect 15926 15204 15930 15260
rect 15866 15200 15930 15204
rect 15946 15260 16010 15264
rect 15946 15204 15950 15260
rect 15950 15204 16006 15260
rect 16006 15204 16010 15260
rect 15946 15200 16010 15204
rect 16026 15260 16090 15264
rect 16026 15204 16030 15260
rect 16030 15204 16086 15260
rect 16086 15204 16090 15260
rect 16026 15200 16090 15204
rect 20731 15260 20795 15264
rect 20731 15204 20735 15260
rect 20735 15204 20791 15260
rect 20791 15204 20795 15260
rect 20731 15200 20795 15204
rect 20811 15260 20875 15264
rect 20811 15204 20815 15260
rect 20815 15204 20871 15260
rect 20871 15204 20875 15260
rect 20811 15200 20875 15204
rect 20891 15260 20955 15264
rect 20891 15204 20895 15260
rect 20895 15204 20951 15260
rect 20951 15204 20955 15260
rect 20891 15200 20955 15204
rect 20971 15260 21035 15264
rect 20971 15204 20975 15260
rect 20975 15204 21031 15260
rect 21031 15204 21035 15260
rect 20971 15200 21035 15204
rect 3424 14716 3488 14720
rect 3424 14660 3428 14716
rect 3428 14660 3484 14716
rect 3484 14660 3488 14716
rect 3424 14656 3488 14660
rect 3504 14716 3568 14720
rect 3504 14660 3508 14716
rect 3508 14660 3564 14716
rect 3564 14660 3568 14716
rect 3504 14656 3568 14660
rect 3584 14716 3648 14720
rect 3584 14660 3588 14716
rect 3588 14660 3644 14716
rect 3644 14660 3648 14716
rect 3584 14656 3648 14660
rect 3664 14716 3728 14720
rect 3664 14660 3668 14716
rect 3668 14660 3724 14716
rect 3724 14660 3728 14716
rect 3664 14656 3728 14660
rect 8369 14716 8433 14720
rect 8369 14660 8373 14716
rect 8373 14660 8429 14716
rect 8429 14660 8433 14716
rect 8369 14656 8433 14660
rect 8449 14716 8513 14720
rect 8449 14660 8453 14716
rect 8453 14660 8509 14716
rect 8509 14660 8513 14716
rect 8449 14656 8513 14660
rect 8529 14716 8593 14720
rect 8529 14660 8533 14716
rect 8533 14660 8589 14716
rect 8589 14660 8593 14716
rect 8529 14656 8593 14660
rect 8609 14716 8673 14720
rect 8609 14660 8613 14716
rect 8613 14660 8669 14716
rect 8669 14660 8673 14716
rect 8609 14656 8673 14660
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 13554 14716 13618 14720
rect 13554 14660 13558 14716
rect 13558 14660 13614 14716
rect 13614 14660 13618 14716
rect 13554 14656 13618 14660
rect 18259 14716 18323 14720
rect 18259 14660 18263 14716
rect 18263 14660 18319 14716
rect 18319 14660 18323 14716
rect 18259 14656 18323 14660
rect 18339 14716 18403 14720
rect 18339 14660 18343 14716
rect 18343 14660 18399 14716
rect 18399 14660 18403 14716
rect 18339 14656 18403 14660
rect 18419 14716 18483 14720
rect 18419 14660 18423 14716
rect 18423 14660 18479 14716
rect 18479 14660 18483 14716
rect 18419 14656 18483 14660
rect 18499 14716 18563 14720
rect 18499 14660 18503 14716
rect 18503 14660 18559 14716
rect 18559 14660 18563 14716
rect 18499 14656 18563 14660
rect 5896 14172 5960 14176
rect 5896 14116 5900 14172
rect 5900 14116 5956 14172
rect 5956 14116 5960 14172
rect 5896 14112 5960 14116
rect 5976 14172 6040 14176
rect 5976 14116 5980 14172
rect 5980 14116 6036 14172
rect 6036 14116 6040 14172
rect 5976 14112 6040 14116
rect 6056 14172 6120 14176
rect 6056 14116 6060 14172
rect 6060 14116 6116 14172
rect 6116 14116 6120 14172
rect 6056 14112 6120 14116
rect 6136 14172 6200 14176
rect 6136 14116 6140 14172
rect 6140 14116 6196 14172
rect 6196 14116 6200 14172
rect 6136 14112 6200 14116
rect 10841 14172 10905 14176
rect 10841 14116 10845 14172
rect 10845 14116 10901 14172
rect 10901 14116 10905 14172
rect 10841 14112 10905 14116
rect 10921 14172 10985 14176
rect 10921 14116 10925 14172
rect 10925 14116 10981 14172
rect 10981 14116 10985 14172
rect 10921 14112 10985 14116
rect 11001 14172 11065 14176
rect 11001 14116 11005 14172
rect 11005 14116 11061 14172
rect 11061 14116 11065 14172
rect 11001 14112 11065 14116
rect 11081 14172 11145 14176
rect 11081 14116 11085 14172
rect 11085 14116 11141 14172
rect 11141 14116 11145 14172
rect 11081 14112 11145 14116
rect 15786 14172 15850 14176
rect 15786 14116 15790 14172
rect 15790 14116 15846 14172
rect 15846 14116 15850 14172
rect 15786 14112 15850 14116
rect 15866 14172 15930 14176
rect 15866 14116 15870 14172
rect 15870 14116 15926 14172
rect 15926 14116 15930 14172
rect 15866 14112 15930 14116
rect 15946 14172 16010 14176
rect 15946 14116 15950 14172
rect 15950 14116 16006 14172
rect 16006 14116 16010 14172
rect 15946 14112 16010 14116
rect 16026 14172 16090 14176
rect 16026 14116 16030 14172
rect 16030 14116 16086 14172
rect 16086 14116 16090 14172
rect 16026 14112 16090 14116
rect 20731 14172 20795 14176
rect 20731 14116 20735 14172
rect 20735 14116 20791 14172
rect 20791 14116 20795 14172
rect 20731 14112 20795 14116
rect 20811 14172 20875 14176
rect 20811 14116 20815 14172
rect 20815 14116 20871 14172
rect 20871 14116 20875 14172
rect 20811 14112 20875 14116
rect 20891 14172 20955 14176
rect 20891 14116 20895 14172
rect 20895 14116 20951 14172
rect 20951 14116 20955 14172
rect 20891 14112 20955 14116
rect 20971 14172 21035 14176
rect 20971 14116 20975 14172
rect 20975 14116 21031 14172
rect 21031 14116 21035 14172
rect 20971 14112 21035 14116
rect 3424 13628 3488 13632
rect 3424 13572 3428 13628
rect 3428 13572 3484 13628
rect 3484 13572 3488 13628
rect 3424 13568 3488 13572
rect 3504 13628 3568 13632
rect 3504 13572 3508 13628
rect 3508 13572 3564 13628
rect 3564 13572 3568 13628
rect 3504 13568 3568 13572
rect 3584 13628 3648 13632
rect 3584 13572 3588 13628
rect 3588 13572 3644 13628
rect 3644 13572 3648 13628
rect 3584 13568 3648 13572
rect 3664 13628 3728 13632
rect 3664 13572 3668 13628
rect 3668 13572 3724 13628
rect 3724 13572 3728 13628
rect 3664 13568 3728 13572
rect 8369 13628 8433 13632
rect 8369 13572 8373 13628
rect 8373 13572 8429 13628
rect 8429 13572 8433 13628
rect 8369 13568 8433 13572
rect 8449 13628 8513 13632
rect 8449 13572 8453 13628
rect 8453 13572 8509 13628
rect 8509 13572 8513 13628
rect 8449 13568 8513 13572
rect 8529 13628 8593 13632
rect 8529 13572 8533 13628
rect 8533 13572 8589 13628
rect 8589 13572 8593 13628
rect 8529 13568 8593 13572
rect 8609 13628 8673 13632
rect 8609 13572 8613 13628
rect 8613 13572 8669 13628
rect 8669 13572 8673 13628
rect 8609 13568 8673 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 13554 13628 13618 13632
rect 13554 13572 13558 13628
rect 13558 13572 13614 13628
rect 13614 13572 13618 13628
rect 13554 13568 13618 13572
rect 18259 13628 18323 13632
rect 18259 13572 18263 13628
rect 18263 13572 18319 13628
rect 18319 13572 18323 13628
rect 18259 13568 18323 13572
rect 18339 13628 18403 13632
rect 18339 13572 18343 13628
rect 18343 13572 18399 13628
rect 18399 13572 18403 13628
rect 18339 13568 18403 13572
rect 18419 13628 18483 13632
rect 18419 13572 18423 13628
rect 18423 13572 18479 13628
rect 18479 13572 18483 13628
rect 18419 13568 18483 13572
rect 18499 13628 18563 13632
rect 18499 13572 18503 13628
rect 18503 13572 18559 13628
rect 18559 13572 18563 13628
rect 18499 13568 18563 13572
rect 5896 13084 5960 13088
rect 5896 13028 5900 13084
rect 5900 13028 5956 13084
rect 5956 13028 5960 13084
rect 5896 13024 5960 13028
rect 5976 13084 6040 13088
rect 5976 13028 5980 13084
rect 5980 13028 6036 13084
rect 6036 13028 6040 13084
rect 5976 13024 6040 13028
rect 6056 13084 6120 13088
rect 6056 13028 6060 13084
rect 6060 13028 6116 13084
rect 6116 13028 6120 13084
rect 6056 13024 6120 13028
rect 6136 13084 6200 13088
rect 6136 13028 6140 13084
rect 6140 13028 6196 13084
rect 6196 13028 6200 13084
rect 6136 13024 6200 13028
rect 10841 13084 10905 13088
rect 10841 13028 10845 13084
rect 10845 13028 10901 13084
rect 10901 13028 10905 13084
rect 10841 13024 10905 13028
rect 10921 13084 10985 13088
rect 10921 13028 10925 13084
rect 10925 13028 10981 13084
rect 10981 13028 10985 13084
rect 10921 13024 10985 13028
rect 11001 13084 11065 13088
rect 11001 13028 11005 13084
rect 11005 13028 11061 13084
rect 11061 13028 11065 13084
rect 11001 13024 11065 13028
rect 11081 13084 11145 13088
rect 11081 13028 11085 13084
rect 11085 13028 11141 13084
rect 11141 13028 11145 13084
rect 11081 13024 11145 13028
rect 15786 13084 15850 13088
rect 15786 13028 15790 13084
rect 15790 13028 15846 13084
rect 15846 13028 15850 13084
rect 15786 13024 15850 13028
rect 15866 13084 15930 13088
rect 15866 13028 15870 13084
rect 15870 13028 15926 13084
rect 15926 13028 15930 13084
rect 15866 13024 15930 13028
rect 15946 13084 16010 13088
rect 15946 13028 15950 13084
rect 15950 13028 16006 13084
rect 16006 13028 16010 13084
rect 15946 13024 16010 13028
rect 16026 13084 16090 13088
rect 16026 13028 16030 13084
rect 16030 13028 16086 13084
rect 16086 13028 16090 13084
rect 16026 13024 16090 13028
rect 20731 13084 20795 13088
rect 20731 13028 20735 13084
rect 20735 13028 20791 13084
rect 20791 13028 20795 13084
rect 20731 13024 20795 13028
rect 20811 13084 20875 13088
rect 20811 13028 20815 13084
rect 20815 13028 20871 13084
rect 20871 13028 20875 13084
rect 20811 13024 20875 13028
rect 20891 13084 20955 13088
rect 20891 13028 20895 13084
rect 20895 13028 20951 13084
rect 20951 13028 20955 13084
rect 20891 13024 20955 13028
rect 20971 13084 21035 13088
rect 20971 13028 20975 13084
rect 20975 13028 21031 13084
rect 21031 13028 21035 13084
rect 20971 13024 21035 13028
rect 3424 12540 3488 12544
rect 3424 12484 3428 12540
rect 3428 12484 3484 12540
rect 3484 12484 3488 12540
rect 3424 12480 3488 12484
rect 3504 12540 3568 12544
rect 3504 12484 3508 12540
rect 3508 12484 3564 12540
rect 3564 12484 3568 12540
rect 3504 12480 3568 12484
rect 3584 12540 3648 12544
rect 3584 12484 3588 12540
rect 3588 12484 3644 12540
rect 3644 12484 3648 12540
rect 3584 12480 3648 12484
rect 3664 12540 3728 12544
rect 3664 12484 3668 12540
rect 3668 12484 3724 12540
rect 3724 12484 3728 12540
rect 3664 12480 3728 12484
rect 8369 12540 8433 12544
rect 8369 12484 8373 12540
rect 8373 12484 8429 12540
rect 8429 12484 8433 12540
rect 8369 12480 8433 12484
rect 8449 12540 8513 12544
rect 8449 12484 8453 12540
rect 8453 12484 8509 12540
rect 8509 12484 8513 12540
rect 8449 12480 8513 12484
rect 8529 12540 8593 12544
rect 8529 12484 8533 12540
rect 8533 12484 8589 12540
rect 8589 12484 8593 12540
rect 8529 12480 8593 12484
rect 8609 12540 8673 12544
rect 8609 12484 8613 12540
rect 8613 12484 8669 12540
rect 8669 12484 8673 12540
rect 8609 12480 8673 12484
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 13554 12540 13618 12544
rect 13554 12484 13558 12540
rect 13558 12484 13614 12540
rect 13614 12484 13618 12540
rect 13554 12480 13618 12484
rect 18259 12540 18323 12544
rect 18259 12484 18263 12540
rect 18263 12484 18319 12540
rect 18319 12484 18323 12540
rect 18259 12480 18323 12484
rect 18339 12540 18403 12544
rect 18339 12484 18343 12540
rect 18343 12484 18399 12540
rect 18399 12484 18403 12540
rect 18339 12480 18403 12484
rect 18419 12540 18483 12544
rect 18419 12484 18423 12540
rect 18423 12484 18479 12540
rect 18479 12484 18483 12540
rect 18419 12480 18483 12484
rect 18499 12540 18563 12544
rect 18499 12484 18503 12540
rect 18503 12484 18559 12540
rect 18559 12484 18563 12540
rect 18499 12480 18563 12484
rect 5896 11996 5960 12000
rect 5896 11940 5900 11996
rect 5900 11940 5956 11996
rect 5956 11940 5960 11996
rect 5896 11936 5960 11940
rect 5976 11996 6040 12000
rect 5976 11940 5980 11996
rect 5980 11940 6036 11996
rect 6036 11940 6040 11996
rect 5976 11936 6040 11940
rect 6056 11996 6120 12000
rect 6056 11940 6060 11996
rect 6060 11940 6116 11996
rect 6116 11940 6120 11996
rect 6056 11936 6120 11940
rect 6136 11996 6200 12000
rect 6136 11940 6140 11996
rect 6140 11940 6196 11996
rect 6196 11940 6200 11996
rect 6136 11936 6200 11940
rect 10841 11996 10905 12000
rect 10841 11940 10845 11996
rect 10845 11940 10901 11996
rect 10901 11940 10905 11996
rect 10841 11936 10905 11940
rect 10921 11996 10985 12000
rect 10921 11940 10925 11996
rect 10925 11940 10981 11996
rect 10981 11940 10985 11996
rect 10921 11936 10985 11940
rect 11001 11996 11065 12000
rect 11001 11940 11005 11996
rect 11005 11940 11061 11996
rect 11061 11940 11065 11996
rect 11001 11936 11065 11940
rect 11081 11996 11145 12000
rect 11081 11940 11085 11996
rect 11085 11940 11141 11996
rect 11141 11940 11145 11996
rect 11081 11936 11145 11940
rect 15786 11996 15850 12000
rect 15786 11940 15790 11996
rect 15790 11940 15846 11996
rect 15846 11940 15850 11996
rect 15786 11936 15850 11940
rect 15866 11996 15930 12000
rect 15866 11940 15870 11996
rect 15870 11940 15926 11996
rect 15926 11940 15930 11996
rect 15866 11936 15930 11940
rect 15946 11996 16010 12000
rect 15946 11940 15950 11996
rect 15950 11940 16006 11996
rect 16006 11940 16010 11996
rect 15946 11936 16010 11940
rect 16026 11996 16090 12000
rect 16026 11940 16030 11996
rect 16030 11940 16086 11996
rect 16086 11940 16090 11996
rect 16026 11936 16090 11940
rect 20731 11996 20795 12000
rect 20731 11940 20735 11996
rect 20735 11940 20791 11996
rect 20791 11940 20795 11996
rect 20731 11936 20795 11940
rect 20811 11996 20875 12000
rect 20811 11940 20815 11996
rect 20815 11940 20871 11996
rect 20871 11940 20875 11996
rect 20811 11936 20875 11940
rect 20891 11996 20955 12000
rect 20891 11940 20895 11996
rect 20895 11940 20951 11996
rect 20951 11940 20955 11996
rect 20891 11936 20955 11940
rect 20971 11996 21035 12000
rect 20971 11940 20975 11996
rect 20975 11940 21031 11996
rect 21031 11940 21035 11996
rect 20971 11936 21035 11940
rect 3424 11452 3488 11456
rect 3424 11396 3428 11452
rect 3428 11396 3484 11452
rect 3484 11396 3488 11452
rect 3424 11392 3488 11396
rect 3504 11452 3568 11456
rect 3504 11396 3508 11452
rect 3508 11396 3564 11452
rect 3564 11396 3568 11452
rect 3504 11392 3568 11396
rect 3584 11452 3648 11456
rect 3584 11396 3588 11452
rect 3588 11396 3644 11452
rect 3644 11396 3648 11452
rect 3584 11392 3648 11396
rect 3664 11452 3728 11456
rect 3664 11396 3668 11452
rect 3668 11396 3724 11452
rect 3724 11396 3728 11452
rect 3664 11392 3728 11396
rect 8369 11452 8433 11456
rect 8369 11396 8373 11452
rect 8373 11396 8429 11452
rect 8429 11396 8433 11452
rect 8369 11392 8433 11396
rect 8449 11452 8513 11456
rect 8449 11396 8453 11452
rect 8453 11396 8509 11452
rect 8509 11396 8513 11452
rect 8449 11392 8513 11396
rect 8529 11452 8593 11456
rect 8529 11396 8533 11452
rect 8533 11396 8589 11452
rect 8589 11396 8593 11452
rect 8529 11392 8593 11396
rect 8609 11452 8673 11456
rect 8609 11396 8613 11452
rect 8613 11396 8669 11452
rect 8669 11396 8673 11452
rect 8609 11392 8673 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 13554 11452 13618 11456
rect 13554 11396 13558 11452
rect 13558 11396 13614 11452
rect 13614 11396 13618 11452
rect 13554 11392 13618 11396
rect 18259 11452 18323 11456
rect 18259 11396 18263 11452
rect 18263 11396 18319 11452
rect 18319 11396 18323 11452
rect 18259 11392 18323 11396
rect 18339 11452 18403 11456
rect 18339 11396 18343 11452
rect 18343 11396 18399 11452
rect 18399 11396 18403 11452
rect 18339 11392 18403 11396
rect 18419 11452 18483 11456
rect 18419 11396 18423 11452
rect 18423 11396 18479 11452
rect 18479 11396 18483 11452
rect 18419 11392 18483 11396
rect 18499 11452 18563 11456
rect 18499 11396 18503 11452
rect 18503 11396 18559 11452
rect 18559 11396 18563 11452
rect 18499 11392 18563 11396
rect 5896 10908 5960 10912
rect 5896 10852 5900 10908
rect 5900 10852 5956 10908
rect 5956 10852 5960 10908
rect 5896 10848 5960 10852
rect 5976 10908 6040 10912
rect 5976 10852 5980 10908
rect 5980 10852 6036 10908
rect 6036 10852 6040 10908
rect 5976 10848 6040 10852
rect 6056 10908 6120 10912
rect 6056 10852 6060 10908
rect 6060 10852 6116 10908
rect 6116 10852 6120 10908
rect 6056 10848 6120 10852
rect 6136 10908 6200 10912
rect 6136 10852 6140 10908
rect 6140 10852 6196 10908
rect 6196 10852 6200 10908
rect 6136 10848 6200 10852
rect 10841 10908 10905 10912
rect 10841 10852 10845 10908
rect 10845 10852 10901 10908
rect 10901 10852 10905 10908
rect 10841 10848 10905 10852
rect 10921 10908 10985 10912
rect 10921 10852 10925 10908
rect 10925 10852 10981 10908
rect 10981 10852 10985 10908
rect 10921 10848 10985 10852
rect 11001 10908 11065 10912
rect 11001 10852 11005 10908
rect 11005 10852 11061 10908
rect 11061 10852 11065 10908
rect 11001 10848 11065 10852
rect 11081 10908 11145 10912
rect 11081 10852 11085 10908
rect 11085 10852 11141 10908
rect 11141 10852 11145 10908
rect 11081 10848 11145 10852
rect 15786 10908 15850 10912
rect 15786 10852 15790 10908
rect 15790 10852 15846 10908
rect 15846 10852 15850 10908
rect 15786 10848 15850 10852
rect 15866 10908 15930 10912
rect 15866 10852 15870 10908
rect 15870 10852 15926 10908
rect 15926 10852 15930 10908
rect 15866 10848 15930 10852
rect 15946 10908 16010 10912
rect 15946 10852 15950 10908
rect 15950 10852 16006 10908
rect 16006 10852 16010 10908
rect 15946 10848 16010 10852
rect 16026 10908 16090 10912
rect 16026 10852 16030 10908
rect 16030 10852 16086 10908
rect 16086 10852 16090 10908
rect 16026 10848 16090 10852
rect 20731 10908 20795 10912
rect 20731 10852 20735 10908
rect 20735 10852 20791 10908
rect 20791 10852 20795 10908
rect 20731 10848 20795 10852
rect 20811 10908 20875 10912
rect 20811 10852 20815 10908
rect 20815 10852 20871 10908
rect 20871 10852 20875 10908
rect 20811 10848 20875 10852
rect 20891 10908 20955 10912
rect 20891 10852 20895 10908
rect 20895 10852 20951 10908
rect 20951 10852 20955 10908
rect 20891 10848 20955 10852
rect 20971 10908 21035 10912
rect 20971 10852 20975 10908
rect 20975 10852 21031 10908
rect 21031 10852 21035 10908
rect 20971 10848 21035 10852
rect 3424 10364 3488 10368
rect 3424 10308 3428 10364
rect 3428 10308 3484 10364
rect 3484 10308 3488 10364
rect 3424 10304 3488 10308
rect 3504 10364 3568 10368
rect 3504 10308 3508 10364
rect 3508 10308 3564 10364
rect 3564 10308 3568 10364
rect 3504 10304 3568 10308
rect 3584 10364 3648 10368
rect 3584 10308 3588 10364
rect 3588 10308 3644 10364
rect 3644 10308 3648 10364
rect 3584 10304 3648 10308
rect 3664 10364 3728 10368
rect 3664 10308 3668 10364
rect 3668 10308 3724 10364
rect 3724 10308 3728 10364
rect 3664 10304 3728 10308
rect 8369 10364 8433 10368
rect 8369 10308 8373 10364
rect 8373 10308 8429 10364
rect 8429 10308 8433 10364
rect 8369 10304 8433 10308
rect 8449 10364 8513 10368
rect 8449 10308 8453 10364
rect 8453 10308 8509 10364
rect 8509 10308 8513 10364
rect 8449 10304 8513 10308
rect 8529 10364 8593 10368
rect 8529 10308 8533 10364
rect 8533 10308 8589 10364
rect 8589 10308 8593 10364
rect 8529 10304 8593 10308
rect 8609 10364 8673 10368
rect 8609 10308 8613 10364
rect 8613 10308 8669 10364
rect 8669 10308 8673 10364
rect 8609 10304 8673 10308
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 13554 10364 13618 10368
rect 13554 10308 13558 10364
rect 13558 10308 13614 10364
rect 13614 10308 13618 10364
rect 13554 10304 13618 10308
rect 18259 10364 18323 10368
rect 18259 10308 18263 10364
rect 18263 10308 18319 10364
rect 18319 10308 18323 10364
rect 18259 10304 18323 10308
rect 18339 10364 18403 10368
rect 18339 10308 18343 10364
rect 18343 10308 18399 10364
rect 18399 10308 18403 10364
rect 18339 10304 18403 10308
rect 18419 10364 18483 10368
rect 18419 10308 18423 10364
rect 18423 10308 18479 10364
rect 18479 10308 18483 10364
rect 18419 10304 18483 10308
rect 18499 10364 18563 10368
rect 18499 10308 18503 10364
rect 18503 10308 18559 10364
rect 18559 10308 18563 10364
rect 18499 10304 18563 10308
rect 5896 9820 5960 9824
rect 5896 9764 5900 9820
rect 5900 9764 5956 9820
rect 5956 9764 5960 9820
rect 5896 9760 5960 9764
rect 5976 9820 6040 9824
rect 5976 9764 5980 9820
rect 5980 9764 6036 9820
rect 6036 9764 6040 9820
rect 5976 9760 6040 9764
rect 6056 9820 6120 9824
rect 6056 9764 6060 9820
rect 6060 9764 6116 9820
rect 6116 9764 6120 9820
rect 6056 9760 6120 9764
rect 6136 9820 6200 9824
rect 6136 9764 6140 9820
rect 6140 9764 6196 9820
rect 6196 9764 6200 9820
rect 6136 9760 6200 9764
rect 10841 9820 10905 9824
rect 10841 9764 10845 9820
rect 10845 9764 10901 9820
rect 10901 9764 10905 9820
rect 10841 9760 10905 9764
rect 10921 9820 10985 9824
rect 10921 9764 10925 9820
rect 10925 9764 10981 9820
rect 10981 9764 10985 9820
rect 10921 9760 10985 9764
rect 11001 9820 11065 9824
rect 11001 9764 11005 9820
rect 11005 9764 11061 9820
rect 11061 9764 11065 9820
rect 11001 9760 11065 9764
rect 11081 9820 11145 9824
rect 11081 9764 11085 9820
rect 11085 9764 11141 9820
rect 11141 9764 11145 9820
rect 11081 9760 11145 9764
rect 15786 9820 15850 9824
rect 15786 9764 15790 9820
rect 15790 9764 15846 9820
rect 15846 9764 15850 9820
rect 15786 9760 15850 9764
rect 15866 9820 15930 9824
rect 15866 9764 15870 9820
rect 15870 9764 15926 9820
rect 15926 9764 15930 9820
rect 15866 9760 15930 9764
rect 15946 9820 16010 9824
rect 15946 9764 15950 9820
rect 15950 9764 16006 9820
rect 16006 9764 16010 9820
rect 15946 9760 16010 9764
rect 16026 9820 16090 9824
rect 16026 9764 16030 9820
rect 16030 9764 16086 9820
rect 16086 9764 16090 9820
rect 16026 9760 16090 9764
rect 20731 9820 20795 9824
rect 20731 9764 20735 9820
rect 20735 9764 20791 9820
rect 20791 9764 20795 9820
rect 20731 9760 20795 9764
rect 20811 9820 20875 9824
rect 20811 9764 20815 9820
rect 20815 9764 20871 9820
rect 20871 9764 20875 9820
rect 20811 9760 20875 9764
rect 20891 9820 20955 9824
rect 20891 9764 20895 9820
rect 20895 9764 20951 9820
rect 20951 9764 20955 9820
rect 20891 9760 20955 9764
rect 20971 9820 21035 9824
rect 20971 9764 20975 9820
rect 20975 9764 21031 9820
rect 21031 9764 21035 9820
rect 20971 9760 21035 9764
rect 3424 9276 3488 9280
rect 3424 9220 3428 9276
rect 3428 9220 3484 9276
rect 3484 9220 3488 9276
rect 3424 9216 3488 9220
rect 3504 9276 3568 9280
rect 3504 9220 3508 9276
rect 3508 9220 3564 9276
rect 3564 9220 3568 9276
rect 3504 9216 3568 9220
rect 3584 9276 3648 9280
rect 3584 9220 3588 9276
rect 3588 9220 3644 9276
rect 3644 9220 3648 9276
rect 3584 9216 3648 9220
rect 3664 9276 3728 9280
rect 3664 9220 3668 9276
rect 3668 9220 3724 9276
rect 3724 9220 3728 9276
rect 3664 9216 3728 9220
rect 8369 9276 8433 9280
rect 8369 9220 8373 9276
rect 8373 9220 8429 9276
rect 8429 9220 8433 9276
rect 8369 9216 8433 9220
rect 8449 9276 8513 9280
rect 8449 9220 8453 9276
rect 8453 9220 8509 9276
rect 8509 9220 8513 9276
rect 8449 9216 8513 9220
rect 8529 9276 8593 9280
rect 8529 9220 8533 9276
rect 8533 9220 8589 9276
rect 8589 9220 8593 9276
rect 8529 9216 8593 9220
rect 8609 9276 8673 9280
rect 8609 9220 8613 9276
rect 8613 9220 8669 9276
rect 8669 9220 8673 9276
rect 8609 9216 8673 9220
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 13554 9276 13618 9280
rect 13554 9220 13558 9276
rect 13558 9220 13614 9276
rect 13614 9220 13618 9276
rect 13554 9216 13618 9220
rect 18259 9276 18323 9280
rect 18259 9220 18263 9276
rect 18263 9220 18319 9276
rect 18319 9220 18323 9276
rect 18259 9216 18323 9220
rect 18339 9276 18403 9280
rect 18339 9220 18343 9276
rect 18343 9220 18399 9276
rect 18399 9220 18403 9276
rect 18339 9216 18403 9220
rect 18419 9276 18483 9280
rect 18419 9220 18423 9276
rect 18423 9220 18479 9276
rect 18479 9220 18483 9276
rect 18419 9216 18483 9220
rect 18499 9276 18563 9280
rect 18499 9220 18503 9276
rect 18503 9220 18559 9276
rect 18559 9220 18563 9276
rect 18499 9216 18563 9220
rect 5896 8732 5960 8736
rect 5896 8676 5900 8732
rect 5900 8676 5956 8732
rect 5956 8676 5960 8732
rect 5896 8672 5960 8676
rect 5976 8732 6040 8736
rect 5976 8676 5980 8732
rect 5980 8676 6036 8732
rect 6036 8676 6040 8732
rect 5976 8672 6040 8676
rect 6056 8732 6120 8736
rect 6056 8676 6060 8732
rect 6060 8676 6116 8732
rect 6116 8676 6120 8732
rect 6056 8672 6120 8676
rect 6136 8732 6200 8736
rect 6136 8676 6140 8732
rect 6140 8676 6196 8732
rect 6196 8676 6200 8732
rect 6136 8672 6200 8676
rect 10841 8732 10905 8736
rect 10841 8676 10845 8732
rect 10845 8676 10901 8732
rect 10901 8676 10905 8732
rect 10841 8672 10905 8676
rect 10921 8732 10985 8736
rect 10921 8676 10925 8732
rect 10925 8676 10981 8732
rect 10981 8676 10985 8732
rect 10921 8672 10985 8676
rect 11001 8732 11065 8736
rect 11001 8676 11005 8732
rect 11005 8676 11061 8732
rect 11061 8676 11065 8732
rect 11001 8672 11065 8676
rect 11081 8732 11145 8736
rect 11081 8676 11085 8732
rect 11085 8676 11141 8732
rect 11141 8676 11145 8732
rect 11081 8672 11145 8676
rect 15786 8732 15850 8736
rect 15786 8676 15790 8732
rect 15790 8676 15846 8732
rect 15846 8676 15850 8732
rect 15786 8672 15850 8676
rect 15866 8732 15930 8736
rect 15866 8676 15870 8732
rect 15870 8676 15926 8732
rect 15926 8676 15930 8732
rect 15866 8672 15930 8676
rect 15946 8732 16010 8736
rect 15946 8676 15950 8732
rect 15950 8676 16006 8732
rect 16006 8676 16010 8732
rect 15946 8672 16010 8676
rect 16026 8732 16090 8736
rect 16026 8676 16030 8732
rect 16030 8676 16086 8732
rect 16086 8676 16090 8732
rect 16026 8672 16090 8676
rect 20731 8732 20795 8736
rect 20731 8676 20735 8732
rect 20735 8676 20791 8732
rect 20791 8676 20795 8732
rect 20731 8672 20795 8676
rect 20811 8732 20875 8736
rect 20811 8676 20815 8732
rect 20815 8676 20871 8732
rect 20871 8676 20875 8732
rect 20811 8672 20875 8676
rect 20891 8732 20955 8736
rect 20891 8676 20895 8732
rect 20895 8676 20951 8732
rect 20951 8676 20955 8732
rect 20891 8672 20955 8676
rect 20971 8732 21035 8736
rect 20971 8676 20975 8732
rect 20975 8676 21031 8732
rect 21031 8676 21035 8732
rect 20971 8672 21035 8676
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 3584 8188 3648 8192
rect 3584 8132 3588 8188
rect 3588 8132 3644 8188
rect 3644 8132 3648 8188
rect 3584 8128 3648 8132
rect 3664 8188 3728 8192
rect 3664 8132 3668 8188
rect 3668 8132 3724 8188
rect 3724 8132 3728 8188
rect 3664 8128 3728 8132
rect 8369 8188 8433 8192
rect 8369 8132 8373 8188
rect 8373 8132 8429 8188
rect 8429 8132 8433 8188
rect 8369 8128 8433 8132
rect 8449 8188 8513 8192
rect 8449 8132 8453 8188
rect 8453 8132 8509 8188
rect 8509 8132 8513 8188
rect 8449 8128 8513 8132
rect 8529 8188 8593 8192
rect 8529 8132 8533 8188
rect 8533 8132 8589 8188
rect 8589 8132 8593 8188
rect 8529 8128 8593 8132
rect 8609 8188 8673 8192
rect 8609 8132 8613 8188
rect 8613 8132 8669 8188
rect 8669 8132 8673 8188
rect 8609 8128 8673 8132
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 13554 8188 13618 8192
rect 13554 8132 13558 8188
rect 13558 8132 13614 8188
rect 13614 8132 13618 8188
rect 13554 8128 13618 8132
rect 18259 8188 18323 8192
rect 18259 8132 18263 8188
rect 18263 8132 18319 8188
rect 18319 8132 18323 8188
rect 18259 8128 18323 8132
rect 18339 8188 18403 8192
rect 18339 8132 18343 8188
rect 18343 8132 18399 8188
rect 18399 8132 18403 8188
rect 18339 8128 18403 8132
rect 18419 8188 18483 8192
rect 18419 8132 18423 8188
rect 18423 8132 18479 8188
rect 18479 8132 18483 8188
rect 18419 8128 18483 8132
rect 18499 8188 18563 8192
rect 18499 8132 18503 8188
rect 18503 8132 18559 8188
rect 18559 8132 18563 8188
rect 18499 8128 18563 8132
rect 5896 7644 5960 7648
rect 5896 7588 5900 7644
rect 5900 7588 5956 7644
rect 5956 7588 5960 7644
rect 5896 7584 5960 7588
rect 5976 7644 6040 7648
rect 5976 7588 5980 7644
rect 5980 7588 6036 7644
rect 6036 7588 6040 7644
rect 5976 7584 6040 7588
rect 6056 7644 6120 7648
rect 6056 7588 6060 7644
rect 6060 7588 6116 7644
rect 6116 7588 6120 7644
rect 6056 7584 6120 7588
rect 6136 7644 6200 7648
rect 6136 7588 6140 7644
rect 6140 7588 6196 7644
rect 6196 7588 6200 7644
rect 6136 7584 6200 7588
rect 10841 7644 10905 7648
rect 10841 7588 10845 7644
rect 10845 7588 10901 7644
rect 10901 7588 10905 7644
rect 10841 7584 10905 7588
rect 10921 7644 10985 7648
rect 10921 7588 10925 7644
rect 10925 7588 10981 7644
rect 10981 7588 10985 7644
rect 10921 7584 10985 7588
rect 11001 7644 11065 7648
rect 11001 7588 11005 7644
rect 11005 7588 11061 7644
rect 11061 7588 11065 7644
rect 11001 7584 11065 7588
rect 11081 7644 11145 7648
rect 11081 7588 11085 7644
rect 11085 7588 11141 7644
rect 11141 7588 11145 7644
rect 11081 7584 11145 7588
rect 15786 7644 15850 7648
rect 15786 7588 15790 7644
rect 15790 7588 15846 7644
rect 15846 7588 15850 7644
rect 15786 7584 15850 7588
rect 15866 7644 15930 7648
rect 15866 7588 15870 7644
rect 15870 7588 15926 7644
rect 15926 7588 15930 7644
rect 15866 7584 15930 7588
rect 15946 7644 16010 7648
rect 15946 7588 15950 7644
rect 15950 7588 16006 7644
rect 16006 7588 16010 7644
rect 15946 7584 16010 7588
rect 16026 7644 16090 7648
rect 16026 7588 16030 7644
rect 16030 7588 16086 7644
rect 16086 7588 16090 7644
rect 16026 7584 16090 7588
rect 20731 7644 20795 7648
rect 20731 7588 20735 7644
rect 20735 7588 20791 7644
rect 20791 7588 20795 7644
rect 20731 7584 20795 7588
rect 20811 7644 20875 7648
rect 20811 7588 20815 7644
rect 20815 7588 20871 7644
rect 20871 7588 20875 7644
rect 20811 7584 20875 7588
rect 20891 7644 20955 7648
rect 20891 7588 20895 7644
rect 20895 7588 20951 7644
rect 20951 7588 20955 7644
rect 20891 7584 20955 7588
rect 20971 7644 21035 7648
rect 20971 7588 20975 7644
rect 20975 7588 21031 7644
rect 21031 7588 21035 7644
rect 20971 7584 21035 7588
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 3584 7100 3648 7104
rect 3584 7044 3588 7100
rect 3588 7044 3644 7100
rect 3644 7044 3648 7100
rect 3584 7040 3648 7044
rect 3664 7100 3728 7104
rect 3664 7044 3668 7100
rect 3668 7044 3724 7100
rect 3724 7044 3728 7100
rect 3664 7040 3728 7044
rect 8369 7100 8433 7104
rect 8369 7044 8373 7100
rect 8373 7044 8429 7100
rect 8429 7044 8433 7100
rect 8369 7040 8433 7044
rect 8449 7100 8513 7104
rect 8449 7044 8453 7100
rect 8453 7044 8509 7100
rect 8509 7044 8513 7100
rect 8449 7040 8513 7044
rect 8529 7100 8593 7104
rect 8529 7044 8533 7100
rect 8533 7044 8589 7100
rect 8589 7044 8593 7100
rect 8529 7040 8593 7044
rect 8609 7100 8673 7104
rect 8609 7044 8613 7100
rect 8613 7044 8669 7100
rect 8669 7044 8673 7100
rect 8609 7040 8673 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 13554 7100 13618 7104
rect 13554 7044 13558 7100
rect 13558 7044 13614 7100
rect 13614 7044 13618 7100
rect 13554 7040 13618 7044
rect 18259 7100 18323 7104
rect 18259 7044 18263 7100
rect 18263 7044 18319 7100
rect 18319 7044 18323 7100
rect 18259 7040 18323 7044
rect 18339 7100 18403 7104
rect 18339 7044 18343 7100
rect 18343 7044 18399 7100
rect 18399 7044 18403 7100
rect 18339 7040 18403 7044
rect 18419 7100 18483 7104
rect 18419 7044 18423 7100
rect 18423 7044 18479 7100
rect 18479 7044 18483 7100
rect 18419 7040 18483 7044
rect 18499 7100 18563 7104
rect 18499 7044 18503 7100
rect 18503 7044 18559 7100
rect 18559 7044 18563 7100
rect 18499 7040 18563 7044
rect 5896 6556 5960 6560
rect 5896 6500 5900 6556
rect 5900 6500 5956 6556
rect 5956 6500 5960 6556
rect 5896 6496 5960 6500
rect 5976 6556 6040 6560
rect 5976 6500 5980 6556
rect 5980 6500 6036 6556
rect 6036 6500 6040 6556
rect 5976 6496 6040 6500
rect 6056 6556 6120 6560
rect 6056 6500 6060 6556
rect 6060 6500 6116 6556
rect 6116 6500 6120 6556
rect 6056 6496 6120 6500
rect 6136 6556 6200 6560
rect 6136 6500 6140 6556
rect 6140 6500 6196 6556
rect 6196 6500 6200 6556
rect 6136 6496 6200 6500
rect 10841 6556 10905 6560
rect 10841 6500 10845 6556
rect 10845 6500 10901 6556
rect 10901 6500 10905 6556
rect 10841 6496 10905 6500
rect 10921 6556 10985 6560
rect 10921 6500 10925 6556
rect 10925 6500 10981 6556
rect 10981 6500 10985 6556
rect 10921 6496 10985 6500
rect 11001 6556 11065 6560
rect 11001 6500 11005 6556
rect 11005 6500 11061 6556
rect 11061 6500 11065 6556
rect 11001 6496 11065 6500
rect 11081 6556 11145 6560
rect 11081 6500 11085 6556
rect 11085 6500 11141 6556
rect 11141 6500 11145 6556
rect 11081 6496 11145 6500
rect 15786 6556 15850 6560
rect 15786 6500 15790 6556
rect 15790 6500 15846 6556
rect 15846 6500 15850 6556
rect 15786 6496 15850 6500
rect 15866 6556 15930 6560
rect 15866 6500 15870 6556
rect 15870 6500 15926 6556
rect 15926 6500 15930 6556
rect 15866 6496 15930 6500
rect 15946 6556 16010 6560
rect 15946 6500 15950 6556
rect 15950 6500 16006 6556
rect 16006 6500 16010 6556
rect 15946 6496 16010 6500
rect 16026 6556 16090 6560
rect 16026 6500 16030 6556
rect 16030 6500 16086 6556
rect 16086 6500 16090 6556
rect 16026 6496 16090 6500
rect 20731 6556 20795 6560
rect 20731 6500 20735 6556
rect 20735 6500 20791 6556
rect 20791 6500 20795 6556
rect 20731 6496 20795 6500
rect 20811 6556 20875 6560
rect 20811 6500 20815 6556
rect 20815 6500 20871 6556
rect 20871 6500 20875 6556
rect 20811 6496 20875 6500
rect 20891 6556 20955 6560
rect 20891 6500 20895 6556
rect 20895 6500 20951 6556
rect 20951 6500 20955 6556
rect 20891 6496 20955 6500
rect 20971 6556 21035 6560
rect 20971 6500 20975 6556
rect 20975 6500 21031 6556
rect 21031 6500 21035 6556
rect 20971 6496 21035 6500
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 3584 6012 3648 6016
rect 3584 5956 3588 6012
rect 3588 5956 3644 6012
rect 3644 5956 3648 6012
rect 3584 5952 3648 5956
rect 3664 6012 3728 6016
rect 3664 5956 3668 6012
rect 3668 5956 3724 6012
rect 3724 5956 3728 6012
rect 3664 5952 3728 5956
rect 8369 6012 8433 6016
rect 8369 5956 8373 6012
rect 8373 5956 8429 6012
rect 8429 5956 8433 6012
rect 8369 5952 8433 5956
rect 8449 6012 8513 6016
rect 8449 5956 8453 6012
rect 8453 5956 8509 6012
rect 8509 5956 8513 6012
rect 8449 5952 8513 5956
rect 8529 6012 8593 6016
rect 8529 5956 8533 6012
rect 8533 5956 8589 6012
rect 8589 5956 8593 6012
rect 8529 5952 8593 5956
rect 8609 6012 8673 6016
rect 8609 5956 8613 6012
rect 8613 5956 8669 6012
rect 8669 5956 8673 6012
rect 8609 5952 8673 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 13554 6012 13618 6016
rect 13554 5956 13558 6012
rect 13558 5956 13614 6012
rect 13614 5956 13618 6012
rect 13554 5952 13618 5956
rect 18259 6012 18323 6016
rect 18259 5956 18263 6012
rect 18263 5956 18319 6012
rect 18319 5956 18323 6012
rect 18259 5952 18323 5956
rect 18339 6012 18403 6016
rect 18339 5956 18343 6012
rect 18343 5956 18399 6012
rect 18399 5956 18403 6012
rect 18339 5952 18403 5956
rect 18419 6012 18483 6016
rect 18419 5956 18423 6012
rect 18423 5956 18479 6012
rect 18479 5956 18483 6012
rect 18419 5952 18483 5956
rect 18499 6012 18563 6016
rect 18499 5956 18503 6012
rect 18503 5956 18559 6012
rect 18559 5956 18563 6012
rect 18499 5952 18563 5956
rect 5896 5468 5960 5472
rect 5896 5412 5900 5468
rect 5900 5412 5956 5468
rect 5956 5412 5960 5468
rect 5896 5408 5960 5412
rect 5976 5468 6040 5472
rect 5976 5412 5980 5468
rect 5980 5412 6036 5468
rect 6036 5412 6040 5468
rect 5976 5408 6040 5412
rect 6056 5468 6120 5472
rect 6056 5412 6060 5468
rect 6060 5412 6116 5468
rect 6116 5412 6120 5468
rect 6056 5408 6120 5412
rect 6136 5468 6200 5472
rect 6136 5412 6140 5468
rect 6140 5412 6196 5468
rect 6196 5412 6200 5468
rect 6136 5408 6200 5412
rect 10841 5468 10905 5472
rect 10841 5412 10845 5468
rect 10845 5412 10901 5468
rect 10901 5412 10905 5468
rect 10841 5408 10905 5412
rect 10921 5468 10985 5472
rect 10921 5412 10925 5468
rect 10925 5412 10981 5468
rect 10981 5412 10985 5468
rect 10921 5408 10985 5412
rect 11001 5468 11065 5472
rect 11001 5412 11005 5468
rect 11005 5412 11061 5468
rect 11061 5412 11065 5468
rect 11001 5408 11065 5412
rect 11081 5468 11145 5472
rect 11081 5412 11085 5468
rect 11085 5412 11141 5468
rect 11141 5412 11145 5468
rect 11081 5408 11145 5412
rect 15786 5468 15850 5472
rect 15786 5412 15790 5468
rect 15790 5412 15846 5468
rect 15846 5412 15850 5468
rect 15786 5408 15850 5412
rect 15866 5468 15930 5472
rect 15866 5412 15870 5468
rect 15870 5412 15926 5468
rect 15926 5412 15930 5468
rect 15866 5408 15930 5412
rect 15946 5468 16010 5472
rect 15946 5412 15950 5468
rect 15950 5412 16006 5468
rect 16006 5412 16010 5468
rect 15946 5408 16010 5412
rect 16026 5468 16090 5472
rect 16026 5412 16030 5468
rect 16030 5412 16086 5468
rect 16086 5412 16090 5468
rect 16026 5408 16090 5412
rect 20731 5468 20795 5472
rect 20731 5412 20735 5468
rect 20735 5412 20791 5468
rect 20791 5412 20795 5468
rect 20731 5408 20795 5412
rect 20811 5468 20875 5472
rect 20811 5412 20815 5468
rect 20815 5412 20871 5468
rect 20871 5412 20875 5468
rect 20811 5408 20875 5412
rect 20891 5468 20955 5472
rect 20891 5412 20895 5468
rect 20895 5412 20951 5468
rect 20951 5412 20955 5468
rect 20891 5408 20955 5412
rect 20971 5468 21035 5472
rect 20971 5412 20975 5468
rect 20975 5412 21031 5468
rect 21031 5412 21035 5468
rect 20971 5408 21035 5412
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 3584 4924 3648 4928
rect 3584 4868 3588 4924
rect 3588 4868 3644 4924
rect 3644 4868 3648 4924
rect 3584 4864 3648 4868
rect 3664 4924 3728 4928
rect 3664 4868 3668 4924
rect 3668 4868 3724 4924
rect 3724 4868 3728 4924
rect 3664 4864 3728 4868
rect 8369 4924 8433 4928
rect 8369 4868 8373 4924
rect 8373 4868 8429 4924
rect 8429 4868 8433 4924
rect 8369 4864 8433 4868
rect 8449 4924 8513 4928
rect 8449 4868 8453 4924
rect 8453 4868 8509 4924
rect 8509 4868 8513 4924
rect 8449 4864 8513 4868
rect 8529 4924 8593 4928
rect 8529 4868 8533 4924
rect 8533 4868 8589 4924
rect 8589 4868 8593 4924
rect 8529 4864 8593 4868
rect 8609 4924 8673 4928
rect 8609 4868 8613 4924
rect 8613 4868 8669 4924
rect 8669 4868 8673 4924
rect 8609 4864 8673 4868
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 13554 4924 13618 4928
rect 13554 4868 13558 4924
rect 13558 4868 13614 4924
rect 13614 4868 13618 4924
rect 13554 4864 13618 4868
rect 18259 4924 18323 4928
rect 18259 4868 18263 4924
rect 18263 4868 18319 4924
rect 18319 4868 18323 4924
rect 18259 4864 18323 4868
rect 18339 4924 18403 4928
rect 18339 4868 18343 4924
rect 18343 4868 18399 4924
rect 18399 4868 18403 4924
rect 18339 4864 18403 4868
rect 18419 4924 18483 4928
rect 18419 4868 18423 4924
rect 18423 4868 18479 4924
rect 18479 4868 18483 4924
rect 18419 4864 18483 4868
rect 18499 4924 18563 4928
rect 18499 4868 18503 4924
rect 18503 4868 18559 4924
rect 18559 4868 18563 4924
rect 18499 4864 18563 4868
rect 5896 4380 5960 4384
rect 5896 4324 5900 4380
rect 5900 4324 5956 4380
rect 5956 4324 5960 4380
rect 5896 4320 5960 4324
rect 5976 4380 6040 4384
rect 5976 4324 5980 4380
rect 5980 4324 6036 4380
rect 6036 4324 6040 4380
rect 5976 4320 6040 4324
rect 6056 4380 6120 4384
rect 6056 4324 6060 4380
rect 6060 4324 6116 4380
rect 6116 4324 6120 4380
rect 6056 4320 6120 4324
rect 6136 4380 6200 4384
rect 6136 4324 6140 4380
rect 6140 4324 6196 4380
rect 6196 4324 6200 4380
rect 6136 4320 6200 4324
rect 10841 4380 10905 4384
rect 10841 4324 10845 4380
rect 10845 4324 10901 4380
rect 10901 4324 10905 4380
rect 10841 4320 10905 4324
rect 10921 4380 10985 4384
rect 10921 4324 10925 4380
rect 10925 4324 10981 4380
rect 10981 4324 10985 4380
rect 10921 4320 10985 4324
rect 11001 4380 11065 4384
rect 11001 4324 11005 4380
rect 11005 4324 11061 4380
rect 11061 4324 11065 4380
rect 11001 4320 11065 4324
rect 11081 4380 11145 4384
rect 11081 4324 11085 4380
rect 11085 4324 11141 4380
rect 11141 4324 11145 4380
rect 11081 4320 11145 4324
rect 15786 4380 15850 4384
rect 15786 4324 15790 4380
rect 15790 4324 15846 4380
rect 15846 4324 15850 4380
rect 15786 4320 15850 4324
rect 15866 4380 15930 4384
rect 15866 4324 15870 4380
rect 15870 4324 15926 4380
rect 15926 4324 15930 4380
rect 15866 4320 15930 4324
rect 15946 4380 16010 4384
rect 15946 4324 15950 4380
rect 15950 4324 16006 4380
rect 16006 4324 16010 4380
rect 15946 4320 16010 4324
rect 16026 4380 16090 4384
rect 16026 4324 16030 4380
rect 16030 4324 16086 4380
rect 16086 4324 16090 4380
rect 16026 4320 16090 4324
rect 20731 4380 20795 4384
rect 20731 4324 20735 4380
rect 20735 4324 20791 4380
rect 20791 4324 20795 4380
rect 20731 4320 20795 4324
rect 20811 4380 20875 4384
rect 20811 4324 20815 4380
rect 20815 4324 20871 4380
rect 20871 4324 20875 4380
rect 20811 4320 20875 4324
rect 20891 4380 20955 4384
rect 20891 4324 20895 4380
rect 20895 4324 20951 4380
rect 20951 4324 20955 4380
rect 20891 4320 20955 4324
rect 20971 4380 21035 4384
rect 20971 4324 20975 4380
rect 20975 4324 21031 4380
rect 21031 4324 21035 4380
rect 20971 4320 21035 4324
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 3584 3836 3648 3840
rect 3584 3780 3588 3836
rect 3588 3780 3644 3836
rect 3644 3780 3648 3836
rect 3584 3776 3648 3780
rect 3664 3836 3728 3840
rect 3664 3780 3668 3836
rect 3668 3780 3724 3836
rect 3724 3780 3728 3836
rect 3664 3776 3728 3780
rect 8369 3836 8433 3840
rect 8369 3780 8373 3836
rect 8373 3780 8429 3836
rect 8429 3780 8433 3836
rect 8369 3776 8433 3780
rect 8449 3836 8513 3840
rect 8449 3780 8453 3836
rect 8453 3780 8509 3836
rect 8509 3780 8513 3836
rect 8449 3776 8513 3780
rect 8529 3836 8593 3840
rect 8529 3780 8533 3836
rect 8533 3780 8589 3836
rect 8589 3780 8593 3836
rect 8529 3776 8593 3780
rect 8609 3836 8673 3840
rect 8609 3780 8613 3836
rect 8613 3780 8669 3836
rect 8669 3780 8673 3836
rect 8609 3776 8673 3780
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 13554 3836 13618 3840
rect 13554 3780 13558 3836
rect 13558 3780 13614 3836
rect 13614 3780 13618 3836
rect 13554 3776 13618 3780
rect 18259 3836 18323 3840
rect 18259 3780 18263 3836
rect 18263 3780 18319 3836
rect 18319 3780 18323 3836
rect 18259 3776 18323 3780
rect 18339 3836 18403 3840
rect 18339 3780 18343 3836
rect 18343 3780 18399 3836
rect 18399 3780 18403 3836
rect 18339 3776 18403 3780
rect 18419 3836 18483 3840
rect 18419 3780 18423 3836
rect 18423 3780 18479 3836
rect 18479 3780 18483 3836
rect 18419 3776 18483 3780
rect 18499 3836 18563 3840
rect 18499 3780 18503 3836
rect 18503 3780 18559 3836
rect 18559 3780 18563 3836
rect 18499 3776 18563 3780
rect 5896 3292 5960 3296
rect 5896 3236 5900 3292
rect 5900 3236 5956 3292
rect 5956 3236 5960 3292
rect 5896 3232 5960 3236
rect 5976 3292 6040 3296
rect 5976 3236 5980 3292
rect 5980 3236 6036 3292
rect 6036 3236 6040 3292
rect 5976 3232 6040 3236
rect 6056 3292 6120 3296
rect 6056 3236 6060 3292
rect 6060 3236 6116 3292
rect 6116 3236 6120 3292
rect 6056 3232 6120 3236
rect 6136 3292 6200 3296
rect 6136 3236 6140 3292
rect 6140 3236 6196 3292
rect 6196 3236 6200 3292
rect 6136 3232 6200 3236
rect 10841 3292 10905 3296
rect 10841 3236 10845 3292
rect 10845 3236 10901 3292
rect 10901 3236 10905 3292
rect 10841 3232 10905 3236
rect 10921 3292 10985 3296
rect 10921 3236 10925 3292
rect 10925 3236 10981 3292
rect 10981 3236 10985 3292
rect 10921 3232 10985 3236
rect 11001 3292 11065 3296
rect 11001 3236 11005 3292
rect 11005 3236 11061 3292
rect 11061 3236 11065 3292
rect 11001 3232 11065 3236
rect 11081 3292 11145 3296
rect 11081 3236 11085 3292
rect 11085 3236 11141 3292
rect 11141 3236 11145 3292
rect 11081 3232 11145 3236
rect 15786 3292 15850 3296
rect 15786 3236 15790 3292
rect 15790 3236 15846 3292
rect 15846 3236 15850 3292
rect 15786 3232 15850 3236
rect 15866 3292 15930 3296
rect 15866 3236 15870 3292
rect 15870 3236 15926 3292
rect 15926 3236 15930 3292
rect 15866 3232 15930 3236
rect 15946 3292 16010 3296
rect 15946 3236 15950 3292
rect 15950 3236 16006 3292
rect 16006 3236 16010 3292
rect 15946 3232 16010 3236
rect 16026 3292 16090 3296
rect 16026 3236 16030 3292
rect 16030 3236 16086 3292
rect 16086 3236 16090 3292
rect 16026 3232 16090 3236
rect 20731 3292 20795 3296
rect 20731 3236 20735 3292
rect 20735 3236 20791 3292
rect 20791 3236 20795 3292
rect 20731 3232 20795 3236
rect 20811 3292 20875 3296
rect 20811 3236 20815 3292
rect 20815 3236 20871 3292
rect 20871 3236 20875 3292
rect 20811 3232 20875 3236
rect 20891 3292 20955 3296
rect 20891 3236 20895 3292
rect 20895 3236 20951 3292
rect 20951 3236 20955 3292
rect 20891 3232 20955 3236
rect 20971 3292 21035 3296
rect 20971 3236 20975 3292
rect 20975 3236 21031 3292
rect 21031 3236 21035 3292
rect 20971 3232 21035 3236
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 3584 2748 3648 2752
rect 3584 2692 3588 2748
rect 3588 2692 3644 2748
rect 3644 2692 3648 2748
rect 3584 2688 3648 2692
rect 3664 2748 3728 2752
rect 3664 2692 3668 2748
rect 3668 2692 3724 2748
rect 3724 2692 3728 2748
rect 3664 2688 3728 2692
rect 8369 2748 8433 2752
rect 8369 2692 8373 2748
rect 8373 2692 8429 2748
rect 8429 2692 8433 2748
rect 8369 2688 8433 2692
rect 8449 2748 8513 2752
rect 8449 2692 8453 2748
rect 8453 2692 8509 2748
rect 8509 2692 8513 2748
rect 8449 2688 8513 2692
rect 8529 2748 8593 2752
rect 8529 2692 8533 2748
rect 8533 2692 8589 2748
rect 8589 2692 8593 2748
rect 8529 2688 8593 2692
rect 8609 2748 8673 2752
rect 8609 2692 8613 2748
rect 8613 2692 8669 2748
rect 8669 2692 8673 2748
rect 8609 2688 8673 2692
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 13554 2748 13618 2752
rect 13554 2692 13558 2748
rect 13558 2692 13614 2748
rect 13614 2692 13618 2748
rect 13554 2688 13618 2692
rect 18259 2748 18323 2752
rect 18259 2692 18263 2748
rect 18263 2692 18319 2748
rect 18319 2692 18323 2748
rect 18259 2688 18323 2692
rect 18339 2748 18403 2752
rect 18339 2692 18343 2748
rect 18343 2692 18399 2748
rect 18399 2692 18403 2748
rect 18339 2688 18403 2692
rect 18419 2748 18483 2752
rect 18419 2692 18423 2748
rect 18423 2692 18479 2748
rect 18479 2692 18483 2748
rect 18419 2688 18483 2692
rect 18499 2748 18563 2752
rect 18499 2692 18503 2748
rect 18503 2692 18559 2748
rect 18559 2692 18563 2748
rect 18499 2688 18563 2692
rect 5896 2204 5960 2208
rect 5896 2148 5900 2204
rect 5900 2148 5956 2204
rect 5956 2148 5960 2204
rect 5896 2144 5960 2148
rect 5976 2204 6040 2208
rect 5976 2148 5980 2204
rect 5980 2148 6036 2204
rect 6036 2148 6040 2204
rect 5976 2144 6040 2148
rect 6056 2204 6120 2208
rect 6056 2148 6060 2204
rect 6060 2148 6116 2204
rect 6116 2148 6120 2204
rect 6056 2144 6120 2148
rect 6136 2204 6200 2208
rect 6136 2148 6140 2204
rect 6140 2148 6196 2204
rect 6196 2148 6200 2204
rect 6136 2144 6200 2148
rect 10841 2204 10905 2208
rect 10841 2148 10845 2204
rect 10845 2148 10901 2204
rect 10901 2148 10905 2204
rect 10841 2144 10905 2148
rect 10921 2204 10985 2208
rect 10921 2148 10925 2204
rect 10925 2148 10981 2204
rect 10981 2148 10985 2204
rect 10921 2144 10985 2148
rect 11001 2204 11065 2208
rect 11001 2148 11005 2204
rect 11005 2148 11061 2204
rect 11061 2148 11065 2204
rect 11001 2144 11065 2148
rect 11081 2204 11145 2208
rect 11081 2148 11085 2204
rect 11085 2148 11141 2204
rect 11141 2148 11145 2204
rect 11081 2144 11145 2148
rect 15786 2204 15850 2208
rect 15786 2148 15790 2204
rect 15790 2148 15846 2204
rect 15846 2148 15850 2204
rect 15786 2144 15850 2148
rect 15866 2204 15930 2208
rect 15866 2148 15870 2204
rect 15870 2148 15926 2204
rect 15926 2148 15930 2204
rect 15866 2144 15930 2148
rect 15946 2204 16010 2208
rect 15946 2148 15950 2204
rect 15950 2148 16006 2204
rect 16006 2148 16010 2204
rect 15946 2144 16010 2148
rect 16026 2204 16090 2208
rect 16026 2148 16030 2204
rect 16030 2148 16086 2204
rect 16086 2148 16090 2204
rect 16026 2144 16090 2148
rect 20731 2204 20795 2208
rect 20731 2148 20735 2204
rect 20735 2148 20791 2204
rect 20791 2148 20795 2204
rect 20731 2144 20795 2148
rect 20811 2204 20875 2208
rect 20811 2148 20815 2204
rect 20815 2148 20871 2204
rect 20871 2148 20875 2204
rect 20811 2144 20875 2148
rect 20891 2204 20955 2208
rect 20891 2148 20895 2204
rect 20895 2148 20951 2204
rect 20951 2148 20955 2204
rect 20891 2144 20955 2148
rect 20971 2204 21035 2208
rect 20971 2148 20975 2204
rect 20975 2148 21031 2204
rect 21031 2148 21035 2204
rect 20971 2144 21035 2148
<< metal4 >>
rect 3416 19072 3736 19632
rect 3416 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3736 19072
rect 3416 17984 3736 19008
rect 3416 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3736 17984
rect 3416 16896 3736 17920
rect 3416 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3736 16896
rect 3416 15808 3736 16832
rect 3416 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3736 15808
rect 3416 14720 3736 15744
rect 3416 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3736 14720
rect 3416 13632 3736 14656
rect 3416 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3736 13632
rect 3416 12544 3736 13568
rect 3416 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3736 12544
rect 3416 11456 3736 12480
rect 3416 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3736 11456
rect 3416 10368 3736 11392
rect 3416 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3736 10368
rect 3416 9280 3736 10304
rect 3416 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3736 9280
rect 3416 8192 3736 9216
rect 3416 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3736 8192
rect 3416 7104 3736 8128
rect 3416 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3736 7104
rect 3416 6016 3736 7040
rect 3416 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3736 6016
rect 3416 4928 3736 5952
rect 3416 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3736 4928
rect 3416 3840 3736 4864
rect 3416 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3736 3840
rect 3416 2752 3736 3776
rect 3416 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3736 2752
rect 3416 2128 3736 2688
rect 5888 19616 6208 19632
rect 5888 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6208 19616
rect 5888 18528 6208 19552
rect 5888 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6208 18528
rect 5888 17440 6208 18464
rect 5888 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6208 17440
rect 5888 16352 6208 17376
rect 5888 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6208 16352
rect 5888 15264 6208 16288
rect 5888 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6208 15264
rect 5888 14176 6208 15200
rect 5888 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6208 14176
rect 5888 13088 6208 14112
rect 5888 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6208 13088
rect 5888 12000 6208 13024
rect 5888 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6208 12000
rect 5888 10912 6208 11936
rect 5888 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6208 10912
rect 5888 9824 6208 10848
rect 5888 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6208 9824
rect 5888 8736 6208 9760
rect 5888 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6208 8736
rect 5888 7648 6208 8672
rect 5888 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6208 7648
rect 5888 6560 6208 7584
rect 5888 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6208 6560
rect 5888 5472 6208 6496
rect 5888 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6208 5472
rect 5888 4384 6208 5408
rect 5888 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6208 4384
rect 5888 3296 6208 4320
rect 5888 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6208 3296
rect 5888 2208 6208 3232
rect 5888 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6208 2208
rect 5888 2128 6208 2144
rect 8361 19072 8681 19632
rect 8361 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8681 19072
rect 8361 17984 8681 19008
rect 8361 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8681 17984
rect 8361 16896 8681 17920
rect 8361 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8681 16896
rect 8361 15808 8681 16832
rect 8361 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8681 15808
rect 8361 14720 8681 15744
rect 8361 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8681 14720
rect 8361 13632 8681 14656
rect 8361 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8681 13632
rect 8361 12544 8681 13568
rect 8361 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8681 12544
rect 8361 11456 8681 12480
rect 8361 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8681 11456
rect 8361 10368 8681 11392
rect 8361 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8681 10368
rect 8361 9280 8681 10304
rect 8361 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8681 9280
rect 8361 8192 8681 9216
rect 8361 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8681 8192
rect 8361 7104 8681 8128
rect 8361 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8681 7104
rect 8361 6016 8681 7040
rect 8361 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8681 6016
rect 8361 4928 8681 5952
rect 8361 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8681 4928
rect 8361 3840 8681 4864
rect 8361 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8681 3840
rect 8361 2752 8681 3776
rect 8361 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8681 2752
rect 8361 2128 8681 2688
rect 10833 19616 11153 19632
rect 10833 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11153 19616
rect 10833 18528 11153 19552
rect 10833 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11153 18528
rect 10833 17440 11153 18464
rect 10833 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11153 17440
rect 10833 16352 11153 17376
rect 10833 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11153 16352
rect 10833 15264 11153 16288
rect 10833 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11153 15264
rect 10833 14176 11153 15200
rect 10833 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11153 14176
rect 10833 13088 11153 14112
rect 10833 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11153 13088
rect 10833 12000 11153 13024
rect 10833 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11153 12000
rect 10833 10912 11153 11936
rect 10833 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11153 10912
rect 10833 9824 11153 10848
rect 10833 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11153 9824
rect 10833 8736 11153 9760
rect 10833 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11153 8736
rect 10833 7648 11153 8672
rect 10833 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11153 7648
rect 10833 6560 11153 7584
rect 10833 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11153 6560
rect 10833 5472 11153 6496
rect 10833 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11153 5472
rect 10833 4384 11153 5408
rect 10833 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11153 4384
rect 10833 3296 11153 4320
rect 10833 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11153 3296
rect 10833 2208 11153 3232
rect 10833 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11153 2208
rect 10833 2128 11153 2144
rect 13306 19072 13626 19632
rect 13306 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13626 19072
rect 13306 17984 13626 19008
rect 13306 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13626 17984
rect 13306 16896 13626 17920
rect 13306 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13626 16896
rect 13306 15808 13626 16832
rect 13306 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13626 15808
rect 13306 14720 13626 15744
rect 13306 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13626 14720
rect 13306 13632 13626 14656
rect 13306 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13626 13632
rect 13306 12544 13626 13568
rect 13306 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13626 12544
rect 13306 11456 13626 12480
rect 13306 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13626 11456
rect 13306 10368 13626 11392
rect 13306 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13626 10368
rect 13306 9280 13626 10304
rect 13306 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13626 9280
rect 13306 8192 13626 9216
rect 13306 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13626 8192
rect 13306 7104 13626 8128
rect 13306 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13626 7104
rect 13306 6016 13626 7040
rect 13306 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13626 6016
rect 13306 4928 13626 5952
rect 13306 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13626 4928
rect 13306 3840 13626 4864
rect 13306 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13626 3840
rect 13306 2752 13626 3776
rect 13306 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13626 2752
rect 13306 2128 13626 2688
rect 15778 19616 16098 19632
rect 15778 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16098 19616
rect 15778 18528 16098 19552
rect 15778 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16098 18528
rect 15778 17440 16098 18464
rect 15778 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16098 17440
rect 15778 16352 16098 17376
rect 15778 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16098 16352
rect 15778 15264 16098 16288
rect 15778 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16098 15264
rect 15778 14176 16098 15200
rect 15778 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16098 14176
rect 15778 13088 16098 14112
rect 15778 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16098 13088
rect 15778 12000 16098 13024
rect 15778 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16098 12000
rect 15778 10912 16098 11936
rect 15778 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16098 10912
rect 15778 9824 16098 10848
rect 15778 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16098 9824
rect 15778 8736 16098 9760
rect 15778 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16098 8736
rect 15778 7648 16098 8672
rect 15778 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16098 7648
rect 15778 6560 16098 7584
rect 15778 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16098 6560
rect 15778 5472 16098 6496
rect 15778 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16098 5472
rect 15778 4384 16098 5408
rect 15778 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16098 4384
rect 15778 3296 16098 4320
rect 15778 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16098 3296
rect 15778 2208 16098 3232
rect 15778 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16098 2208
rect 15778 2128 16098 2144
rect 18251 19072 18571 19632
rect 18251 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18571 19072
rect 18251 17984 18571 19008
rect 18251 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18571 17984
rect 18251 16896 18571 17920
rect 18251 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18571 16896
rect 18251 15808 18571 16832
rect 18251 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18571 15808
rect 18251 14720 18571 15744
rect 18251 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18571 14720
rect 18251 13632 18571 14656
rect 18251 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18571 13632
rect 18251 12544 18571 13568
rect 18251 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18571 12544
rect 18251 11456 18571 12480
rect 18251 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18571 11456
rect 18251 10368 18571 11392
rect 18251 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18571 10368
rect 18251 9280 18571 10304
rect 18251 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18571 9280
rect 18251 8192 18571 9216
rect 18251 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18571 8192
rect 18251 7104 18571 8128
rect 18251 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18571 7104
rect 18251 6016 18571 7040
rect 18251 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18571 6016
rect 18251 4928 18571 5952
rect 18251 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18571 4928
rect 18251 3840 18571 4864
rect 18251 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18571 3840
rect 18251 2752 18571 3776
rect 18251 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18571 2752
rect 18251 2128 18571 2688
rect 20723 19616 21043 19632
rect 20723 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21043 19616
rect 20723 18528 21043 19552
rect 20723 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21043 18528
rect 20723 17440 21043 18464
rect 20723 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21043 17440
rect 20723 16352 21043 17376
rect 20723 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21043 16352
rect 20723 15264 21043 16288
rect 20723 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21043 15264
rect 20723 14176 21043 15200
rect 20723 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21043 14176
rect 20723 13088 21043 14112
rect 20723 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21043 13088
rect 20723 12000 21043 13024
rect 20723 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21043 12000
rect 20723 10912 21043 11936
rect 20723 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21043 10912
rect 20723 9824 21043 10848
rect 20723 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21043 9824
rect 20723 8736 21043 9760
rect 20723 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21043 8736
rect 20723 7648 21043 8672
rect 20723 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21043 7648
rect 20723 6560 21043 7584
rect 20723 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21043 6560
rect 20723 5472 21043 6496
rect 20723 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21043 5472
rect 20723 4384 21043 5408
rect 20723 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21043 4384
rect 20723 3296 21043 4320
rect 20723 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21043 3296
rect 20723 2208 21043 3232
rect 20723 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21043 2208
rect 20723 2128 21043 2144
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99
timestamp 1676037725
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_157
timestamp 1676037725
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_186
timestamp 1676037725
transform 1 0 18216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1676037725
transform 1 0 19780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_33
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_211
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1676037725
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_37
timestamp 1676037725
transform 1 0 4508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1676037725
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1676037725
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1676037725
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1676037725
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1676037725
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1676037725
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_156
timestamp 1676037725
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_168
timestamp 1676037725
transform 1 0 16560 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1676037725
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_13
timestamp 1676037725
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_25
timestamp 1676037725
transform 1 0 3404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1676037725
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1676037725
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_90
timestamp 1676037725
transform 1 0 9384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1676037725
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1676037725
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1676037725
transform 1 0 12880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1676037725
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1676037725
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_194
timestamp 1676037725
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_206
timestamp 1676037725
transform 1 0 20056 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1676037725
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_50
timestamp 1676037725
transform 1 0 5704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_54
timestamp 1676037725
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1676037725
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_105
timestamp 1676037725
transform 1 0 10764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_123
timestamp 1676037725
transform 1 0 12420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1676037725
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1676037725
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_148
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_156
timestamp 1676037725
transform 1 0 15456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_166
timestamp 1676037725
transform 1 0 16376 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_172
timestamp 1676037725
transform 1 0 16928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1676037725
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1676037725
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_32
timestamp 1676037725
transform 1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1676037725
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_75
timestamp 1676037725
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1676037725
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_122
timestamp 1676037725
transform 1 0 12328 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1676037725
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_143
timestamp 1676037725
transform 1 0 14260 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1676037725
transform 1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1676037725
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_184
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_196
timestamp 1676037725
transform 1 0 19136 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1676037725
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_49
timestamp 1676037725
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_58
timestamp 1676037725
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_70
timestamp 1676037725
transform 1 0 7544 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_107
timestamp 1676037725
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_119
timestamp 1676037725
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_154
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_166
timestamp 1676037725
transform 1 0 16376 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_175
timestamp 1676037725
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1676037725
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_33
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1676037725
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_70
timestamp 1676037725
transform 1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_83
timestamp 1676037725
transform 1 0 8740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1676037725
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1676037725
transform 1 0 12420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1676037725
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_180
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_192
timestamp 1676037725
transform 1 0 18768 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_204
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1676037725
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1676037725
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1676037725
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_50
timestamp 1676037725
transform 1 0 5704 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_56
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1676037725
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1676037725
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_94
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1676037725
transform 1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_111
timestamp 1676037725
transform 1 0 11316 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1676037725
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1676037725
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1676037725
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_154
timestamp 1676037725
transform 1 0 15272 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1676037725
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_179
timestamp 1676037725
transform 1 0 17572 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_187
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1676037725
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_16
timestamp 1676037725
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_82
timestamp 1676037725
transform 1 0 8648 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_94
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1676037725
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_126
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_138
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1676037725
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1676037725
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_186
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1676037725
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1676037725
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1676037725
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1676037725
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1676037725
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_164
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_180
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_202
timestamp 1676037725
transform 1 0 19688 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1676037725
transform 1 0 20424 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_133
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_183
timestamp 1676037725
transform 1 0 17940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_195
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_202
timestamp 1676037725
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_167
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_173
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_14
timestamp 1676037725
transform 1 0 2392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_26
timestamp 1676037725
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1676037725
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_200
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1676037725
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1676037725
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 1676037725
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_103
timestamp 1676037725
transform 1 0 10580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_115
timestamp 1676037725
transform 1 0 11684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_156
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_14
timestamp 1676037725
transform 1 0 2392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1676037725
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1676037725
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1676037725
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_102
timestamp 1676037725
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_134
timestamp 1676037725
transform 1 0 13432 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1676037725
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1676037725
transform 1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_203
timestamp 1676037725
transform 1 0 19780 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1676037725
transform 1 0 20516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1676037725
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1676037725
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_50
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_62
timestamp 1676037725
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1676037725
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1676037725
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_123
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_155
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_206
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_12
timestamp 1676037725
transform 1 0 2208 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_24
timestamp 1676037725
transform 1 0 3312 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1676037725
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_75
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_87
timestamp 1676037725
transform 1 0 9108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_99
timestamp 1676037725
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_132
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_184
timestamp 1676037725
transform 1 0 18032 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1676037725
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1676037725
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1676037725
transform 1 0 2392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_47
timestamp 1676037725
transform 1 0 5428 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1676037725
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1676037725
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1676037725
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_16
timestamp 1676037725
transform 1 0 2576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1676037725
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_132
timestamp 1676037725
transform 1 0 13248 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_144
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_156
timestamp 1676037725
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_192
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1676037725
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_12
timestamp 1676037725
transform 1 0 2208 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1676037725
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_47
timestamp 1676037725
transform 1 0 5428 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1676037725
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1676037725
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1676037725
transform 1 0 16560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1676037725
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_206
timestamp 1676037725
transform 1 0 20056 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_145
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1676037725
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_186
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1676037725
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_16
timestamp 1676037725
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_173
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1676037725
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1676037725
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 1676037725
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1676037725
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_14
timestamp 1676037725
transform 1 0 2392 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_26
timestamp 1676037725
transform 1 0 3496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1676037725
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1676037725
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_134
timestamp 1676037725
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_155
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_180
timestamp 1676037725
transform 1 0 17664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_202
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1676037725
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_12
timestamp 1676037725
transform 1 0 2208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1676037725
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_105
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_185
timestamp 1676037725
transform 1 0 18124 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1676037725
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_24
timestamp 1676037725
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1676037725
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1676037725
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_178
timestamp 1676037725
transform 1 0 17480 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_190
timestamp 1676037725
transform 1 0 18584 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_16
timestamp 1676037725
transform 1 0 2576 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_47
timestamp 1676037725
transform 1 0 5428 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 1676037725
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_63
timestamp 1676037725
transform 1 0 6900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1676037725
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1676037725
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1676037725
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1676037725
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_155
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_167
timestamp 1676037725
transform 1 0 16468 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1676037725
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_180
timestamp 1676037725
transform 1 0 17664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1676037725
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_17
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_70
timestamp 1676037725
transform 1 0 7544 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_90
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_102
timestamp 1676037725
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1676037725
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1676037725
transform 1 0 15364 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_185
timestamp 1676037725
transform 1 0 18124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_197
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_209
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1676037725
transform 1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_49
timestamp 1676037725
transform 1 0 5612 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_66
timestamp 1676037725
transform 1 0 7176 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1676037725
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1676037725
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1676037725
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_78
timestamp 1676037725
transform 1 0 8280 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_132
timestamp 1676037725
transform 1 0 13248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_141
timestamp 1676037725
transform 1 0 14076 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_150
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_175
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_203
timestamp 1676037725
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1676037725
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1676037725
transform -1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1676037725
transform 1 0 15640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1676037725
transform 1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1676037725
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4140 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2760 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _193_
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18308 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _198_
timestamp 1676037725
transform -1 0 17388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 1676037725
transform 1 0 14904 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_4  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform -1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15640 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _209_
timestamp 1676037725
transform -1 0 15456 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15640 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _212_
timestamp 1676037725
transform -1 0 17480 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _213_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1676037725
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _218_
timestamp 1676037725
transform -1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15916 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ai_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14628 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _225_
timestamp 1676037725
transform -1 0 15272 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _229_
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _231_
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18584 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _233_
timestamp 1676037725
transform 1 0 18124 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1676037725
transform -1 0 5244 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1676037725
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 1676037725
transform -1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _239_
timestamp 1676037725
transform 1 0 5612 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _240_
timestamp 1676037725
transform 1 0 8096 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_4  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1676037725
transform -1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1676037725
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _248_
timestamp 1676037725
transform -1 0 8648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9384 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _250_
timestamp 1676037725
transform 1 0 8004 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 1676037725
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1676037725
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1676037725
transform 1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _257_
timestamp 1676037725
transform -1 0 6440 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1676037725
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _260_
timestamp 1676037725
transform -1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1676037725
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1676037725
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _263_
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _267_
timestamp 1676037725
transform -1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _268_
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1676037725
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _270_
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _273_
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _274_
timestamp 1676037725
transform -1 0 14720 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp 1676037725
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12972 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _277_
timestamp 1676037725
transform 1 0 12972 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _279_
timestamp 1676037725
transform 1 0 11776 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13892 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and4_2  _284_
timestamp 1676037725
transform -1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _286_
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _289_
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1676037725
transform -1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _291_
timestamp 1676037725
transform -1 0 12696 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _292_
timestamp 1676037725
transform 1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _295_
timestamp 1676037725
transform -1 0 19964 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1676037725
transform -1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _297_
timestamp 1676037725
transform 1 0 16928 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp 1676037725
transform -1 0 17572 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _300_
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _301_
timestamp 1676037725
transform -1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _302_
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1676037725
transform -1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _304_
timestamp 1676037725
transform -1 0 17940 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _305_
timestamp 1676037725
transform -1 0 18308 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1676037725
transform -1 0 19504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20056 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _309_
timestamp 1676037725
transform -1 0 19780 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _310_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _311_
timestamp 1676037725
transform -1 0 20056 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _312_
timestamp 1676037725
transform -1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 1676037725
transform -1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _314_
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _315_
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _316_
timestamp 1676037725
transform -1 0 20240 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _317_
timestamp 1676037725
transform -1 0 20056 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1676037725
transform -1 0 19412 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _320_
timestamp 1676037725
transform -1 0 17572 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _321_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1676037725
transform -1 0 18216 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _323_
timestamp 1676037725
transform 1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _324_
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _325_
timestamp 1676037725
transform -1 0 20148 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _327_
timestamp 1676037725
transform -1 0 17572 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _328_
timestamp 1676037725
transform -1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _330_
timestamp 1676037725
transform 1 0 16928 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _331_
timestamp 1676037725
transform -1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _332_
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1676037725
transform -1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _334_
timestamp 1676037725
transform -1 0 18032 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _335_
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _336_
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16100 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _340_
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _342_
timestamp 1676037725
transform -1 0 14904 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _344_
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _345_
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform -1 0 3404 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 1676037725
transform -1 0 2576 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 1676037725
transform -1 0 14996 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _349_
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _350_
timestamp 1676037725
transform -1 0 2668 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1676037725
transform 1 0 2024 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _352_
timestamp 1676037725
transform 1 0 2852 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _353_
timestamp 1676037725
transform 1 0 1840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _354_
timestamp 1676037725
transform -1 0 2392 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1676037725
transform 1 0 1840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _357_
timestamp 1676037725
transform -1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _358_
timestamp 1676037725
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _359_
timestamp 1676037725
transform -1 0 2392 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 1676037725
transform 1 0 2760 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8648 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5704 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _364_
timestamp 1676037725
transform -1 0 5520 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5520 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1676037725
transform -1 0 8004 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1676037725
transform 1 0 6440 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _374_
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _375_
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _376_
timestamp 1676037725
transform 1 0 6716 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _377_
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _378_
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _379_
timestamp 1676037725
transform 1 0 8740 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _381_
timestamp 1676037725
transform 1 0 9752 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _382_
timestamp 1676037725
transform 1 0 11776 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1676037725
transform 1 0 11776 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1676037725
transform 1 0 7636 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _390_
timestamp 1676037725
transform 1 0 9200 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1676037725
transform 1 0 9108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1676037725
transform 1 0 11776 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _394_
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1676037725
transform 1 0 9568 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1676037725
transform 1 0 11776 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _397_
timestamp 1676037725
transform -1 0 5704 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _398_
timestamp 1676037725
transform -1 0 5612 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _399_
timestamp 1676037725
transform -1 0 5336 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform -1 0 5428 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1676037725
transform -1 0 5244 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1676037725
transform -1 0 8464 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform 1 0 5704 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform -1 0 5428 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform -1 0 8004 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform -1 0 5428 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform -1 0 8004 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform -1 0 7452 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1676037725
transform -1 0 5428 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1676037725
transform -1 0 8004 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform -1 0 5428 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 6900 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5336 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1676037725
transform 1 0 19504 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout15
timestamp 1676037725
transform -1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout17
timestamp 1676037725
transform -1 0 8280 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1676037725
transform -1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1676037725
transform -1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform -1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform -1 0 11224 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output3
timestamp 1676037725
transform -1 0 2208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1676037725
transform -1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform -1 0 7544 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 17664 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 19872 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 3698 21200 3754 22000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 18234 21200 18290 22000 0 FreeSans 224 90 0 0 io_in
port 1 nsew signal input
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 io_out[0]
port 2 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 io_out[1]
port 3 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 io_out[2]
port 4 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 io_out[3]
port 5 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_out[4]
port 6 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_out[5]
port 7 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 io_out[6]
port 8 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[7]
port 9 nsew signal tristate
flabel metal2 s 10966 21200 11022 22000 0 FreeSans 224 90 0 0 rst
port 10 nsew signal input
flabel metal4 s 3416 2128 3736 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 8361 2128 8681 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 13306 2128 13626 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 18251 2128 18571 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 5888 2128 6208 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 10833 2128 11153 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 15778 2128 16098 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 20723 2128 21043 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
<< end >>
